module d01_example_adder (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire _07_;
	wire _08_;
	wire _09_;
	wire _10_;
	wire _11_;
	wire _12_;
	wire _13_;
	wire _14_;
	wire _15_;
	wire _16_;
	wire _17_;
	wire _18_;
	wire _19_;
	wire _20_;
	wire _21_;
	wire _22_;
	wire _23_;
	wire _24_;
	wire _25_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _00_ = io_in[5] ^ io_in[11];
	assign _01_ = ~(io_in[4] ^ io_in[10]);
	assign _02_ = _00_ & ~_01_;
	assign _03_ = ~(io_in[3] & io_in[9]);
	assign _04_ = io_in[3] ^ io_in[9];
	assign _05_ = ~(io_in[2] & io_in[8]);
	assign _06_ = _04_ & ~_05_;
	assign _07_ = _03_ & ~_06_;
	assign _08_ = ~(io_in[2] ^ io_in[8]);
	assign _09_ = _04_ & ~_08_;
	assign _10_ = ~(io_in[1] & io_in[7]);
	assign _11_ = io_in[1] ^ io_in[7];
	assign _12_ = ~(io_in[0] & io_in[6]);
	assign _13_ = _11_ & ~_12_;
	assign _14_ = _10_ & ~_13_;
	assign _15_ = _09_ & ~_14_;
	assign _16_ = _07_ & ~_15_;
	assign _17_ = _02_ & ~_16_;
	assign _18_ = ~(io_in[4] & io_in[10]);
	assign _19_ = _00_ & ~_18_;
	assign _20_ = io_in[5] & io_in[11];
	assign _21_ = _20_ | _19_;
	assign io_out[6] = _21_ | _17_;
	assign io_out[1] = ~(_12_ ^ _11_);
	assign io_out[2] = _14_ ^ _08_;
	assign _22_ = ~(_14_ | _08_);
	assign _23_ = _22_ | ~_05_;
	assign io_out[3] = _23_ ^ _04_;
	assign io_out[4] = _16_ ^ _01_;
	assign _24_ = ~(_16_ | _01_);
	assign _25_ = _24_ | ~_18_;
	assign io_out[5] = _25_ ^ _00_;
	assign io_out[0] = io_in[0] ^ io_in[6];
	assign io_out[13:7] = 7'h00;
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {5'h00, io_out[6:0]};
	assign \mchip.reset  = io_in[13];
endmodule
module d02_example_counter (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire [11:0] _059_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire \mchip.enable ;
	wire [11:0] \mchip.io_in ;
	reg [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire \mchip.updown ;
	assign _059_[0] = ~\mchip.io_out [0];
	assign _001_ = ~(io_in[1] & io_in[0]);
	assign _002_ = io_in[1] | ~io_in[0];
	assign _000_ = ~(_002_ & _001_);
	assign _003_ = _001_ ^ \mchip.io_out [1];
	assign _059_[1] = _003_ ^ _059_[0];
	assign _004_ = \mchip.io_out [1] & ~_001_;
	assign _005_ = \mchip.io_out [0] & ~_003_;
	assign _006_ = _005_ | _004_;
	assign _007_ = _001_ ^ \mchip.io_out [2];
	assign _059_[2] = ~(_007_ ^ _006_);
	assign _008_ = \mchip.io_out [2] & ~_001_;
	assign _009_ = _006_ & ~_007_;
	assign _010_ = ~(_009_ | _008_);
	assign _011_ = _001_ ^ \mchip.io_out [3];
	assign _059_[3] = _011_ ^ _010_;
	assign _012_ = _011_ | _007_;
	assign _013_ = _006_ & ~_012_;
	assign _014_ = \mchip.io_out [3] & ~_001_;
	assign _015_ = _008_ & ~_011_;
	assign _016_ = _015_ | _014_;
	assign _017_ = _016_ | _013_;
	assign _018_ = _001_ ^ \mchip.io_out [4];
	assign _059_[4] = ~(_018_ ^ _017_);
	assign _019_ = \mchip.io_out [4] & ~_001_;
	assign _020_ = _017_ & ~_018_;
	assign _021_ = ~(_020_ | _019_);
	assign _022_ = _001_ ^ \mchip.io_out [5];
	assign _059_[5] = _022_ ^ _021_;
	assign _023_ = _022_ | _018_;
	assign _024_ = _017_ & ~_023_;
	assign _025_ = \mchip.io_out [5] & ~_001_;
	assign _026_ = _019_ & ~_022_;
	assign _027_ = _026_ | _025_;
	assign _028_ = _027_ | _024_;
	assign _029_ = _001_ ^ \mchip.io_out [6];
	assign _059_[6] = ~(_029_ ^ _028_);
	assign _030_ = \mchip.io_out [6] & ~_001_;
	assign _031_ = _028_ & ~_029_;
	assign _032_ = ~(_031_ | _030_);
	assign _033_ = _001_ ^ \mchip.io_out [7];
	assign _059_[7] = _033_ ^ _032_;
	assign _034_ = \mchip.io_out [7] & ~_001_;
	assign _035_ = _030_ & ~_033_;
	assign _036_ = _035_ | _034_;
	assign _037_ = _033_ | _029_;
	assign _038_ = _027_ & ~_037_;
	assign _039_ = _038_ | _036_;
	assign _040_ = _037_ | _023_;
	assign _041_ = _017_ & ~_040_;
	assign _042_ = _041_ | _039_;
	assign _043_ = ~(_001_ ^ \mchip.io_out [8]);
	assign _059_[8] = _043_ ^ _042_;
	assign _044_ = \mchip.io_out [8] & ~_001_;
	assign _045_ = _043_ & _042_;
	assign _046_ = _045_ | _044_;
	assign _047_ = ~(_001_ ^ \mchip.io_out [9]);
	assign _059_[9] = _047_ ^ _046_;
	assign _048_ = \mchip.io_out [9] & ~_001_;
	assign _049_ = _047_ & _044_;
	assign _050_ = _049_ | _048_;
	assign _051_ = ~(_047_ & _043_);
	assign _052_ = _042_ & ~_051_;
	assign _053_ = _052_ | _050_;
	assign _054_ = ~(_001_ ^ \mchip.io_out [10]);
	assign _059_[10] = _054_ ^ _053_;
	assign _055_ = \mchip.io_out [10] & ~_001_;
	assign _056_ = _054_ & _053_;
	assign _057_ = _056_ | _055_;
	assign _058_ = ~(_001_ ^ \mchip.io_out [11]);
	assign _059_[11] = _058_ ^ _057_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [0] <= 1'h0;
		else if (_000_)
			\mchip.io_out [0] <= _059_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [1] <= 1'h0;
		else if (_000_)
			\mchip.io_out [1] <= _059_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [2] <= 1'h0;
		else if (_000_)
			\mchip.io_out [2] <= _059_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [3] <= 1'h0;
		else if (_000_)
			\mchip.io_out [3] <= _059_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [4] <= 1'h0;
		else if (_000_)
			\mchip.io_out [4] <= _059_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [5] <= 1'h0;
		else if (_000_)
			\mchip.io_out [5] <= _059_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [6] <= 1'h0;
		else if (_000_)
			\mchip.io_out [6] <= _059_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [7] <= 1'h0;
		else if (_000_)
			\mchip.io_out [7] <= _059_[7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [8] <= 1'h0;
		else if (_000_)
			\mchip.io_out [8] <= _059_[8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [9] <= 1'h0;
		else if (_000_)
			\mchip.io_out [9] <= _059_[9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [10] <= 1'h0;
		else if (_000_)
			\mchip.io_out [10] <= _059_[10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [11] <= 1'h0;
		else if (_000_)
			\mchip.io_out [11] <= _059_[11];
	assign io_out = {2'h0, \mchip.io_out };
	assign \mchip.clock  = io_in[12];
	assign \mchip.enable  = io_in[0];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.reset  = io_in[13];
	assign \mchip.updown  = io_in[1];
endmodule
module d03_example_iotest (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire [3:0] _091_;
	wire [3:0] _092_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	reg [3:0] \mchip.idx ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire [11:0] \mchip.shift_bit ;
	assign _091_[0] = ~\mchip.idx [0];
	assign _035_ = \mchip.idx [1] & \mchip.idx [0];
	assign _036_ = \mchip.idx [2] | ~\mchip.idx [3];
	assign _037_ = _035_ & ~_036_;
	assign _000_ = _037_ | io_in[13];
	assign _038_ = ~(\mchip.idx [3] | \mchip.idx [2]);
	assign _039_ = \mchip.idx [1] | \mchip.idx [0];
	assign _040_ = _038_ & ~_039_;
	assign _041_ = ~\mchip.idx [2];
	assign _042_ = _041_ & ~_039_;
	assign _043_ = _042_ ^ \mchip.idx [3];
	assign _044_ = _039_ ^ _041_;
	assign _045_ = \mchip.idx [1] | ~\mchip.idx [0];
	assign _046_ = _045_ | _044_;
	assign _047_ = ~(_046_ | _043_);
	assign _048_ = _047_ & ~_040_;
	assign io_out[0] = _048_ & ~_040_;
	assign _049_ = io_in[6] ^ io_in[7];
	assign _050_ = io_in[4] ^ io_in[5];
	assign _051_ = _050_ ^ _049_;
	assign _052_ = ~_040_;
	assign _053_ = ~_044_;
	assign _054_ = _039_ & ~_035_;
	assign _055_ = _040_ | \mchip.idx [0];
	assign _056_ = _055_ | _054_;
	assign _057_ = _056_ | _053_;
	assign _058_ = _057_ | _043_;
	assign _059_ = _058_ | _040_;
	assign _060_ = _052_ & ~_059_;
	assign io_out[7] = _060_ ^ _051_;
	assign _061_ = io_in[2] ^ io_in[3];
	assign _062_ = io_in[0] ^ io_in[1];
	assign _063_ = _062_ ^ _061_;
	assign _064_ = _063_ ^ _050_;
	assign _065_ = \mchip.idx [0] | ~\mchip.idx [1];
	assign _066_ = _065_ | _044_;
	assign _067_ = _066_ | ~_043_;
	assign _068_ = _067_ | _040_;
	assign _069_ = _052_ & ~_068_;
	assign io_out[9] = _069_ ^ _064_;
	assign _070_ = io_in[10] ^ io_in[11];
	assign _071_ = io_in[8] ^ io_in[9];
	assign _072_ = _071_ ^ _070_;
	assign _073_ = _072_ ^ _063_;
	assign _074_ = ~(\mchip.idx [1] & \mchip.idx [0]);
	assign _075_ = _074_ | ~_044_;
	assign _076_ = _075_ | _043_;
	assign _077_ = _076_ | _040_;
	assign _078_ = _052_ & ~_077_;
	assign io_out[6] = _078_ ^ _073_;
	assign _079_ = _072_ ^ _049_;
	assign _080_ = _046_ | ~_043_;
	assign _081_ = _080_ | _040_;
	assign _082_ = _052_ & ~_081_;
	assign io_out[8] = _082_ ^ _079_;
	assign _083_ = _062_ ^ _050_;
	assign _084_ = _083_ ^ _071_;
	assign _085_ = _065_ | ~_044_;
	assign _086_ = _085_ | _043_;
	assign _087_ = _086_ | _040_;
	assign _088_ = _052_ & ~_087_;
	assign io_out[5] = _088_ ^ _084_;
	assign _089_ = _061_ ^ _049_;
	assign _090_ = _089_ ^ _070_;
	assign _001_ = _045_ | ~_044_;
	assign _002_ = _001_ | _043_;
	assign _003_ = _002_ | _040_;
	assign _004_ = _052_ & ~_003_;
	assign io_out[4] = _004_ ^ _090_;
	assign _005_ = _074_ | _044_;
	assign _006_ = _005_ | ~_043_;
	assign _007_ = _006_ | _040_;
	assign _008_ = _052_ & ~_007_;
	assign io_out[10] = _008_ ^ _072_;
	assign _009_ = ~(io_in[10] ^ io_in[8]);
	assign _010_ = ~(io_in[6] ^ io_in[4]);
	assign _011_ = io_in[2] ^ io_in[0];
	assign _012_ = _011_ ^ _010_;
	assign _013_ = _012_ ^ _009_;
	assign _014_ = _056_ | _044_;
	assign _015_ = _014_ | _043_;
	assign _016_ = _015_ | _040_;
	assign _017_ = _052_ & ~_016_;
	assign io_out[3] = _017_ ^ _013_;
	assign _018_ = ~(io_in[11] ^ io_in[9]);
	assign _019_ = ~(io_in[7] ^ io_in[5]);
	assign _020_ = io_in[3] ^ io_in[1];
	assign _021_ = _020_ ^ _019_;
	assign _022_ = _021_ ^ _018_;
	assign _023_ = _005_ | _043_;
	assign _024_ = _023_ | _040_;
	assign _025_ = _052_ & ~_024_;
	assign io_out[2] = _025_ ^ _022_;
	assign _026_ = _063_ ^ _051_;
	assign _027_ = _026_ ^ _072_;
	assign _028_ = _066_ | _043_;
	assign _029_ = _028_ | _040_;
	assign _030_ = _052_ & ~_029_;
	assign io_out[1] = _030_ ^ _027_;
	assign _031_ = _014_ | ~_043_;
	assign _032_ = _031_ | _040_;
	assign _033_ = _052_ & ~_032_;
	assign io_out[11] = _033_ ^ _051_;
	assign _092_[1] = \mchip.idx [1] ^ \mchip.idx [0];
	assign _092_[2] = _035_ ^ \mchip.idx [2];
	assign _034_ = _035_ & ~_041_;
	assign _092_[3] = _034_ ^ \mchip.idx [3];
	always @(posedge io_in[12])
		if (_000_)
			\mchip.idx [0] <= 1'h0;
		else
			\mchip.idx [0] <= _091_[0];
	always @(posedge io_in[12])
		if (_000_)
			\mchip.idx [1] <= 1'h0;
		else
			\mchip.idx [1] <= _092_[1];
	always @(posedge io_in[12])
		if (_000_)
			\mchip.idx [2] <= 1'h0;
		else
			\mchip.idx [2] <= _092_[2];
	always @(posedge io_in[12])
		if (_000_)
			\mchip.idx [3] <= 1'h0;
		else
			\mchip.idx [3] <= _092_[3];
	assign _091_[3:1] = \mchip.idx [3:1];
	assign _092_[0] = _091_[0];
	assign io_out[13:12] = 2'h0;
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = io_out[11:0];
	assign \mchip.reset  = io_in[13];
	assign \mchip.shift_bit  = {11'h000, io_out[0]};
endmodule
module d05_meta_info (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire _2025_;
	wire _2026_;
	wire _2027_;
	wire _2028_;
	wire _2029_;
	wire _2030_;
	wire _2031_;
	wire _2032_;
	wire _2033_;
	wire _2034_;
	wire _2035_;
	wire _2036_;
	wire _2037_;
	wire _2038_;
	wire _2039_;
	wire _2040_;
	wire _2041_;
	wire _2042_;
	wire _2043_;
	wire _2044_;
	wire _2045_;
	wire _2046_;
	wire _2047_;
	wire _2048_;
	wire _2049_;
	wire _2050_;
	wire _2051_;
	wire _2052_;
	wire _2053_;
	wire _2054_;
	wire _2055_;
	wire _2056_;
	wire _2057_;
	wire _2058_;
	wire _2059_;
	wire _2060_;
	wire _2061_;
	wire _2062_;
	wire _2063_;
	wire _2064_;
	wire _2065_;
	wire _2066_;
	wire _2067_;
	wire _2068_;
	wire _2069_;
	wire _2070_;
	wire _2071_;
	wire _2072_;
	wire _2073_;
	wire _2074_;
	wire _2075_;
	wire _2076_;
	wire _2077_;
	wire _2078_;
	wire _2079_;
	wire _2080_;
	wire _2081_;
	wire _2082_;
	wire _2083_;
	wire _2084_;
	wire _2085_;
	wire _2086_;
	wire _2087_;
	wire _2088_;
	wire _2089_;
	wire _2090_;
	wire _2091_;
	wire _2092_;
	wire _2093_;
	wire _2094_;
	wire _2095_;
	wire _2096_;
	wire _2097_;
	wire _2098_;
	wire _2099_;
	wire _2100_;
	wire _2101_;
	wire _2102_;
	wire _2103_;
	wire _2104_;
	wire _2105_;
	wire _2106_;
	wire _2107_;
	wire _2108_;
	wire _2109_;
	wire _2110_;
	wire _2111_;
	wire _2112_;
	wire _2113_;
	wire _2114_;
	wire _2115_;
	wire _2116_;
	wire _2117_;
	wire _2118_;
	wire _2119_;
	wire _2120_;
	wire _2121_;
	wire _2122_;
	wire _2123_;
	wire _2124_;
	wire _2125_;
	wire _2126_;
	wire _2127_;
	wire _2128_;
	wire _2129_;
	wire _2130_;
	wire _2131_;
	wire _2132_;
	wire _2133_;
	wire _2134_;
	wire _2135_;
	wire _2136_;
	wire _2137_;
	wire _2138_;
	wire _2139_;
	wire _2140_;
	wire _2141_;
	wire _2142_;
	wire _2143_;
	wire _2144_;
	wire _2145_;
	wire _2146_;
	wire _2147_;
	wire _2148_;
	wire _2149_;
	wire _2150_;
	wire _2151_;
	wire _2152_;
	wire _2153_;
	wire _2154_;
	wire _2155_;
	wire _2156_;
	wire _2157_;
	wire _2158_;
	wire _2159_;
	wire _2160_;
	wire _2161_;
	wire _2162_;
	wire _2163_;
	wire _2164_;
	wire _2165_;
	wire _2166_;
	wire _2167_;
	wire _2168_;
	wire _2169_;
	wire _2170_;
	wire _2171_;
	wire _2172_;
	wire _2173_;
	wire _2174_;
	wire _2175_;
	wire _2176_;
	wire _2177_;
	wire _2178_;
	wire _2179_;
	wire _2180_;
	wire _2181_;
	wire _2182_;
	wire _2183_;
	wire _2184_;
	wire _2185_;
	wire _2186_;
	wire _2187_;
	wire _2188_;
	wire _2189_;
	wire _2190_;
	wire _2191_;
	wire _2192_;
	wire _2193_;
	wire _2194_;
	wire _2195_;
	wire _2196_;
	wire _2197_;
	wire _2198_;
	wire _2199_;
	wire _2200_;
	wire _2201_;
	wire _2202_;
	wire _2203_;
	wire _2204_;
	wire _2205_;
	wire _2206_;
	wire _2207_;
	wire _2208_;
	wire _2209_;
	wire _2210_;
	wire _2211_;
	wire _2212_;
	wire _2213_;
	wire _2214_;
	wire _2215_;
	wire _2216_;
	wire _2217_;
	wire _2218_;
	wire _2219_;
	wire _2220_;
	wire _2221_;
	wire _2222_;
	wire _2223_;
	wire _2224_;
	wire _2225_;
	wire _2226_;
	wire _2227_;
	wire _2228_;
	wire _2229_;
	wire _2230_;
	wire _2231_;
	wire _2232_;
	wire _2233_;
	wire _2234_;
	wire _2235_;
	wire _2236_;
	wire _2237_;
	wire _2238_;
	wire _2239_;
	wire _2240_;
	wire _2241_;
	wire _2242_;
	wire _2243_;
	wire _2244_;
	wire _2245_;
	wire _2246_;
	wire _2247_;
	wire _2248_;
	wire _2249_;
	wire _2250_;
	wire _2251_;
	wire _2252_;
	wire _2253_;
	wire _2254_;
	wire _2255_;
	wire _2256_;
	wire _2257_;
	wire _2258_;
	wire _2259_;
	wire _2260_;
	wire _2261_;
	wire _2262_;
	wire _2263_;
	wire _2264_;
	wire _2265_;
	wire _2266_;
	wire _2267_;
	wire _2268_;
	wire _2269_;
	wire _2270_;
	wire _2271_;
	wire _2272_;
	wire _2273_;
	wire _2274_;
	wire _2275_;
	wire _2276_;
	wire _2277_;
	wire _2278_;
	wire _2279_;
	wire _2280_;
	wire _2281_;
	wire _2282_;
	wire _2283_;
	wire _2284_;
	wire _2285_;
	wire _2286_;
	wire _2287_;
	wire _2288_;
	wire _2289_;
	wire _2290_;
	wire _2291_;
	wire _2292_;
	wire _2293_;
	wire _2294_;
	wire _2295_;
	wire _2296_;
	wire _2297_;
	wire _2298_;
	wire _2299_;
	wire _2300_;
	wire _2301_;
	wire _2302_;
	wire _2303_;
	wire _2304_;
	wire _2305_;
	wire _2306_;
	wire _2307_;
	wire _2308_;
	wire _2309_;
	wire _2310_;
	wire _2311_;
	wire _2312_;
	wire _2313_;
	wire _2314_;
	wire _2315_;
	wire _2316_;
	wire _2317_;
	wire _2318_;
	wire _2319_;
	wire _2320_;
	wire _2321_;
	wire _2322_;
	wire _2323_;
	wire _2324_;
	wire _2325_;
	wire _2326_;
	wire _2327_;
	wire _2328_;
	wire _2329_;
	wire _2330_;
	wire _2331_;
	wire _2332_;
	wire _2333_;
	wire _2334_;
	wire _2335_;
	wire _2336_;
	wire _2337_;
	wire _2338_;
	wire _2339_;
	wire _2340_;
	wire _2341_;
	wire _2342_;
	wire _2343_;
	wire _2344_;
	wire _2345_;
	wire _2346_;
	wire _2347_;
	wire _2348_;
	wire _2349_;
	wire _2350_;
	wire _2351_;
	wire _2352_;
	wire _2353_;
	wire _2354_;
	wire _2355_;
	wire _2356_;
	wire _2357_;
	wire _2358_;
	wire _2359_;
	wire _2360_;
	wire _2361_;
	wire _2362_;
	wire _2363_;
	wire _2364_;
	wire _2365_;
	wire _2366_;
	wire _2367_;
	wire _2368_;
	wire _2369_;
	wire _2370_;
	wire _2371_;
	wire _2372_;
	wire _2373_;
	wire _2374_;
	wire _2375_;
	wire _2376_;
	wire _2377_;
	wire _2378_;
	wire _2379_;
	wire _2380_;
	wire _2381_;
	wire _2382_;
	wire _2383_;
	wire _2384_;
	wire _2385_;
	wire _2386_;
	wire _2387_;
	wire _2388_;
	wire _2389_;
	wire _2390_;
	wire _2391_;
	wire _2392_;
	wire _2393_;
	wire _2394_;
	wire _2395_;
	wire _2396_;
	wire _2397_;
	wire _2398_;
	wire _2399_;
	wire _2400_;
	wire _2401_;
	wire _2402_;
	wire _2403_;
	wire _2404_;
	wire _2405_;
	wire _2406_;
	wire _2407_;
	wire _2408_;
	wire _2409_;
	wire _2410_;
	wire _2411_;
	wire _2412_;
	wire _2413_;
	wire _2414_;
	wire _2415_;
	wire _2416_;
	wire _2417_;
	wire _2418_;
	wire _2419_;
	wire _2420_;
	wire _2421_;
	wire _2422_;
	wire _2423_;
	wire _2424_;
	wire _2425_;
	wire _2426_;
	wire _2427_;
	wire _2428_;
	wire _2429_;
	wire _2430_;
	wire _2431_;
	wire _2432_;
	wire _2433_;
	wire _2434_;
	wire _2435_;
	wire _2436_;
	wire _2437_;
	wire _2438_;
	wire _2439_;
	wire _2440_;
	wire _2441_;
	wire _2442_;
	wire _2443_;
	wire _2444_;
	wire _2445_;
	wire _2446_;
	wire _2447_;
	wire _2448_;
	wire _2449_;
	wire _2450_;
	wire _2451_;
	wire _2452_;
	wire _2453_;
	wire _2454_;
	wire _2455_;
	wire _2456_;
	wire _2457_;
	wire _2458_;
	wire _2459_;
	wire _2460_;
	wire _2461_;
	wire _2462_;
	wire _2463_;
	wire _2464_;
	wire _2465_;
	wire _2466_;
	wire _2467_;
	wire _2468_;
	wire _2469_;
	wire _2470_;
	wire _2471_;
	wire _2472_;
	wire _2473_;
	wire _2474_;
	wire _2475_;
	wire _2476_;
	wire _2477_;
	wire _2478_;
	wire _2479_;
	wire _2480_;
	wire _2481_;
	wire _2482_;
	wire _2483_;
	wire _2484_;
	wire _2485_;
	wire _2486_;
	wire _2487_;
	wire _2488_;
	wire _2489_;
	wire _2490_;
	wire _2491_;
	wire _2492_;
	wire _2493_;
	wire _2494_;
	wire _2495_;
	wire _2496_;
	wire _2497_;
	wire _2498_;
	wire _2499_;
	wire _2500_;
	wire _2501_;
	wire _2502_;
	wire _2503_;
	wire _2504_;
	wire _2505_;
	wire _2506_;
	wire _2507_;
	wire _2508_;
	wire _2509_;
	wire _2510_;
	wire _2511_;
	wire _2512_;
	wire _2513_;
	wire _2514_;
	wire _2515_;
	wire _2516_;
	wire _2517_;
	wire _2518_;
	wire _2519_;
	wire _2520_;
	wire _2521_;
	wire _2522_;
	wire _2523_;
	wire _2524_;
	wire _2525_;
	wire _2526_;
	wire _2527_;
	wire _2528_;
	wire _2529_;
	wire _2530_;
	wire _2531_;
	wire _2532_;
	wire _2533_;
	wire _2534_;
	wire _2535_;
	wire _2536_;
	wire _2537_;
	wire _2538_;
	wire _2539_;
	wire _2540_;
	wire _2541_;
	wire _2542_;
	wire _2543_;
	wire _2544_;
	wire _2545_;
	wire _2546_;
	wire _2547_;
	wire _2548_;
	wire _2549_;
	wire _2550_;
	wire _2551_;
	wire _2552_;
	wire _2553_;
	wire _2554_;
	wire _2555_;
	wire _2556_;
	wire _2557_;
	wire _2558_;
	wire _2559_;
	wire _2560_;
	wire _2561_;
	wire _2562_;
	wire _2563_;
	wire _2564_;
	wire _2565_;
	wire _2566_;
	wire _2567_;
	wire _2568_;
	wire _2569_;
	wire _2570_;
	wire _2571_;
	wire _2572_;
	wire _2573_;
	wire _2574_;
	wire _2575_;
	wire _2576_;
	wire _2577_;
	wire _2578_;
	wire _2579_;
	wire _2580_;
	wire _2581_;
	wire _2582_;
	wire _2583_;
	wire _2584_;
	wire _2585_;
	wire _2586_;
	wire _2587_;
	wire _2588_;
	wire _2589_;
	wire _2590_;
	wire _2591_;
	wire _2592_;
	wire _2593_;
	wire _2594_;
	wire _2595_;
	wire _2596_;
	wire _2597_;
	wire _2598_;
	wire _2599_;
	wire _2600_;
	wire _2601_;
	wire _2602_;
	wire _2603_;
	wire _2604_;
	wire _2605_;
	wire _2606_;
	wire _2607_;
	wire _2608_;
	wire _2609_;
	wire _2610_;
	wire _2611_;
	wire _2612_;
	wire _2613_;
	wire _2614_;
	wire _2615_;
	wire _2616_;
	wire _2617_;
	wire _2618_;
	wire _2619_;
	wire _2620_;
	wire _2621_;
	wire _2622_;
	wire _2623_;
	wire _2624_;
	wire _2625_;
	wire _2626_;
	wire _2627_;
	wire _2628_;
	wire _2629_;
	wire _2630_;
	wire _2631_;
	wire _2632_;
	wire _2633_;
	wire _2634_;
	wire _2635_;
	wire _2636_;
	wire _2637_;
	wire _2638_;
	wire _2639_;
	wire _2640_;
	wire _2641_;
	wire _2642_;
	wire _2643_;
	wire _2644_;
	wire _2645_;
	wire _2646_;
	wire _2647_;
	wire _2648_;
	wire _2649_;
	wire _2650_;
	wire _2651_;
	wire _2652_;
	wire _2653_;
	wire _2654_;
	wire _2655_;
	wire _2656_;
	wire _2657_;
	wire _2658_;
	wire _2659_;
	wire _2660_;
	wire _2661_;
	wire _2662_;
	wire _2663_;
	wire _2664_;
	wire _2665_;
	wire _2666_;
	wire _2667_;
	wire _2668_;
	wire _2669_;
	wire _2670_;
	wire _2671_;
	wire _2672_;
	wire _2673_;
	wire _2674_;
	wire _2675_;
	wire _2676_;
	wire _2677_;
	wire _2678_;
	wire _2679_;
	wire _2680_;
	wire _2681_;
	wire _2682_;
	wire _2683_;
	wire _2684_;
	wire _2685_;
	wire _2686_;
	wire _2687_;
	wire _2688_;
	wire _2689_;
	wire _2690_;
	wire _2691_;
	wire _2692_;
	wire _2693_;
	wire _2694_;
	wire _2695_;
	wire _2696_;
	wire _2697_;
	wire _2698_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	reg [11:0] \mchip.index ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire [7:0] \mchip.val ;
	assign _1097_ = \mchip.index [0] | ~\mchip.index [2];
	assign _1208_ = \mchip.index [5] & ~_1097_;
	assign _1319_ = ~\mchip.index [9];
	assign _1430_ = ~\mchip.index [7];
	assign _1540_ = ~\mchip.index [6];
	assign _1651_ = ~(\mchip.index [0] & \mchip.index [2]);
	assign _1762_ = _1651_ | \mchip.index [3];
	assign _1873_ = _1762_ | _1540_;
	assign _1909_ = _1873_ | _1430_;
	assign _1920_ = _1319_ & ~_1909_;
	assign _1931_ = ~\mchip.index [10];
	assign _1942_ = \mchip.index [2] | ~\mchip.index [1];
	assign _1953_ = _1942_ | \mchip.index [7];
	assign _1964_ = _1953_ | _1319_;
	assign _1975_ = _1931_ & ~_1964_;
	assign _1986_ = \mchip.index [1] | ~\mchip.index [2];
	assign _1997_ = _1986_ | \mchip.index [3];
	assign _2008_ = _1997_ | \mchip.index [8];
	assign _2019_ = \mchip.index [9] & ~_2008_;
	assign _2030_ = ~\mchip.index [4];
	assign _2041_ = _1762_ | _2030_;
	assign _2052_ = _2041_ | \mchip.index [6];
	assign _2063_ = \mchip.index [9] & ~_2052_;
	assign _2074_ = _1986_ | \mchip.index [4];
	assign _2085_ = _2074_ | \mchip.index [6];
	assign _2096_ = \mchip.index [7] & ~_2085_;
	assign _2107_ = _2096_ & ~\mchip.index [10];
	assign _2118_ = \mchip.index [0] | ~\mchip.index [5];
	assign _2129_ = _2118_ | \mchip.index [6];
	assign _2139_ = _2129_ | _1430_;
	assign _2150_ = \mchip.index [8] & ~_2139_;
	assign _2161_ = ~\mchip.index [5];
	assign _2172_ = \mchip.index [4] | ~\mchip.index [1];
	assign _2183_ = _2172_ | _2161_;
	assign _2194_ = _2183_ | _1430_;
	assign _2205_ = \mchip.index [8] & ~_2194_;
	assign _2216_ = _1651_ | \mchip.index [4];
	assign _2227_ = _2216_ | \mchip.index [5];
	assign _2238_ = _2227_ | \mchip.index [7];
	assign _2249_ = _2238_ | _1319_;
	assign _2260_ = _1931_ & ~_2249_;
	assign _2271_ = ~\mchip.index [11];
	assign _2282_ = \mchip.index [1] | ~\mchip.index [5];
	assign _2293_ = _2282_ | _1540_;
	assign _2304_ = _2271_ & ~_2293_;
	assign _2315_ = ~(\mchip.index [3] & \mchip.index [2]);
	assign _2326_ = _2315_ | \mchip.index [6];
	assign _2337_ = _2326_ | \mchip.index [8];
	assign _2348_ = \mchip.index [10] & ~_2337_;
	assign _2359_ = ~\mchip.index [8];
	assign _2370_ = \mchip.index [3] | ~\mchip.index [0];
	assign _2381_ = _2370_ | _2030_;
	assign _2392_ = _2381_ | \mchip.index [5];
	assign _2403_ = _2392_ | \mchip.index [7];
	assign _2414_ = _2403_ | _2359_;
	assign _2425_ = \mchip.index [10] & ~_2414_;
	assign _2436_ = \mchip.index [3] | ~\mchip.index [1];
	assign _2446_ = _2436_ | _2030_;
	assign _2457_ = _2446_ | _1540_;
	assign _2468_ = _2457_ | \mchip.index [8];
	assign _2479_ = \mchip.index [10] & ~_2468_;
	assign _2490_ = \mchip.index [0] | \mchip.index [2];
	assign _2501_ = _2490_ | \mchip.index [3];
	assign _2512_ = _2501_ | \mchip.index [4];
	assign _2523_ = _2512_ | _1430_;
	assign _2534_ = _2523_ | _1319_;
	assign _2545_ = _2534_ | \mchip.index [10];
	assign _2556_ = _2271_ & ~_2545_;
	assign _2567_ = ~\mchip.index [3];
	assign _2578_ = ~\mchip.index [2];
	assign _2589_ = \mchip.index [0] | ~\mchip.index [1];
	assign _2600_ = _2589_ | _2578_;
	assign _2611_ = _2600_ | _2567_;
	assign _2622_ = _2611_ | \mchip.index [4];
	assign _2633_ = _1430_ & ~_2622_;
	assign _2644_ = _1986_ | _2030_;
	assign _2655_ = _2644_ | _1540_;
	assign _2666_ = _2655_ | \mchip.index [7];
	assign _2677_ = _1319_ & ~_2666_;
	assign _2688_ = \mchip.index [1] | ~\mchip.index [0];
	assign _0000_ = _2688_ | _2578_;
	assign _0011_ = _0000_ | _2567_;
	assign _0022_ = _0011_ | _1540_;
	assign _0033_ = _0022_ | \mchip.index [7];
	assign _0044_ = ~(\mchip.index [1] & \mchip.index [0]);
	assign _0055_ = _0044_ | _2578_;
	assign _0066_ = _0055_ | _1931_;
	assign _0077_ = _2271_ & ~_0066_;
	assign _0088_ = _1942_ | \mchip.index [3];
	assign _0099_ = _0088_ | \mchip.index [4];
	assign _0110_ = _0099_ | \mchip.index [7];
	assign _0121_ = _1931_ & ~_0110_;
	assign _0132_ = _0088_ | \mchip.index [5];
	assign _0143_ = _0132_ | \mchip.index [6];
	assign _0154_ = \mchip.index [9] & ~_0143_;
	assign _0165_ = \mchip.index [1] | \mchip.index [0];
	assign _0176_ = _0165_ | \mchip.index [2];
	assign _0187_ = _0176_ | _2567_;
	assign _0198_ = _0187_ | \mchip.index [4];
	assign _0208_ = _1430_ & ~_0198_;
	assign _0219_ = _1097_ | _1540_;
	assign _0230_ = _0219_ | \mchip.index [8];
	assign _0241_ = _1931_ & ~_0230_;
	assign _0252_ = \mchip.index [3] | \mchip.index [2];
	assign _0263_ = _0252_ | _1540_;
	assign _0274_ = _0263_ | \mchip.index [7];
	assign _0285_ = _0274_ | \mchip.index [8];
	assign _0296_ = _0285_ | \mchip.index [9];
	assign _0307_ = _0296_ | _1931_;
	assign _0318_ = _2271_ & ~_0307_;
	assign _0329_ = _0165_ | \mchip.index [3];
	assign _0340_ = _0329_ | _2030_;
	assign _0351_ = _0340_ | _1540_;
	assign _0362_ = _0351_ | \mchip.index [7];
	assign _0373_ = _1319_ & ~_0362_;
	assign _0384_ = _1762_ | \mchip.index [5];
	assign _0395_ = _0384_ | \mchip.index [6];
	assign _0406_ = _0395_ | _2359_;
	assign _0417_ = _2271_ & ~_0406_;
	assign _0428_ = \mchip.index [2] | ~\mchip.index [0];
	assign _0439_ = _0428_ | \mchip.index [4];
	assign _0450_ = _0439_ | _2161_;
	assign _0461_ = _1430_ & ~_0450_;
	assign _0472_ = _2589_ | \mchip.index [3];
	assign _0483_ = _0472_ | \mchip.index [6];
	assign _0494_ = _0483_ | \mchip.index [7];
	assign _0505_ = \mchip.index [9] & ~_0494_;
	assign _0516_ = _2490_ | _2030_;
	assign _0527_ = _0516_ | _1540_;
	assign _0538_ = _0527_ | _1430_;
	assign _0549_ = _2359_ & ~_0538_;
	assign _0560_ = _2446_ | \mchip.index [5];
	assign _0571_ = _0560_ | \mchip.index [6];
	assign _0582_ = \mchip.index [8] & ~_0571_;
	assign _0593_ = _0055_ | \mchip.index [3];
	assign _0604_ = _0593_ | \mchip.index [4];
	assign _0615_ = _0604_ | \mchip.index [5];
	assign _0626_ = _0615_ | _1540_;
	assign _0637_ = \mchip.index [9] & ~_0626_;
	assign _0648_ = _0472_ | \mchip.index [4];
	assign _0659_ = _0648_ | _1540_;
	assign _0669_ = _0659_ | _1430_;
	assign _0680_ = \mchip.index [9] & ~_0669_;
	assign _0691_ = _2370_ | \mchip.index [4];
	assign _0702_ = _0691_ | \mchip.index [6];
	assign _0713_ = _0702_ | \mchip.index [7];
	assign _0724_ = _2359_ & ~_0713_;
	assign _0735_ = _0648_ | \mchip.index [8];
	assign _0746_ = \mchip.index [9] & ~_0735_;
	assign _0757_ = ~(\mchip.index [2] & \mchip.index [4]);
	assign _0768_ = _0757_ | \mchip.index [6];
	assign _0779_ = _0768_ | _1430_;
	assign _0790_ = _0779_ | \mchip.index [8];
	assign _0801_ = \mchip.index [10] & ~_0790_;
	assign _0812_ = _0252_ | \mchip.index [4];
	assign _0823_ = _0812_ | _1540_;
	assign _0834_ = _0823_ | \mchip.index [7];
	assign _0845_ = _0834_ | _2359_;
	assign _0856_ = _0845_ | \mchip.index [10];
	assign _0867_ = _2271_ & ~_0856_;
	assign _0878_ = _0165_ | _2578_;
	assign _0889_ = _0878_ | _2567_;
	assign _0900_ = _0889_ | \mchip.index [6];
	assign _0911_ = \mchip.index [7] & ~_0900_;
	assign _0922_ = _0472_ | _2161_;
	assign _0933_ = \mchip.index [9] & ~_0922_;
	assign _0944_ = _1097_ | \mchip.index [3];
	assign _0955_ = _0944_ | _2030_;
	assign _0966_ = _0955_ | _1540_;
	assign _0977_ = _1931_ & ~_0966_;
	assign _0988_ = \mchip.index [2] | ~\mchip.index [4];
	assign _0999_ = _0988_ | _1430_;
	assign _1010_ = _0999_ | \mchip.index [9];
	assign _1021_ = _1931_ & ~_1010_;
	assign _1032_ = \mchip.index [1] | \mchip.index [2];
	assign _1043_ = _1032_ | _2567_;
	assign _1054_ = _1043_ | _1540_;
	assign _1065_ = _1054_ | _1430_;
	assign _1076_ = _2271_ & ~_1065_;
	assign _1087_ = ~(\mchip.index [0] & \mchip.index [3]);
	assign _1098_ = _1087_ | _2030_;
	assign _1109_ = _1098_ | \mchip.index [7];
	assign _1120_ = _2271_ & ~_1109_;
	assign _1131_ = _0252_ | _2030_;
	assign _1142_ = _1131_ | \mchip.index [5];
	assign _1153_ = _1142_ | _1540_;
	assign _1164_ = _1153_ | \mchip.index [7];
	assign _1175_ = \mchip.index [10] & ~_1164_;
	assign _1186_ = _2688_ | _2567_;
	assign _1197_ = _1186_ | \mchip.index [9];
	assign _1209_ = _1931_ & ~_1197_;
	assign _1220_ = _0516_ | \mchip.index [6];
	assign _1231_ = _1220_ | _1430_;
	assign _1242_ = \mchip.index [9] & ~_1231_;
	assign _1253_ = _1651_ | _2030_;
	assign _1264_ = _1253_ | _1430_;
	assign _1275_ = _1264_ | _2359_;
	assign _1286_ = _1931_ & ~_1275_;
	assign _1297_ = \mchip.index [2] | ~\mchip.index [3];
	assign _1308_ = _1297_ | \mchip.index [4];
	assign _1320_ = _1308_ | _1430_;
	assign _1331_ = _1319_ & ~_1320_;
	assign _1342_ = _0044_ | _2567_;
	assign _1353_ = _1342_ | \mchip.index [8];
	assign _1364_ = \mchip.index [9] & ~_1353_;
	assign _1375_ = _0044_ | \mchip.index [2];
	assign _1386_ = _1375_ | \mchip.index [3];
	assign _1397_ = _1386_ | \mchip.index [7];
	assign _1408_ = _2271_ & ~_1397_;
	assign _1419_ = _0428_ | \mchip.index [3];
	assign _1431_ = _1419_ | \mchip.index [4];
	assign _1442_ = _1431_ | \mchip.index [6];
	assign _1453_ = \mchip.index [9] & ~_1442_;
	assign _1464_ = _2688_ | _2030_;
	assign _1474_ = _1464_ | _1540_;
	assign _1485_ = _1474_ | _1430_;
	assign _1496_ = _1931_ & ~_1485_;
	assign _1507_ = _2589_ | \mchip.index [2];
	assign _1518_ = _1507_ | _2030_;
	assign _1529_ = _1518_ | _1430_;
	assign _1541_ = _2271_ & ~_1529_;
	assign _1552_ = _0878_ | \mchip.index [4];
	assign _1563_ = _1552_ | \mchip.index [6];
	assign _1574_ = \mchip.index [10] & ~_1563_;
	assign _1585_ = _1953_ | \mchip.index [8];
	assign _1596_ = \mchip.index [10] & ~_1585_;
	assign _1607_ = \mchip.index [1] | \mchip.index [3];
	assign _1618_ = _1607_ | \mchip.index [4];
	assign _1629_ = _1618_ | \mchip.index [5];
	assign _1640_ = _1629_ | _1430_;
	assign _1652_ = _1640_ | _2359_;
	assign _1663_ = _1652_ | _1319_;
	assign _1674_ = _1663_ | _1931_;
	assign _1685_ = \mchip.index [11] & ~_1674_;
	assign _1696_ = \mchip.index [0] | \mchip.index [3];
	assign _1707_ = _1696_ | _2030_;
	assign _1718_ = _1707_ | \mchip.index [7];
	assign _1729_ = _1718_ | \mchip.index [8];
	assign _1740_ = \mchip.index [10] & ~_1729_;
	assign _1751_ = _2688_ | \mchip.index [4];
	assign _1763_ = _1751_ | _1540_;
	assign _1774_ = _1763_ | _2359_;
	assign _1785_ = _1319_ & ~_1774_;
	assign _1796_ = _0044_ | \mchip.index [4];
	assign _1807_ = _1796_ | \mchip.index [6];
	assign _1818_ = _1807_ | _1430_;
	assign _1829_ = \mchip.index [8] & ~_1818_;
	assign _1840_ = \mchip.index [7] & ~_1552_;
	assign _1851_ = _1651_ | _2567_;
	assign _1862_ = _1851_ | \mchip.index [7];
	assign _1874_ = _1931_ & ~_1862_;
	assign _1885_ = _2315_ | _2030_;
	assign _1896_ = _1885_ | _1430_;
	assign _1902_ = _1319_ & ~_1896_;
	assign _1903_ = \mchip.index [1] | ~\mchip.index [3];
	assign _1904_ = _1903_ | _2030_;
	assign _1905_ = _1904_ | _1540_;
	assign _1906_ = _1905_ | \mchip.index [7];
	assign _1907_ = \mchip.index [11] & ~_1906_;
	assign _1908_ = _1342_ | \mchip.index [6];
	assign _1910_ = _1908_ | _1430_;
	assign _1911_ = \mchip.index [10] & ~_1910_;
	assign _1912_ = _0944_ | _1540_;
	assign _1913_ = _1912_ | \mchip.index [7];
	assign _1914_ = _1319_ & ~_1913_;
	assign _1915_ = _2490_ | \mchip.index [4];
	assign _1916_ = _1915_ | _2359_;
	assign _1917_ = _1916_ | _1319_;
	assign _1918_ = _1917_ | \mchip.index [10];
	assign _1919_ = _2271_ & ~_1918_;
	assign _1921_ = _1931_ & ~_1220_;
	assign _1922_ = ~(\mchip.index [5] & \mchip.index [3]);
	assign _1923_ = \mchip.index [7] & ~_1922_;
	assign _1924_ = _1308_ | _1540_;
	assign _1925_ = _1924_ | _1430_;
	assign _1926_ = \mchip.index [10] & ~_1925_;
	assign _1927_ = _1942_ | _2567_;
	assign _1928_ = _1927_ | \mchip.index [6];
	assign _1929_ = _2359_ & ~_1928_;
	assign _1930_ = _2490_ | _2567_;
	assign _1932_ = _1930_ | \mchip.index [5];
	assign _1933_ = _1932_ | \mchip.index [7];
	assign _1934_ = \mchip.index [9] & ~_1933_;
	assign _1935_ = _0428_ | _2567_;
	assign _1936_ = _1935_ | \mchip.index [4];
	assign _1937_ = _1936_ | _2359_;
	assign _1938_ = \mchip.index [10] & ~_1937_;
	assign _1939_ = _1419_ | _2030_;
	assign _1940_ = _1939_ | _1540_;
	assign _1941_ = _1940_ | \mchip.index [7];
	assign _1943_ = \mchip.index [9] & ~_1941_;
	assign _1944_ = _1903_ | _1430_;
	assign _1945_ = _1944_ | _2359_;
	assign _1946_ = _1931_ & ~_1945_;
	assign _1947_ = _1043_ | _2030_;
	assign _1948_ = _1947_ | \mchip.index [6];
	assign _1949_ = \mchip.index [9] & ~_1948_;
	assign _1950_ = \mchip.index [0] | ~\mchip.index [3];
	assign _1951_ = _1950_ | _1430_;
	assign _1952_ = _1951_ | \mchip.index [9];
	assign _1954_ = \mchip.index [10] & ~_1952_;
	assign _1955_ = _1431_ | _2359_;
	assign _1956_ = _1931_ & ~_1955_;
	assign _1957_ = ~(\mchip.index [1] & \mchip.index [2]);
	assign _1958_ = _1957_ | _2567_;
	assign _1959_ = _1958_ | \mchip.index [4];
	assign _1960_ = _1959_ | _2359_;
	assign _1961_ = _2271_ & ~_1960_;
	assign _1962_ = \mchip.index [2] | \mchip.index [4];
	assign _1963_ = _1962_ | \mchip.index [5];
	assign _1965_ = _1963_ | \mchip.index [6];
	assign _1966_ = _1965_ | _1430_;
	assign _1967_ = _1966_ | \mchip.index [8];
	assign _1968_ = _1967_ | \mchip.index [9];
	assign _1969_ = _1968_ | _1931_;
	assign _1970_ = _2271_ & ~_1969_;
	assign _1971_ = _2074_ | _2161_;
	assign _1972_ = _1971_ | \mchip.index [7];
	assign _1973_ = \mchip.index [11] & ~_1972_;
	assign _1974_ = _2688_ | \mchip.index [2];
	assign _1976_ = _1974_ | \mchip.index [3];
	assign _1977_ = _1540_ & ~_1976_;
	assign _1978_ = ~(_1977_ & \mchip.index [7]);
	assign _1979_ = \mchip.index [10] & ~_1978_;
	assign _1980_ = _0000_ | \mchip.index [3];
	assign _1981_ = _1980_ | \mchip.index [5];
	assign _1982_ = _1981_ | \mchip.index [6];
	assign _1983_ = \mchip.index [9] & ~_1982_;
	assign _1984_ = _0165_ | \mchip.index [4];
	assign _1985_ = _1984_ | \mchip.index [5];
	assign _1987_ = _1985_ | \mchip.index [6];
	assign _1988_ = _1987_ | _2359_;
	assign _1989_ = _1988_ | _1319_;
	assign _1990_ = _1989_ | _1931_;
	assign _1991_ = \mchip.index [11] & ~_1990_;
	assign _1992_ = _2501_ | \mchip.index [7];
	assign _1993_ = _1992_ | \mchip.index [8];
	assign _1994_ = _1993_ | \mchip.index [9];
	assign _1995_ = _1994_ | _1931_;
	assign _1996_ = _2271_ & ~_1995_;
	assign _1998_ = _1942_ | \mchip.index [4];
	assign _1999_ = _1998_ | \mchip.index [7];
	assign _2000_ = _1999_ | _2359_;
	assign _2001_ = _1931_ & ~_2000_;
	assign _2002_ = _1957_ | _2030_;
	assign _2003_ = _2002_ | _1540_;
	assign _2004_ = _2003_ | \mchip.index [7];
	assign _2005_ = \mchip.index [11] & ~_2004_;
	assign _2006_ = _1032_ | _2030_;
	assign _2007_ = _2006_ | _2359_;
	assign _2009_ = _2007_ | \mchip.index [9];
	assign _2010_ = \mchip.index [10] & ~_2009_;
	assign _2011_ = \mchip.index [1] | ~\mchip.index [4];
	assign _2012_ = _2011_ | _2161_;
	assign _2013_ = _1540_ & ~_2012_;
	assign _2014_ = _0878_ | _1540_;
	assign _2015_ = _2014_ | _1319_;
	assign _2016_ = _2271_ & ~_2015_;
	assign _2017_ = _1957_ | \mchip.index [6];
	assign _2018_ = _2017_ | _1430_;
	assign _2020_ = _2018_ | _1931_;
	assign _2021_ = _2271_ & ~_2020_;
	assign _2022_ = _1904_ | _2359_;
	assign _2023_ = _2022_ | _1319_;
	assign _2024_ = _2271_ & ~_2023_;
	assign _2025_ = _0044_ | \mchip.index [3];
	assign _2026_ = _2025_ | \mchip.index [4];
	assign _2027_ = _2026_ | \mchip.index [8];
	assign _2028_ = _1319_ & ~_2027_;
	assign _2029_ = _1087_ | \mchip.index [4];
	assign _2031_ = _2029_ | \mchip.index [6];
	assign _2032_ = _2031_ | \mchip.index [7];
	assign _2033_ = \mchip.index [11] & ~_2032_;
	assign _2034_ = _2033_ | _2028_;
	assign _2035_ = _2034_ | _2024_;
	assign _2036_ = _2035_ | _2021_;
	assign _2037_ = _2036_ | _2016_;
	assign _2038_ = _2037_ | _2013_;
	assign _2039_ = _2038_ | _2010_;
	assign _2040_ = _2039_ | _2005_;
	assign _2042_ = _2040_ | _2001_;
	assign _2043_ = _2042_ | _1996_;
	assign _2044_ = _2043_ | _1991_;
	assign _2045_ = _2044_ | _1983_;
	assign _2046_ = _2045_ | _1979_;
	assign _2047_ = _2046_ | _1973_;
	assign _2048_ = _2047_ | _1970_;
	assign _2049_ = _2048_ | _1961_;
	assign _2050_ = _2049_ | _1956_;
	assign _2051_ = _2050_ | _1954_;
	assign _2053_ = _2051_ | _1949_;
	assign _2054_ = _2053_ | _1946_;
	assign _2055_ = _2054_ | _1943_;
	assign _2056_ = _2055_ | _1938_;
	assign _2057_ = _2056_ | _1934_;
	assign _2058_ = _2057_ | _1929_;
	assign _2059_ = _2058_ | _1926_;
	assign _2060_ = _2059_ | _1923_;
	assign _2061_ = _2060_ | _1921_;
	assign _2062_ = _2061_ | _1919_;
	assign _2064_ = _2062_ | _1914_;
	assign _2065_ = _2064_ | _1911_;
	assign _2066_ = _2065_ | _1907_;
	assign _2067_ = _2066_ | _1902_;
	assign _2068_ = _2067_ | _1874_;
	assign _2069_ = _2068_ | _1840_;
	assign _2070_ = _2069_ | _1829_;
	assign _2071_ = _2070_ | _1785_;
	assign _2072_ = _2071_ | _1740_;
	assign _2073_ = _2072_ | _1685_;
	assign _2075_ = _2073_ | _1596_;
	assign _2076_ = _2075_ | _1574_;
	assign _2077_ = _2076_ | _1541_;
	assign _2078_ = _2077_ | _1496_;
	assign _2079_ = _2078_ | _1453_;
	assign _2080_ = _2079_ | _1408_;
	assign _2081_ = _2080_ | _1364_;
	assign _2082_ = _2081_ | _1331_;
	assign _2083_ = _2082_ | _1286_;
	assign _2084_ = _2083_ | _1242_;
	assign _2086_ = _2084_ | _1209_;
	assign _2087_ = _2086_ | _1175_;
	assign _2088_ = _2087_ | _1120_;
	assign _2089_ = _2088_ | _1076_;
	assign _2090_ = _2089_ | _1021_;
	assign _2091_ = _2090_ | _0977_;
	assign _2092_ = _2091_ | _0933_;
	assign _2093_ = _2092_ | _0911_;
	assign _2094_ = _2093_ | _0867_;
	assign _2095_ = _2094_ | _0801_;
	assign _2097_ = _2095_ | _0746_;
	assign _2098_ = _2097_ | _0724_;
	assign _2099_ = _2098_ | _0680_;
	assign _2100_ = _2099_ | _0637_;
	assign _2101_ = _2100_ | _0582_;
	assign _2102_ = _2101_ | _0549_;
	assign _2103_ = _2102_ | _0505_;
	assign _2104_ = _2103_ | _0461_;
	assign _2105_ = _2104_ | _0417_;
	assign _2106_ = _2105_ | _0373_;
	assign _2108_ = _2106_ | _0318_;
	assign _2109_ = _2108_ | _0241_;
	assign _2110_ = _2109_ | _0208_;
	assign _2111_ = _2110_ | _0154_;
	assign _2112_ = _2111_ | _0121_;
	assign _2113_ = ~(_2112_ | _0077_);
	assign _2114_ = ~(_2113_ & _0033_);
	assign _2115_ = _2114_ | _2677_;
	assign _2116_ = _2115_ | _2633_;
	assign _2117_ = _2116_ | _2556_;
	assign _2119_ = _2117_ | _2479_;
	assign _2120_ = _2119_ | _2425_;
	assign _2121_ = _2120_ | _2348_;
	assign _2122_ = _2121_ | _2304_;
	assign _2123_ = _2122_ | _2260_;
	assign _2124_ = _2123_ | _2205_;
	assign _2125_ = _2124_ | _2150_;
	assign _2126_ = _2125_ | _2107_;
	assign _2127_ = _2126_ | _2063_;
	assign _2128_ = _2127_ | _2019_;
	assign _2130_ = _2128_ | _1975_;
	assign _2131_ = _2130_ | _1920_;
	assign \mchip.val [6] = _2131_ | _1208_;
	assign _2132_ = _1903_ | \mchip.index [4];
	assign _2133_ = _2132_ | _1430_;
	assign _2134_ = _2359_ & ~_2133_;
	assign _2135_ = \mchip.index [11] & ~_1951_;
	assign _2136_ = \mchip.index [4] | ~\mchip.index [0];
	assign _2137_ = _2136_ | \mchip.index [8];
	assign _2138_ = \mchip.index [9] & ~_2137_;
	assign _2140_ = _1931_ & ~_1935_;
	assign _2141_ = _1997_ | _1540_;
	assign _2142_ = _2141_ | \mchip.index [7];
	assign _2143_ = _1319_ & ~_2142_;
	assign _2144_ = \mchip.index [0] | \mchip.index [4];
	assign _2145_ = _2144_ | _2161_;
	assign _2146_ = _1430_ & ~_2145_;
	assign _2147_ = _1998_ | \mchip.index [6];
	assign _2148_ = _2147_ | _1430_;
	assign _2149_ = \mchip.index [10] & ~_2148_;
	assign _2151_ = \mchip.index [5] | ~\mchip.index [2];
	assign _2152_ = _2151_ | _1540_;
	assign _2153_ = _2152_ | _1430_;
	assign _2154_ = \mchip.index [11] & ~_2153_;
	assign _2155_ = \mchip.index [0] | ~\mchip.index [4];
	assign _2156_ = _2155_ | _1430_;
	assign _2157_ = \mchip.index [11] & ~_2156_;
	assign _2158_ = _1974_ | \mchip.index [4];
	assign _2159_ = _2359_ & ~_2158_;
	assign _2160_ = _2359_ & ~_1924_;
	assign _2162_ = ~(\mchip.index [0] & \mchip.index [4]);
	assign _2163_ = _2162_ | _1540_;
	assign _2164_ = _2163_ | _1430_;
	assign _2165_ = \mchip.index [8] & ~_2164_;
	assign _2166_ = _0088_ | _2030_;
	assign _2167_ = \mchip.index [6] & ~_2166_;
	assign _2168_ = _1297_ | _1540_;
	assign _2169_ = \mchip.index [7] & ~_2168_;
	assign _2170_ = _0088_ | \mchip.index [7];
	assign _2171_ = _2170_ | _2359_;
	assign _2173_ = \mchip.index [10] & ~_2171_;
	assign _2174_ = _1851_ | _2030_;
	assign _2175_ = \mchip.index [6] & ~_2174_;
	assign _2176_ = \mchip.index [8] & ~_0560_;
	assign _2177_ = \mchip.index [1] | \mchip.index [4];
	assign _2178_ = _2177_ | _1540_;
	assign _2179_ = _2178_ | _1430_;
	assign _2180_ = _2179_ | \mchip.index [8];
	assign _2181_ = _2180_ | \mchip.index [9];
	assign _2182_ = _2181_ | _1931_;
	assign _2184_ = _2271_ & ~_2182_;
	assign _2185_ = _1651_ | _2161_;
	assign _2186_ = _2185_ | \mchip.index [6];
	assign _2187_ = \mchip.index [10] & ~_2186_;
	assign _2188_ = _0428_ | _1540_;
	assign _2189_ = _2188_ | _1430_;
	assign _2190_ = _2271_ & ~_2189_;
	assign _2191_ = _0055_ | \mchip.index [7];
	assign _2192_ = _2359_ & ~_2191_;
	assign _2193_ = _1342_ | \mchip.index [4];
	assign _2195_ = _2193_ | \mchip.index [5];
	assign _2196_ = _1430_ & ~_2195_;
	assign _2197_ = _1319_ & ~_2337_;
	assign _2198_ = _2006_ | _1430_;
	assign _2199_ = \mchip.index [9] & ~_2198_;
	assign _2200_ = _2688_ | \mchip.index [3];
	assign _2201_ = _2200_ | \mchip.index [8];
	assign _2202_ = \mchip.index [9] & ~_2201_;
	assign _2203_ = \mchip.index [3] | ~\mchip.index [4];
	assign _2204_ = _2203_ | _1540_;
	assign _2206_ = _2204_ | \mchip.index [7];
	assign _2207_ = _1319_ & ~_2206_;
	assign _2208_ = _1186_ | _2030_;
	assign _2209_ = \mchip.index [8] & ~_2208_;
	assign _2210_ = _1540_ & ~_2006_;
	assign _2211_ = _1957_ | \mchip.index [4];
	assign _2212_ = _2211_ | \mchip.index [7];
	assign _2213_ = _2212_ | _2359_;
	assign _2214_ = _1931_ & ~_2213_;
	assign _2215_ = ~(\mchip.index [1] & \mchip.index [6]);
	assign _2217_ = _2215_ | _2359_;
	assign _2218_ = _1319_ & ~_2217_;
	assign _2219_ = _0944_ | \mchip.index [6];
	assign _2220_ = _1931_ & ~_2219_;
	assign _2221_ = \mchip.index [9] & ~_1043_;
	assign _2222_ = _1097_ | _2567_;
	assign _2223_ = _2222_ | \mchip.index [7];
	assign _2224_ = _2223_ | _2359_;
	assign _2225_ = _1931_ & ~_2224_;
	assign _2226_ = _1931_ & ~_1718_;
	assign _2228_ = _0560_ | _1430_;
	assign _2229_ = \mchip.index [10] & ~_2228_;
	assign _2230_ = _0165_ | _2567_;
	assign _2231_ = _2230_ | \mchip.index [6];
	assign _2232_ = _2359_ & ~_2231_;
	assign _2233_ = \mchip.index [6] | ~\mchip.index [0];
	assign _2234_ = _2233_ | _1430_;
	assign _2235_ = _2234_ | _1931_;
	assign _2236_ = _2271_ & ~_2235_;
	assign _2237_ = _1696_ | \mchip.index [6];
	assign _2239_ = _2237_ | \mchip.index [7];
	assign _2240_ = _2239_ | _2359_;
	assign _2241_ = _2240_ | \mchip.index [9];
	assign _2242_ = _2241_ | _1931_;
	assign _2243_ = _2271_ & ~_2242_;
	assign _2244_ = _0648_ | \mchip.index [6];
	assign _2245_ = _1430_ & ~_2244_;
	assign _2246_ = _1942_ | _1430_;
	assign _2247_ = _2246_ | _2359_;
	assign _2248_ = _1931_ & ~_2247_;
	assign _2250_ = _1998_ | \mchip.index [5];
	assign _2251_ = _2250_ | \mchip.index [6];
	assign _2252_ = \mchip.index [8] & ~_2251_;
	assign _2253_ = _0044_ | _2030_;
	assign _2254_ = _1319_ & ~_2253_;
	assign _2255_ = _2136_ | _1540_;
	assign _2256_ = _2255_ | \mchip.index [8];
	assign _2257_ = _1931_ & ~_2256_;
	assign _2258_ = _2370_ | _1540_;
	assign _2259_ = _2258_ | \mchip.index [7];
	assign _2261_ = _1319_ & ~_2259_;
	assign _2262_ = _1997_ | \mchip.index [4];
	assign _2263_ = _2262_ | \mchip.index [5];
	assign _2264_ = _2263_ | _1430_;
	assign _2265_ = \mchip.index [8] & ~_2264_;
	assign _2266_ = _0165_ | _2030_;
	assign _2267_ = _2266_ | \mchip.index [7];
	assign _2268_ = _2267_ | \mchip.index [9];
	assign _2269_ = \mchip.index [10] & ~_2268_;
	assign _2270_ = _0944_ | \mchip.index [5];
	assign _2272_ = _2270_ | _1540_;
	assign _2273_ = _2272_ | _1430_;
	assign _2274_ = \mchip.index [10] & ~_2273_;
	assign _2275_ = _2074_ | \mchip.index [7];
	assign _2276_ = _2275_ | _2359_;
	assign _2277_ = \mchip.index [10] & ~_2276_;
	assign _2278_ = _1931_ & ~_2193_;
	assign _2279_ = _1851_ | _1540_;
	assign _2280_ = \mchip.index [9] & ~_2279_;
	assign _2281_ = _2144_ | _1540_;
	assign _2283_ = _2281_ | \mchip.index [7];
	assign _2284_ = _2283_ | _2359_;
	assign _2285_ = _2284_ | _1319_;
	assign _2286_ = _2285_ | _1931_;
	assign _2287_ = \mchip.index [11] & ~_2286_;
	assign _2288_ = _1959_ | _1540_;
	assign _2289_ = _1430_ & ~_2288_;
	assign _2290_ = _2436_ | \mchip.index [6];
	assign _2291_ = _2290_ | \mchip.index [7];
	assign _2292_ = \mchip.index [9] & ~_2291_;
	assign _2294_ = _1942_ | \mchip.index [5];
	assign _2295_ = _2294_ | _1540_;
	assign _2296_ = _2295_ | _1931_;
	assign _2297_ = _2271_ & ~_2296_;
	assign _2298_ = _0889_ | \mchip.index [4];
	assign _2299_ = \mchip.index [10] & ~_2298_;
	assign _2300_ = _0099_ | \mchip.index [6];
	assign _2301_ = \mchip.index [9] & ~_2300_;
	assign _2302_ = _1375_ | \mchip.index [5];
	assign _2303_ = _2302_ | _1430_;
	assign _2305_ = \mchip.index [9] & ~_2303_;
	assign _2306_ = _2270_ | _2359_;
	assign _2307_ = \mchip.index [10] & ~_2306_;
	assign _2308_ = \mchip.index [8] & ~_2288_;
	assign _2309_ = ~(\mchip.index [1] & \mchip.index [4]);
	assign _2310_ = _2309_ | _1540_;
	assign _2311_ = _2310_ | _1430_;
	assign _2312_ = \mchip.index [10] & ~_2311_;
	assign _2313_ = _1032_ | _2161_;
	assign _2314_ = _2313_ | _1430_;
	assign _2316_ = \mchip.index [8] & ~_2314_;
	assign _2317_ = _1903_ | \mchip.index [6];
	assign _2318_ = \mchip.index [11] & ~_2317_;
	assign _2319_ = \mchip.index [0] | \mchip.index [6];
	assign _2320_ = _2319_ | _1430_;
	assign _2321_ = _2320_ | \mchip.index [8];
	assign _2322_ = _2321_ | \mchip.index [9];
	assign _2323_ = _2322_ | \mchip.index [10];
	assign _2324_ = _2271_ & ~_2323_;
	assign _2325_ = _2600_ | \mchip.index [3];
	assign _2327_ = _2325_ | \mchip.index [8];
	assign _2328_ = \mchip.index [9] & ~_2327_;
	assign _2329_ = _2255_ | _1430_;
	assign _2330_ = _1931_ & ~_2329_;
	assign _2331_ = _1097_ | \mchip.index [4];
	assign _2332_ = _2331_ | \mchip.index [6];
	assign _2333_ = _1931_ & ~_2332_;
	assign _2334_ = _1297_ | _2030_;
	assign _2335_ = _2334_ | \mchip.index [5];
	assign _2336_ = \mchip.index [9] & ~_2335_;
	assign _2338_ = _2185_ | \mchip.index [7];
	assign _2339_ = \mchip.index [10] & ~_2338_;
	assign _2340_ = _0428_ | \mchip.index [5];
	assign _2341_ = _2340_ | \mchip.index [7];
	assign _2342_ = \mchip.index [11] & ~_2341_;
	assign _2343_ = _1607_ | _1540_;
	assign _2344_ = _2343_ | \mchip.index [7];
	assign _2345_ = _2344_ | \mchip.index [8];
	assign _2346_ = _2345_ | \mchip.index [9];
	assign _2347_ = _2346_ | \mchip.index [10];
	assign _2349_ = _2271_ & ~_2347_;
	assign _2350_ = ~(\mchip.index [1] & \mchip.index [3]);
	assign _2351_ = _2350_ | \mchip.index [5];
	assign _2352_ = _2351_ | \mchip.index [7];
	assign _2353_ = \mchip.index [11] & ~_2352_;
	assign _2354_ = _0165_ | _2161_;
	assign _2355_ = _2354_ | _1540_;
	assign _2356_ = _1430_ & ~_2355_;
	assign _2357_ = _2356_ | _2353_;
	assign _2358_ = _2357_ | _2349_;
	assign _2360_ = _2358_ | _2342_;
	assign _2361_ = _2360_ | _2339_;
	assign _2362_ = _2361_ | _2336_;
	assign _2363_ = _2362_ | _2333_;
	assign _2364_ = _2363_ | _2330_;
	assign _2365_ = _2364_ | _2328_;
	assign _2366_ = _2365_ | _2324_;
	assign _2367_ = _2366_ | _2318_;
	assign _2368_ = _2367_ | _2316_;
	assign _2369_ = _2368_ | _2312_;
	assign _2371_ = _2369_ | _1977_;
	assign _2372_ = _2371_ | _2308_;
	assign _2373_ = _2372_ | _2307_;
	assign _2374_ = _2373_ | _2305_;
	assign _2375_ = _2374_ | _2301_;
	assign _2376_ = _2375_ | _2299_;
	assign _2377_ = _2376_ | _2297_;
	assign _2378_ = _2377_ | _2292_;
	assign _2379_ = _2378_ | _2289_;
	assign _2380_ = _2379_ | _2287_;
	assign _2382_ = _2380_ | _2280_;
	assign _2383_ = _2382_ | _2278_;
	assign _2384_ = _2383_ | _2277_;
	assign _2385_ = _2384_ | _2274_;
	assign _2386_ = _2385_ | _2269_;
	assign _2387_ = _2386_ | _2265_;
	assign _2388_ = _2387_ | _2261_;
	assign _2389_ = _2388_ | _2257_;
	assign _2390_ = _2389_ | _2254_;
	assign _2391_ = _2390_ | _2252_;
	assign _2393_ = _2391_ | _2248_;
	assign _2394_ = _2393_ | _2245_;
	assign _2395_ = _2394_ | _2243_;
	assign _2396_ = _2395_ | _2236_;
	assign _2397_ = _2396_ | _2232_;
	assign _2398_ = _2397_ | _2229_;
	assign _2399_ = _2398_ | _2226_;
	assign _2400_ = _2399_ | _2225_;
	assign _2401_ = _2400_ | _2221_;
	assign _2402_ = _2401_ | _2220_;
	assign _2404_ = _2402_ | _2218_;
	assign _2405_ = _2404_ | _2214_;
	assign _2406_ = _2405_ | _2210_;
	assign _2407_ = _2406_ | _2209_;
	assign _2408_ = _2407_ | _2207_;
	assign _2409_ = _2408_ | _2202_;
	assign _2410_ = _2409_ | _2199_;
	assign _2411_ = _2410_ | _2197_;
	assign _2412_ = _2411_ | _2196_;
	assign _2413_ = _2412_ | _2192_;
	assign _2415_ = _2413_ | _2190_;
	assign _2416_ = _2415_ | _2187_;
	assign _2417_ = _2416_ | _2184_;
	assign _2418_ = _2417_ | _2176_;
	assign _2419_ = _2418_ | _2175_;
	assign _2420_ = _2419_ | _2173_;
	assign _2421_ = _2420_ | _2096_;
	assign _2422_ = _2421_ | _2169_;
	assign _2423_ = _2422_ | _2167_;
	assign _2424_ = _2423_ | _2165_;
	assign _2426_ = _2424_ | _2160_;
	assign _2427_ = _2426_ | _2159_;
	assign _2428_ = _2427_ | _2157_;
	assign _2429_ = _2428_ | _2154_;
	assign _2430_ = _2429_ | _2149_;
	assign _2431_ = _2430_ | _2146_;
	assign _2432_ = _2431_ | _2143_;
	assign _2433_ = _2432_ | _2140_;
	assign _2434_ = _2433_ | _2138_;
	assign _2435_ = _2434_ | _2135_;
	assign \mchip.val [5] = _2435_ | _2134_;
	assign _2437_ = _1386_ | \mchip.index [4];
	assign _2438_ = _2437_ | _1540_;
	assign _2439_ = _2438_ | \mchip.index [7];
	assign _2440_ = \mchip.index [11] & ~_2439_;
	assign _2441_ = _2025_ | _2030_;
	assign _2442_ = _2441_ | _1540_;
	assign _2443_ = _2442_ | _1430_;
	assign _2444_ = \mchip.index [10] & ~_2443_;
	assign _2445_ = _2262_ | _2161_;
	assign _2447_ = _2445_ | \mchip.index [6];
	assign _2448_ = _2447_ | \mchip.index [7];
	assign _2449_ = \mchip.index [11] & ~_2448_;
	assign _2450_ = _1974_ | _2161_;
	assign _2451_ = _2271_ & ~_2450_;
	assign _2452_ = _1186_ | \mchip.index [4];
	assign _2453_ = _2452_ | \mchip.index [5];
	assign _2454_ = _2453_ | \mchip.index [6];
	assign _2455_ = _2454_ | _1430_;
	assign _2456_ = \mchip.index [11] & ~_2455_;
	assign _2458_ = _1507_ | _2567_;
	assign _2459_ = _2458_ | \mchip.index [4];
	assign _2460_ = _2459_ | \mchip.index [5];
	assign _2461_ = _2460_ | _1540_;
	assign _2462_ = \mchip.index [8] & ~_2461_;
	assign _2463_ = _1950_ | _2030_;
	assign _2464_ = _2463_ | _1540_;
	assign _2465_ = _2464_ | _1430_;
	assign _2466_ = _1319_ & ~_2465_;
	assign _2467_ = _1958_ | _1540_;
	assign _2469_ = _2467_ | _1430_;
	assign _2470_ = \mchip.index [11] & ~_2469_;
	assign _2471_ = _1629_ | _1540_;
	assign _2472_ = _2471_ | \mchip.index [7];
	assign _2473_ = _2472_ | _2359_;
	assign _2474_ = _2473_ | _1319_;
	assign _2475_ = _2474_ | _1931_;
	assign _2476_ = \mchip.index [11] & ~_2475_;
	assign _2477_ = _1751_ | _1430_;
	assign _2478_ = _2477_ | \mchip.index [9];
	assign _2480_ = _1931_ & ~_2478_;
	assign _2481_ = _0176_ | \mchip.index [3];
	assign _2482_ = _2481_ | \mchip.index [4];
	assign _2483_ = _2482_ | \mchip.index [5];
	assign _2484_ = _2483_ | \mchip.index [6];
	assign _2485_ = _2484_ | \mchip.index [7];
	assign _2486_ = _2485_ | _2359_;
	assign _2487_ = _2486_ | _1319_;
	assign _2488_ = _2487_ | \mchip.index [10];
	assign _2489_ = _2271_ & ~_2488_;
	assign _2491_ = _1980_ | _2030_;
	assign _2492_ = _2491_ | \mchip.index [5];
	assign _2493_ = _2492_ | \mchip.index [6];
	assign _2494_ = \mchip.index [8] & ~_2493_;
	assign _2495_ = _2589_ | _2567_;
	assign _2496_ = _2495_ | _2030_;
	assign _2497_ = _2496_ | _1430_;
	assign _2498_ = _1319_ & ~_2497_;
	assign _2499_ = _2481_ | _2030_;
	assign _2500_ = _2499_ | \mchip.index [7];
	assign _2502_ = _2500_ | \mchip.index [8];
	assign _2503_ = _1931_ & ~_2502_;
	assign _2504_ = _0198_ | \mchip.index [6];
	assign _2505_ = _2504_ | \mchip.index [8];
	assign _2506_ = \mchip.index [9] & ~_2505_;
	assign _2507_ = _2002_ | \mchip.index [5];
	assign _2508_ = _2507_ | \mchip.index [6];
	assign _2509_ = _2508_ | \mchip.index [7];
	assign _2510_ = \mchip.index [11] & ~_2509_;
	assign _2511_ = _0055_ | _2567_;
	assign _2513_ = _2511_ | \mchip.index [4];
	assign _2514_ = _2513_ | \mchip.index [8];
	assign _2515_ = \mchip.index [10] & ~_2514_;
	assign _2516_ = _1507_ | \mchip.index [3];
	assign _2517_ = _2516_ | \mchip.index [6];
	assign _2518_ = _2517_ | _1430_;
	assign _2519_ = \mchip.index [10] & ~_2518_;
	assign _2520_ = _1958_ | \mchip.index [5];
	assign _2521_ = _2520_ | \mchip.index [6];
	assign _2522_ = _2521_ | \mchip.index [7];
	assign _2524_ = \mchip.index [11] & ~_2522_;
	assign _2525_ = _1507_ | \mchip.index [4];
	assign _2526_ = _2525_ | _1540_;
	assign _2527_ = _2526_ | \mchip.index [7];
	assign _2528_ = _2527_ | _2359_;
	assign _2529_ = _2271_ & ~_2528_;
	assign _2530_ = _2481_ | _1540_;
	assign _2531_ = _2530_ | _1430_;
	assign _2532_ = _2531_ | _2359_;
	assign _2533_ = _2532_ | _1319_;
	assign _2535_ = _2533_ | _1931_;
	assign _2536_ = \mchip.index [11] & ~_2535_;
	assign _2537_ = _2350_ | _2030_;
	assign _2538_ = _2537_ | _1540_;
	assign _2539_ = _2538_ | _1430_;
	assign _2540_ = \mchip.index [11] & ~_2539_;
	assign _2541_ = _0187_ | _2030_;
	assign _2542_ = _2541_ | \mchip.index [5];
	assign _2543_ = _2542_ | _1540_;
	assign _2544_ = _2543_ | \mchip.index [7];
	assign _2546_ = \mchip.index [9] & ~_2544_;
	assign _2547_ = _2437_ | _2161_;
	assign _2548_ = _2547_ | \mchip.index [7];
	assign _2549_ = \mchip.index [11] & ~_2548_;
	assign _2550_ = _0878_ | \mchip.index [3];
	assign _2551_ = _2550_ | \mchip.index [4];
	assign _2552_ = _2551_ | \mchip.index [6];
	assign _2553_ = _2552_ | \mchip.index [8];
	assign _2554_ = \mchip.index [10] & ~_2553_;
	assign _2555_ = _0176_ | _2030_;
	assign _2557_ = _2555_ | \mchip.index [6];
	assign _2558_ = _2557_ | _1430_;
	assign _2559_ = _2558_ | _2359_;
	assign _2560_ = _2271_ & ~_2559_;
	assign _2561_ = _1098_ | _1540_;
	assign _2562_ = _2561_ | _1430_;
	assign _2563_ = \mchip.index [11] & ~_2562_;
	assign _2564_ = _1976_ | \mchip.index [4];
	assign _2565_ = _2564_ | _2161_;
	assign _2566_ = _2565_ | \mchip.index [6];
	assign _2568_ = \mchip.index [7] & ~_2566_;
	assign _2569_ = _1974_ | _1540_;
	assign _2570_ = _2569_ | \mchip.index [8];
	assign _2571_ = \mchip.index [9] & ~_2570_;
	assign _2572_ = _2458_ | _2030_;
	assign _2573_ = _2572_ | \mchip.index [7];
	assign _2574_ = _1931_ & ~_2573_;
	assign _2575_ = ~(_0208_ & _1319_);
	assign _2576_ = \mchip.index [10] & ~_2575_;
	assign _2577_ = _1935_ | _1430_;
	assign _2579_ = _2577_ | \mchip.index [9];
	assign _2580_ = _1931_ & ~_2579_;
	assign _2581_ = _2512_ | _1540_;
	assign _2582_ = _2581_ | \mchip.index [7];
	assign _2583_ = _2582_ | _2359_;
	assign _2584_ = _2583_ | \mchip.index [9];
	assign _2585_ = _2584_ | \mchip.index [10];
	assign _2586_ = _2271_ & ~_2585_;
	assign _2587_ = _2555_ | _1540_;
	assign _2588_ = _2587_ | _1430_;
	assign _2590_ = _1319_ & ~_2588_;
	assign _2591_ = _1563_ | _1430_;
	assign _2592_ = \mchip.index [11] & ~_2591_;
	assign _2593_ = _1980_ | \mchip.index [4];
	assign _2594_ = _2593_ | _2359_;
	assign _2595_ = _1319_ & ~_2594_;
	assign _2596_ = _1751_ | \mchip.index [5];
	assign _2597_ = _2596_ | _1540_;
	assign _2598_ = _2597_ | \mchip.index [7];
	assign _2599_ = \mchip.index [11] & ~_2598_;
	assign _2601_ = _1032_ | \mchip.index [3];
	assign _2602_ = _2601_ | \mchip.index [4];
	assign _2603_ = _2602_ | \mchip.index [6];
	assign _2604_ = _2603_ | _1430_;
	assign _2605_ = _2604_ | \mchip.index [8];
	assign _2606_ = _2605_ | \mchip.index [9];
	assign _2607_ = _2606_ | \mchip.index [10];
	assign _2608_ = _2271_ & ~_2607_;
	assign _2609_ = _1032_ | \mchip.index [4];
	assign _2610_ = _2609_ | \mchip.index [5];
	assign _2612_ = _2610_ | \mchip.index [6];
	assign _2613_ = _2612_ | \mchip.index [7];
	assign _2614_ = _2613_ | _2359_;
	assign _2615_ = _2614_ | _1319_;
	assign _2616_ = _2615_ | _1931_;
	assign _2617_ = \mchip.index [11] & ~_2616_;
	assign _2618_ = _0099_ | \mchip.index [5];
	assign _2619_ = _2618_ | \mchip.index [6];
	assign _2620_ = _2619_ | _1430_;
	assign _2621_ = \mchip.index [8] & ~_2620_;
	assign _2623_ = _1507_ | \mchip.index [6];
	assign _2624_ = _2623_ | _1430_;
	assign _2625_ = _2624_ | \mchip.index [8];
	assign _2626_ = \mchip.index [10] & ~_2625_;
	assign _2627_ = _2222_ | _1540_;
	assign _2628_ = _2627_ | \mchip.index [8];
	assign _2629_ = \mchip.index [9] & ~_2628_;
	assign _2630_ = _0648_ | \mchip.index [5];
	assign _2631_ = _2630_ | \mchip.index [6];
	assign _2632_ = _2631_ | \mchip.index [7];
	assign _2634_ = \mchip.index [11] & ~_2632_;
	assign _2635_ = _1930_ | _1540_;
	assign _2636_ = _2635_ | \mchip.index [7];
	assign _2637_ = _2636_ | _1319_;
	assign _2638_ = _1931_ & ~_2637_;
	assign _2639_ = _2222_ | _2359_;
	assign _2640_ = _2639_ | _1931_;
	assign _2641_ = _2271_ & ~_2640_;
	assign _2642_ = _2200_ | \mchip.index [5];
	assign _2643_ = _2642_ | _1540_;
	assign _2645_ = _2643_ | \mchip.index [7];
	assign _2646_ = \mchip.index [11] & ~_2645_;
	assign _2647_ = _2482_ | _1540_;
	assign _2648_ = _2647_ | _1430_;
	assign _2649_ = _2648_ | _2359_;
	assign _2650_ = _2649_ | _1319_;
	assign _2651_ = _2650_ | \mchip.index [10];
	assign _2652_ = _2271_ & ~_2651_;
	assign _2653_ = ~(\mchip.index [1] & \mchip.index [5]);
	assign _2654_ = _2653_ | _1540_;
	assign _2656_ = _2654_ | _1430_;
	assign _2657_ = \mchip.index [9] & ~_2656_;
	assign _2658_ = _1518_ | _1540_;
	assign _2659_ = _2658_ | _1430_;
	assign _2660_ = _2659_ | _2359_;
	assign _2661_ = _1931_ & ~_2660_;
	assign _2662_ = _2622_ | \mchip.index [6];
	assign _2663_ = _2662_ | _1430_;
	assign _2664_ = _2663_ | _2359_;
	assign _2665_ = _2271_ & ~_2664_;
	assign _2667_ = _2325_ | \mchip.index [4];
	assign _2668_ = _2667_ | _1540_;
	assign _2669_ = _2668_ | _1430_;
	assign _2670_ = _2669_ | _2359_;
	assign _2671_ = _2271_ & ~_2670_;
	assign _2672_ = _2511_ | _1540_;
	assign _2673_ = _2672_ | \mchip.index [7];
	assign _2674_ = _2673_ | _1319_;
	assign _2675_ = _1931_ & ~_2674_;
	assign _2676_ = _0329_ | \mchip.index [4];
	assign _2678_ = _2676_ | _1540_;
	assign _2679_ = _2678_ | \mchip.index [7];
	assign _2680_ = _2679_ | \mchip.index [8];
	assign _2681_ = _2680_ | \mchip.index [9];
	assign _2682_ = _2681_ | \mchip.index [10];
	assign _2683_ = _2271_ & ~_2682_;
	assign _2684_ = _2550_ | _2030_;
	assign _2685_ = _2684_ | _1540_;
	assign _2686_ = _2685_ | \mchip.index [7];
	assign _2687_ = _2686_ | _1931_;
	assign _2689_ = _2271_ & ~_2687_;
	assign _2690_ = _0659_ | _2359_;
	assign _2691_ = _1319_ & ~_2690_;
	assign _2692_ = _1342_ | _1540_;
	assign _2693_ = _2692_ | \mchip.index [7];
	assign _2694_ = _2693_ | \mchip.index [8];
	assign _2695_ = \mchip.index [10] & ~_2694_;
	assign _2696_ = _1097_ | _2030_;
	assign _2697_ = _2696_ | _1540_;
	assign _2698_ = _2697_ | _1430_;
	assign _0001_ = \mchip.index [11] & ~_2698_;
	assign _0002_ = _2602_ | \mchip.index [5];
	assign _0003_ = _0002_ | _1540_;
	assign _0004_ = _0003_ | _1430_;
	assign _0005_ = _0004_ | \mchip.index [8];
	assign _0006_ = _0005_ | \mchip.index [9];
	assign _0007_ = _0006_ | _1931_;
	assign _0008_ = _2271_ & ~_0007_;
	assign _0009_ = _0055_ | _2030_;
	assign _0010_ = _0009_ | \mchip.index [5];
	assign _0012_ = _0010_ | _1540_;
	assign _0013_ = \mchip.index [11] & ~_0012_;
	assign _0014_ = _1375_ | \mchip.index [4];
	assign _0015_ = _0014_ | \mchip.index [6];
	assign _0016_ = _0015_ | _1430_;
	assign _0017_ = _0016_ | _2359_;
	assign _0018_ = _2271_ & ~_0017_;
	assign _0019_ = _2441_ | \mchip.index [5];
	assign _0020_ = _0019_ | \mchip.index [6];
	assign _0021_ = _0020_ | \mchip.index [7];
	assign _0023_ = \mchip.index [11] & ~_0021_;
	assign _0024_ = _1974_ | _2030_;
	assign _0025_ = _0024_ | _1540_;
	assign _0026_ = _0025_ | \mchip.index [7];
	assign _0027_ = _0026_ | \mchip.index [9];
	assign _0028_ = \mchip.index [10] & ~_0027_;
	assign _0029_ = _1936_ | _2161_;
	assign _0030_ = \mchip.index [6] & ~_0029_;
	assign _0031_ = _0428_ | _2030_;
	assign _0032_ = _0031_ | _1540_;
	assign _0034_ = _0032_ | _1430_;
	assign _0035_ = \mchip.index [11] & ~_0034_;
	assign _0036_ = _1930_ | \mchip.index [4];
	assign _0037_ = _0036_ | _1540_;
	assign _0038_ = _0037_ | _1430_;
	assign _0039_ = \mchip.index [11] & ~_0038_;
	assign _0040_ = _2609_ | \mchip.index [6];
	assign _0041_ = _0040_ | \mchip.index [7];
	assign _0042_ = _0041_ | _2359_;
	assign _0043_ = _0042_ | \mchip.index [9];
	assign _0045_ = _0043_ | _1931_;
	assign _0046_ = _2271_ & ~_0045_;
	assign _0047_ = _2511_ | _2030_;
	assign _0048_ = \mchip.index [11] & ~_0047_;
	assign _0049_ = _2667_ | \mchip.index [6];
	assign _0050_ = _0049_ | \mchip.index [8];
	assign _0051_ = \mchip.index [9] & ~_0050_;
	assign _0052_ = _2516_ | _2030_;
	assign _0053_ = _0052_ | _1540_;
	assign _0054_ = _0053_ | \mchip.index [7];
	assign _0056_ = _0054_ | _1931_;
	assign _0057_ = _2271_ & ~_0056_;
	assign _0058_ = _0052_ | _2359_;
	assign _0059_ = _0058_ | _1931_;
	assign _0060_ = _2271_ & ~_0059_;
	assign _0061_ = _1980_ | \mchip.index [6];
	assign _0062_ = _0061_ | _1430_;
	assign _0063_ = _0062_ | _2359_;
	assign _0064_ = _1931_ & ~_0063_;
	assign _0065_ = _1974_ | _2567_;
	assign _0067_ = _0065_ | \mchip.index [4];
	assign _0068_ = _0067_ | _1430_;
	assign _0069_ = _1319_ & ~_0068_;
	assign _0070_ = _1386_ | \mchip.index [5];
	assign _0071_ = _0070_ | \mchip.index [6];
	assign _0072_ = _0071_ | _2359_;
	assign _0073_ = _1931_ & ~_0072_;
	assign _0074_ = _0593_ | _2030_;
	assign _0075_ = _0074_ | \mchip.index [8];
	assign _0076_ = \mchip.index [10] & ~_0075_;
	assign _0078_ = _2499_ | \mchip.index [6];
	assign _0079_ = _0078_ | \mchip.index [8];
	assign _0080_ = \mchip.index [9] & ~_0079_;
	assign _0081_ = _0065_ | _2030_;
	assign _0082_ = _0081_ | \mchip.index [7];
	assign _0083_ = _1931_ & ~_0082_;
	assign _0084_ = _1958_ | \mchip.index [6];
	assign _0085_ = _0084_ | \mchip.index [7];
	assign _0086_ = _2359_ & ~_0085_;
	assign _0087_ = _0955_ | \mchip.index [6];
	assign _0089_ = _0087_ | _1430_;
	assign _0090_ = _0089_ | \mchip.index [9];
	assign _0091_ = \mchip.index [10] & ~_0090_;
	assign _0092_ = _1762_ | \mchip.index [4];
	assign _0093_ = _0092_ | _1540_;
	assign _0094_ = _0093_ | _1430_;
	assign _0095_ = _2359_ & ~_0094_;
	assign _0096_ = _1997_ | _2030_;
	assign _0097_ = _0096_ | _1540_;
	assign _0098_ = _0097_ | _1430_;
	assign _0100_ = _0098_ | _2359_;
	assign _0101_ = _1931_ & ~_0100_;
	assign _0102_ = _2441_ | \mchip.index [6];
	assign _0103_ = _0102_ | _1430_;
	assign _0104_ = _0103_ | _2359_;
	assign _0105_ = _1931_ & ~_0104_;
	assign _0106_ = _2452_ | _2161_;
	assign _0107_ = _0106_ | \mchip.index [6];
	assign _0108_ = _1430_ & ~_0107_;
	assign _0109_ = _0889_ | _2161_;
	assign _0111_ = \mchip.index [6] & ~_0109_;
	assign _0112_ = _1885_ | \mchip.index [6];
	assign _0113_ = _0112_ | \mchip.index [7];
	assign _0114_ = \mchip.index [10] & ~_0113_;
	assign _0115_ = _0114_ | _0111_;
	assign _0116_ = _0115_ | _0108_;
	assign _0117_ = _0116_ | _0105_;
	assign _0118_ = _0117_ | _0101_;
	assign _0119_ = _0118_ | _0095_;
	assign _0120_ = _0119_ | _0091_;
	assign _0122_ = _0120_ | _0086_;
	assign _0123_ = _0122_ | _0083_;
	assign _0124_ = _0123_ | _0080_;
	assign _0125_ = _0124_ | _0076_;
	assign _0126_ = _0125_ | _0073_;
	assign _0127_ = _0126_ | _0069_;
	assign _0128_ = _0127_ | _0064_;
	assign _0129_ = _0128_ | _0060_;
	assign _0130_ = _0129_ | _0057_;
	assign _0131_ = _0130_ | _0051_;
	assign _0133_ = _0131_ | _0048_;
	assign _0134_ = _0133_ | _0046_;
	assign _0135_ = _0134_ | _0039_;
	assign _0136_ = _0135_ | _0035_;
	assign _0137_ = _0136_ | _0030_;
	assign _0138_ = _0137_ | _0028_;
	assign _0139_ = _0138_ | _0023_;
	assign _0140_ = _0139_ | _0018_;
	assign _0141_ = _0140_ | _0013_;
	assign _0142_ = _0141_ | _0008_;
	assign _0144_ = _0142_ | _0001_;
	assign _0145_ = _0144_ | _2695_;
	assign _0146_ = _0145_ | _2691_;
	assign _0147_ = _0146_ | _2689_;
	assign _0148_ = _0147_ | _2683_;
	assign _0149_ = _0148_ | _2675_;
	assign _0150_ = _0149_ | _2671_;
	assign _0151_ = _0150_ | _2665_;
	assign _0152_ = _0151_ | _2661_;
	assign _0153_ = _0152_ | _2657_;
	assign _0155_ = _0153_ | _2652_;
	assign _0156_ = _0155_ | _2646_;
	assign _0157_ = _0156_ | _2641_;
	assign _0158_ = _0157_ | _2638_;
	assign _0159_ = _0158_ | _2634_;
	assign _0160_ = _0159_ | _2629_;
	assign _0161_ = _0160_ | _2626_;
	assign _0162_ = _0161_ | _2621_;
	assign _0163_ = _0162_ | _2617_;
	assign _0164_ = _0163_ | _2608_;
	assign _0166_ = _0164_ | _2599_;
	assign _0167_ = _0166_ | _2595_;
	assign _0168_ = _0167_ | _2592_;
	assign _0169_ = _0168_ | _2590_;
	assign _0170_ = _0169_ | _2586_;
	assign _0171_ = _0170_ | _2580_;
	assign _0172_ = _0171_ | _2576_;
	assign _0173_ = _0172_ | _2574_;
	assign _0174_ = _0173_ | _2571_;
	assign _0175_ = _0174_ | _2568_;
	assign _0177_ = _0175_ | _2563_;
	assign _0178_ = _0177_ | _2560_;
	assign _0179_ = _0178_ | _2554_;
	assign _0180_ = _0179_ | _2549_;
	assign _0181_ = _0180_ | _2546_;
	assign _0182_ = _0181_ | _2540_;
	assign _0183_ = _0182_ | _2536_;
	assign _0184_ = _0183_ | _2529_;
	assign _0185_ = _0184_ | _2524_;
	assign _0186_ = _0185_ | _2519_;
	assign _0188_ = _0186_ | _2515_;
	assign _0189_ = _0188_ | _2510_;
	assign _0190_ = _0189_ | _2506_;
	assign _0191_ = _0190_ | _2503_;
	assign _0192_ = _0191_ | _2498_;
	assign _0193_ = _0192_ | _2494_;
	assign _0194_ = _0193_ | _2489_;
	assign _0195_ = _0194_ | _2480_;
	assign _0196_ = _0195_ | _2476_;
	assign _0197_ = _0196_ | _2470_;
	assign _0199_ = _0197_ | _2466_;
	assign _0200_ = _0199_ | _2462_;
	assign _0201_ = _0200_ | _2456_;
	assign _0202_ = _0201_ | _2451_;
	assign _0203_ = _0202_ | _2449_;
	assign _0204_ = _0203_ | _2444_;
	assign \mchip.val [4] = _0204_ | _2440_;
	assign _0205_ = _0011_ | _2030_;
	assign _0206_ = _0205_ | _1540_;
	assign _0207_ = _1430_ & ~_0206_;
	assign _0209_ = _0067_ | \mchip.index [6];
	assign _0210_ = _0209_ | _1430_;
	assign _0211_ = _0210_ | _2359_;
	assign _0212_ = _1931_ & ~_0211_;
	assign _0213_ = _2611_ | _2161_;
	assign _0214_ = _1540_ & ~_0213_;
	assign _0215_ = _2026_ | \mchip.index [6];
	assign _0216_ = _0215_ | \mchip.index [7];
	assign _0217_ = _1931_ & ~_0216_;
	assign _0218_ = _0215_ | \mchip.index [8];
	assign _0220_ = \mchip.index [9] & ~_0218_;
	assign _0221_ = _2511_ | \mchip.index [6];
	assign _0222_ = _0221_ | _1430_;
	assign _0223_ = _0222_ | _2359_;
	assign _0224_ = _2271_ & ~_0223_;
	assign _0225_ = _2564_ | \mchip.index [7];
	assign _0226_ = _2359_ & ~_0225_;
	assign _0227_ = _0198_ | _1540_;
	assign _0228_ = _0227_ | _2359_;
	assign _0229_ = _2271_ & ~_0228_;
	assign _0231_ = _1986_ | _2567_;
	assign _0232_ = _0231_ | _2030_;
	assign _0233_ = _0232_ | _1430_;
	assign _0234_ = _0233_ | _2359_;
	assign _0235_ = _1931_ & ~_0234_;
	assign _0236_ = _2611_ | \mchip.index [5];
	assign _0237_ = _0236_ | _1540_;
	assign _0238_ = _0237_ | \mchip.index [7];
	assign _0239_ = \mchip.index [11] & ~_0238_;
	assign _0240_ = ~(_2633_ & \mchip.index [10]);
	assign _0242_ = _2271_ & ~_0240_;
	assign _0243_ = _1375_ | _2030_;
	assign _0244_ = _0243_ | \mchip.index [7];
	assign _0245_ = _0244_ | _1319_;
	assign _0246_ = _1931_ & ~_0245_;
	assign _0247_ = _0231_ | \mchip.index [4];
	assign _0248_ = _0247_ | \mchip.index [5];
	assign _0249_ = _0248_ | \mchip.index [6];
	assign _0250_ = _0249_ | _1430_;
	assign _0251_ = \mchip.index [10] & ~_0250_;
	assign _0253_ = _0052_ | \mchip.index [5];
	assign _0254_ = _0253_ | \mchip.index [6];
	assign _0255_ = _0254_ | \mchip.index [7];
	assign _0256_ = \mchip.index [11] & ~_0255_;
	assign _0257_ = _1851_ | _2161_;
	assign _0258_ = \mchip.index [6] & ~_0257_;
	assign _0259_ = _2511_ | _1430_;
	assign _0260_ = _0259_ | \mchip.index [9];
	assign _0261_ = _1931_ & ~_0260_;
	assign _0262_ = _2551_ | _1540_;
	assign _0264_ = _0262_ | _2359_;
	assign _0265_ = _2271_ & ~_0264_;
	assign _0266_ = _1796_ | _2161_;
	assign _0267_ = _0266_ | \mchip.index [6];
	assign _0268_ = \mchip.index [7] & ~_0267_;
	assign _0269_ = _0626_ | \mchip.index [7];
	assign _0270_ = \mchip.index [10] & ~_0269_;
	assign _0271_ = _0031_ | \mchip.index [5];
	assign _0272_ = _0271_ | \mchip.index [6];
	assign _0273_ = _0272_ | _1430_;
	assign _0275_ = \mchip.index [11] & ~_0273_;
	assign _0276_ = \mchip.index [10] & ~_2502_;
	assign _0277_ = _0262_ | \mchip.index [8];
	assign _0278_ = \mchip.index [10] & ~_0277_;
	assign _0279_ = _1958_ | _2359_;
	assign _0280_ = _0279_ | _1931_;
	assign _0281_ = _2271_ & ~_0280_;
	assign _0282_ = _2026_ | _1540_;
	assign _0283_ = _0282_ | _1430_;
	assign _0284_ = _0283_ | _2359_;
	assign _0286_ = _2271_ & ~_0284_;
	assign _0287_ = _1552_ | _1540_;
	assign _0288_ = _0287_ | _1430_;
	assign _0289_ = _1319_ & ~_0288_;
	assign _0290_ = _1431_ | \mchip.index [5];
	assign _0291_ = _0290_ | \mchip.index [6];
	assign _0292_ = _0291_ | \mchip.index [7];
	assign _0293_ = _1931_ & ~_0292_;
	assign _0294_ = _0047_ | \mchip.index [6];
	assign _0295_ = _1319_ & ~_0294_;
	assign _0297_ = _0016_ | \mchip.index [8];
	assign _0298_ = \mchip.index [10] & ~_0297_;
	assign _0299_ = _2593_ | \mchip.index [5];
	assign _0300_ = _0299_ | \mchip.index [6];
	assign _0301_ = _0300_ | \mchip.index [7];
	assign _0302_ = \mchip.index [11] & ~_0301_;
	assign _0303_ = _0231_ | _1540_;
	assign _0304_ = _0303_ | \mchip.index [7];
	assign _0305_ = _0304_ | _2359_;
	assign _0306_ = _1931_ & ~_0305_;
	assign _0308_ = _1957_ | \mchip.index [3];
	assign _0309_ = _0308_ | _2030_;
	assign _0310_ = _0309_ | \mchip.index [6];
	assign _0311_ = _0310_ | _1430_;
	assign _0312_ = \mchip.index [8] & ~_0311_;
	assign _0313_ = _2611_ | _2030_;
	assign _0314_ = _0313_ | _1540_;
	assign _0315_ = \mchip.index [11] & ~_0314_;
	assign _0316_ = _2572_ | \mchip.index [6];
	assign _0317_ = _0316_ | _1430_;
	assign _0319_ = _0317_ | _2359_;
	assign _0320_ = _1931_ & ~_0319_;
	assign _0321_ = _0176_ | \mchip.index [4];
	assign _0322_ = _0321_ | \mchip.index [5];
	assign _0323_ = _0322_ | \mchip.index [6];
	assign _0324_ = _0323_ | _1430_;
	assign _0325_ = _0324_ | \mchip.index [8];
	assign _0326_ = _0325_ | \mchip.index [9];
	assign _0327_ = _0326_ | _1931_;
	assign _0328_ = _2271_ & ~_0327_;
	assign _0330_ = _1375_ | _2567_;
	assign _0331_ = _0330_ | _1540_;
	assign _0332_ = _0331_ | \mchip.index [7];
	assign _0333_ = _0332_ | _1319_;
	assign _0334_ = _1931_ & ~_0333_;
	assign _0335_ = _2155_ | \mchip.index [6];
	assign _0336_ = _0335_ | \mchip.index [7];
	assign _0337_ = _2359_ & ~_0336_;
	assign _0338_ = _0009_ | _1430_;
	assign _0339_ = _0338_ | _2359_;
	assign _0341_ = _2271_ & ~_0339_;
	assign _0342_ = _2359_ & ~_2355_;
	assign _0343_ = \mchip.index [6] & ~_0106_;
	assign _0344_ = _0011_ | \mchip.index [7];
	assign _0345_ = _0344_ | _2359_;
	assign _0346_ = _1931_ & ~_0345_;
	assign _0347_ = _0052_ | \mchip.index [6];
	assign _0348_ = _2359_ & ~_0347_;
	assign _0349_ = _2200_ | _2030_;
	assign _0350_ = _0349_ | _2359_;
	assign _0352_ = _0350_ | _1931_;
	assign _0353_ = _2271_ & ~_0352_;
	assign _0354_ = _2622_ | _1540_;
	assign _0355_ = _0354_ | _1430_;
	assign _0356_ = _1931_ & ~_0355_;
	assign _0357_ = _2630_ | _1540_;
	assign _0358_ = _0357_ | _1430_;
	assign _0359_ = \mchip.index [11] & ~_0358_;
	assign _0360_ = _2601_ | _2030_;
	assign _0361_ = _0360_ | \mchip.index [5];
	assign _0363_ = _0361_ | \mchip.index [6];
	assign _0364_ = _0363_ | _1430_;
	assign _0365_ = \mchip.index [11] & ~_0364_;
	assign _0366_ = _2495_ | \mchip.index [4];
	assign _0367_ = _0366_ | \mchip.index [6];
	assign _0368_ = _0367_ | \mchip.index [7];
	assign _0369_ = _1931_ & ~_0368_;
	assign _0370_ = _2516_ | \mchip.index [4];
	assign _0371_ = _0370_ | _2359_;
	assign _0372_ = _0371_ | \mchip.index [9];
	assign _0374_ = \mchip.index [10] & ~_0372_;
	assign _0375_ = _2589_ | _2030_;
	assign _0376_ = _0375_ | \mchip.index [9];
	assign _0377_ = _1931_ & ~_0376_;
	assign _0378_ = _2648_ | \mchip.index [8];
	assign _0379_ = _0378_ | _1319_;
	assign _0380_ = _0379_ | \mchip.index [10];
	assign _0381_ = _2271_ & ~_0380_;
	assign _0382_ = _0889_ | \mchip.index [5];
	assign _0383_ = _0382_ | \mchip.index [6];
	assign _0385_ = _0383_ | _1430_;
	assign _0386_ = \mchip.index [8] & ~_0385_;
	assign _0387_ = _1386_ | _2030_;
	assign _0388_ = _0387_ | _1540_;
	assign _0389_ = _1430_ & ~_0388_;
	assign _0390_ = _0389_ & ~_1931_;
	assign _0391_ = _0088_ | \mchip.index [6];
	assign _0392_ = _0391_ | \mchip.index [8];
	assign _0393_ = \mchip.index [9] & ~_0392_;
	assign _0394_ = _0370_ | _2161_;
	assign _0396_ = _1540_ & ~_0394_;
	assign _0397_ = ~(_0396_ & _1430_);
	assign _0398_ = \mchip.index [11] & ~_0397_;
	assign _0399_ = _1442_ | _1430_;
	assign _0400_ = _0399_ | \mchip.index [8];
	assign _0401_ = \mchip.index [10] & ~_0400_;
	assign _0402_ = _2026_ | \mchip.index [7];
	assign _0403_ = _0402_ | \mchip.index [8];
	assign _0404_ = _1931_ & ~_0403_;
	assign _0405_ = _1948_ | \mchip.index [7];
	assign _0407_ = \mchip.index [11] & ~_0405_;
	assign _0408_ = _2501_ | _2030_;
	assign _0409_ = _0408_ | _1540_;
	assign _0410_ = _0409_ | _2359_;
	assign _0411_ = _1319_ & ~_0410_;
	assign _0412_ = _2600_ | _2030_;
	assign _0413_ = _0412_ | _2359_;
	assign _0414_ = _1319_ & ~_0413_;
	assign _0415_ = \mchip.index [5] & ~_2696_;
	assign _0416_ = _0388_ | \mchip.index [8];
	assign _0418_ = \mchip.index [10] & ~_0416_;
	assign _0419_ = _0096_ | \mchip.index [6];
	assign _0420_ = _0419_ | \mchip.index [8];
	assign _0421_ = \mchip.index [9] & ~_0420_;
	assign _0422_ = _2619_ | \mchip.index [7];
	assign _0423_ = _1931_ & ~_0422_;
	assign _0424_ = _2491_ | _1540_;
	assign _0425_ = _0424_ | _1430_;
	assign _0426_ = \mchip.index [11] & ~_0425_;
	assign _0427_ = _0053_ | _1430_;
	assign _0429_ = \mchip.index [9] & ~_0427_;
	assign _0430_ = _0412_ | _1540_;
	assign _0431_ = _0430_ | \mchip.index [7];
	assign _0432_ = \mchip.index [8] & ~_0431_;
	assign _0433_ = _0024_ | _2161_;
	assign _0434_ = _1540_ & ~_0433_;
	assign _0435_ = \mchip.index [7] & ~_0257_;
	assign _0436_ = _2467_ | \mchip.index [8];
	assign _0437_ = \mchip.index [9] & ~_0436_;
	assign _0438_ = _1507_ | _1430_;
	assign _0440_ = _0438_ | \mchip.index [9];
	assign _0441_ = _1931_ & ~_0440_;
	assign _0442_ = _2557_ | \mchip.index [8];
	assign _0443_ = \mchip.index [9] & ~_0442_;
	assign _0444_ = _0387_ | \mchip.index [6];
	assign _0445_ = _1931_ & ~_0444_;
	assign _0446_ = _1930_ | _2161_;
	assign _0447_ = \mchip.index [7] & ~_0446_;
	assign _0448_ = _0036_ | \mchip.index [8];
	assign _0449_ = _0448_ | \mchip.index [9];
	assign _0451_ = _1931_ & ~_0449_;
	assign _0452_ = _1552_ | _2359_;
	assign _0453_ = _1319_ & ~_0452_;
	assign _0454_ = _2550_ | _1430_;
	assign _0455_ = _0454_ | \mchip.index [9];
	assign _0456_ = _1931_ & ~_0455_;
	assign _0457_ = _2230_ | _2030_;
	assign _0458_ = _0457_ | \mchip.index [6];
	assign _0459_ = _1319_ & ~_0458_;
	assign _0460_ = _2564_ | \mchip.index [5];
	assign _0462_ = _0460_ | _1540_;
	assign _0463_ = _0462_ | _2359_;
	assign _0464_ = \mchip.index [9] & ~_0463_;
	assign _0465_ = _2600_ | _1540_;
	assign _0466_ = _0465_ | \mchip.index [8];
	assign _0467_ = \mchip.index [9] & ~_0466_;
	assign _0468_ = _0944_ | _2161_;
	assign _0469_ = _0468_ | _1540_;
	assign _0470_ = _1430_ & ~_0469_;
	assign _0471_ = _2262_ | \mchip.index [6];
	assign _0473_ = _0471_ | _1430_;
	assign _0474_ = _0473_ | _2359_;
	assign _0475_ = _1931_ & ~_0474_;
	assign _0476_ = _0215_ | _1430_;
	assign _0477_ = _0476_ | \mchip.index [9];
	assign _0478_ = \mchip.index [10] & ~_0477_;
	assign _0479_ = _1442_ | \mchip.index [8];
	assign _0480_ = \mchip.index [9] & ~_0479_;
	assign _0481_ = _0370_ | \mchip.index [5];
	assign _0482_ = _0481_ | _1540_;
	assign _0484_ = \mchip.index [10] & ~_0482_;
	assign _0485_ = _2298_ | \mchip.index [8];
	assign _0486_ = \mchip.index [9] & ~_0485_;
	assign _0487_ = _2166_ | _2161_;
	assign _0488_ = \mchip.index [6] & ~_0487_;
	assign _0489_ = _0032_ | \mchip.index [7];
	assign _0490_ = _0489_ | _1319_;
	assign _0491_ = _2271_ & ~_0490_;
	assign _0492_ = _0330_ | \mchip.index [4];
	assign _0493_ = _0492_ | \mchip.index [5];
	assign _0495_ = _0493_ | _1540_;
	assign _0496_ = _0495_ | \mchip.index [7];
	assign _0497_ = \mchip.index [10] & ~_0496_;
	assign _0498_ = _0340_ | \mchip.index [5];
	assign _0499_ = _0498_ | _1540_;
	assign _0500_ = _0499_ | \mchip.index [7];
	assign _0501_ = \mchip.index [11] & ~_0500_;
	assign _0502_ = _2359_ & ~_2573_;
	assign _0503_ = _2002_ | \mchip.index [9];
	assign _0504_ = _1931_ & ~_0503_;
	assign _0506_ = _0198_ | \mchip.index [5];
	assign _0507_ = _0506_ | _1540_;
	assign _0508_ = _1430_ & ~_0507_;
	assign _0509_ = _0011_ | \mchip.index [6];
	assign _0510_ = _0509_ | \mchip.index [7];
	assign _0511_ = _2359_ & ~_0510_;
	assign _0512_ = _1319_ & ~_2639_;
	assign _0513_ = _2525_ | \mchip.index [5];
	assign _0514_ = _0513_ | _1540_;
	assign _0515_ = _0514_ | _1430_;
	assign _0517_ = _1319_ & ~_0515_;
	assign _0518_ = _1976_ | \mchip.index [5];
	assign _0519_ = _0518_ | \mchip.index [6];
	assign _0520_ = _0519_ | _1430_;
	assign _0521_ = \mchip.index [11] & ~_0520_;
	assign _0522_ = _0232_ | \mchip.index [6];
	assign _0523_ = _0522_ | _1430_;
	assign _0524_ = \mchip.index [8] & ~_0523_;
	assign _0525_ = _2309_ | \mchip.index [6];
	assign _0526_ = _0525_ | \mchip.index [7];
	assign _0528_ = _2359_ & ~_0526_;
	assign _0529_ = _0330_ | _2030_;
	assign _0530_ = _0529_ | _1430_;
	assign _0531_ = \mchip.index [11] & ~_0530_;
	assign _0532_ = _1927_ | \mchip.index [4];
	assign _0533_ = _0532_ | \mchip.index [5];
	assign _0534_ = _0533_ | \mchip.index [6];
	assign _0535_ = _0534_ | \mchip.index [7];
	assign _0536_ = \mchip.index [11] & ~_0535_;
	assign _0537_ = _0000_ | _2030_;
	assign _0539_ = _0537_ | _1540_;
	assign _0540_ = _0539_ | \mchip.index [7];
	assign _0541_ = _1319_ & ~_0540_;
	assign _0542_ = _2002_ | _2161_;
	assign _0543_ = _1540_ & ~_0542_;
	assign _0544_ = _1930_ | \mchip.index [6];
	assign _0545_ = _0544_ | \mchip.index [7];
	assign _0546_ = _2359_ & ~_0545_;
	assign _0547_ = _2676_ | \mchip.index [6];
	assign _0548_ = _0547_ | _1430_;
	assign _0550_ = _0548_ | _2359_;
	assign _0551_ = _0550_ | _1319_;
	assign _0552_ = _0551_ | \mchip.index [10];
	assign _0553_ = _2271_ & ~_0552_;
	assign _0554_ = _0025_ | \mchip.index [8];
	assign _0555_ = \mchip.index [9] & ~_0554_;
	assign _0556_ = _0555_ | _0553_;
	assign _0557_ = _0556_ | _0546_;
	assign _0558_ = _0557_ | _0543_;
	assign _0559_ = _0558_ | _0541_;
	assign _0561_ = _0559_ | _0536_;
	assign _0562_ = _0561_ | _0531_;
	assign _0563_ = _0562_ | _0528_;
	assign _0564_ = _0563_ | _0524_;
	assign _0565_ = _0564_ | _0521_;
	assign _0566_ = _0565_ | _0517_;
	assign _0567_ = _0566_ | _0512_;
	assign _0568_ = _0567_ | _0511_;
	assign _0569_ = _0568_ | _0508_;
	assign _0570_ = _0569_ | _0504_;
	assign _0572_ = _0570_ | _0502_;
	assign _0573_ = _0572_ | _0501_;
	assign _0574_ = _0573_ | _0497_;
	assign _0575_ = _0574_ | _0491_;
	assign _0576_ = _0575_ | _0488_;
	assign _0577_ = _0576_ | _0486_;
	assign _0578_ = _0577_ | _0484_;
	assign _0579_ = _0578_ | _0480_;
	assign _0580_ = _0579_ | _0478_;
	assign _0581_ = _0580_ | _0475_;
	assign _0583_ = _0581_ | _0470_;
	assign _0584_ = _0583_ | _0467_;
	assign _0585_ = _0584_ | _0464_;
	assign _0586_ = _0585_ | _0459_;
	assign _0587_ = _0586_ | _0456_;
	assign _0588_ = _0587_ | _0453_;
	assign _0589_ = _0588_ | _0451_;
	assign _0590_ = _0589_ | _0447_;
	assign _0591_ = _0590_ | _0445_;
	assign _0592_ = _0591_ | _0443_;
	assign _0594_ = _0592_ | _0441_;
	assign _0595_ = _0594_ | _0437_;
	assign _0596_ = _0595_ | _0435_;
	assign _0597_ = _0596_ | _0434_;
	assign _0598_ = _0597_ | _0432_;
	assign _0599_ = _0598_ | _0429_;
	assign _0600_ = _0599_ | _0426_;
	assign _0601_ = _0600_ | _0423_;
	assign _0602_ = _0601_ | _0421_;
	assign _0603_ = _0602_ | _0418_;
	assign _0605_ = _0603_ | _0415_;
	assign _0606_ = _0605_ | _0414_;
	assign _0607_ = _0606_ | _0411_;
	assign _0608_ = _0607_ | _0407_;
	assign _0609_ = _0608_ | _0404_;
	assign _0610_ = _0609_ | _0401_;
	assign _0611_ = _0610_ | _0398_;
	assign _0612_ = _0611_ | _0393_;
	assign _0613_ = _0612_ | _0390_;
	assign _0614_ = _0613_ | _0386_;
	assign _0616_ = _0614_ | _0381_;
	assign _0617_ = _0616_ | _0377_;
	assign _0618_ = _0617_ | _0374_;
	assign _0619_ = _0618_ | _0369_;
	assign _0620_ = _0619_ | _0365_;
	assign _0621_ = _0620_ | _0359_;
	assign _0622_ = _0621_ | _0356_;
	assign _0623_ = _0622_ | _0353_;
	assign _0624_ = _0623_ | _0348_;
	assign _0625_ = _0624_ | _0346_;
	assign _0627_ = _0625_ | _0343_;
	assign _0628_ = _0627_ | _0342_;
	assign _0629_ = _0628_ | _0341_;
	assign _0630_ = _0629_ | _0337_;
	assign _0631_ = _0630_ | _0334_;
	assign _0632_ = _0631_ | _0328_;
	assign _0633_ = _0632_ | _0320_;
	assign _0634_ = _0633_ | _0315_;
	assign _0635_ = _0634_ | _0312_;
	assign _0636_ = _0635_ | _0306_;
	assign _0638_ = _0636_ | _0302_;
	assign _0639_ = _0638_ | _0298_;
	assign _0640_ = _0639_ | _0295_;
	assign _0641_ = _0640_ | _0293_;
	assign _0642_ = _0641_ | _0289_;
	assign _0643_ = _0642_ | _0286_;
	assign _0644_ = _0643_ | _0281_;
	assign _0645_ = _0644_ | _0278_;
	assign _0646_ = _0645_ | _0276_;
	assign _0647_ = _0646_ | _0275_;
	assign _0649_ = _0647_ | _0270_;
	assign _0650_ = _0649_ | _0268_;
	assign _0651_ = _0650_ | _0265_;
	assign _0652_ = _0651_ | _0261_;
	assign _0653_ = _0652_ | _0258_;
	assign _0654_ = _0653_ | _0256_;
	assign _0655_ = _0654_ | _0251_;
	assign _0656_ = _0655_ | _0246_;
	assign _0657_ = _0656_ | _0242_;
	assign _0658_ = _0657_ | _0239_;
	assign _0660_ = _0658_ | _0235_;
	assign _0661_ = _0660_ | _0229_;
	assign _0662_ = _0661_ | _0226_;
	assign _0663_ = _0662_ | _0224_;
	assign _0664_ = _0663_ | _0220_;
	assign _0665_ = _0664_ | _0217_;
	assign _0666_ = _0665_ | _0214_;
	assign _0667_ = _0666_ | _0212_;
	assign \mchip.val [3] = _0667_ | _0207_;
	assign _0668_ = _0065_ | _2359_;
	assign _0670_ = _1319_ & ~_0668_;
	assign _0671_ = _0205_ | _1430_;
	assign _0672_ = \mchip.index [11] & ~_0671_;
	assign _0673_ = _0757_ | _2161_;
	assign _0674_ = _1540_ & ~_0673_;
	assign _0675_ = _2697_ | \mchip.index [7];
	assign _0676_ = _1931_ & ~_0675_;
	assign _0677_ = _0911_ & ~\mchip.index [10];
	assign _0678_ = _2325_ | _2030_;
	assign _0679_ = _0678_ | \mchip.index [7];
	assign _0681_ = _1931_ & ~_0679_;
	assign _0682_ = _0036_ | \mchip.index [6];
	assign _0683_ = _0682_ | \mchip.index [7];
	assign _0684_ = _1931_ & ~_0683_;
	assign _0685_ = _0529_ | \mchip.index [6];
	assign _0686_ = _0685_ | _1430_;
	assign _0687_ = \mchip.index [11] & ~_0686_;
	assign _0688_ = _0024_ | \mchip.index [5];
	assign _0689_ = _0688_ | \mchip.index [6];
	assign _0690_ = _0689_ | \mchip.index [7];
	assign _0692_ = \mchip.index [11] & ~_0690_;
	assign _0693_ = _1707_ | _2161_;
	assign _0694_ = _0693_ | \mchip.index [6];
	assign _0695_ = _1430_ & ~_0694_;
	assign _0696_ = _0321_ | _1540_;
	assign _0697_ = _0696_ | \mchip.index [7];
	assign _0698_ = _0697_ | \mchip.index [9];
	assign _0699_ = _0698_ | \mchip.index [10];
	assign _0700_ = _2271_ & ~_0699_;
	assign _0701_ = _0532_ | _1540_;
	assign _0703_ = _0701_ | _1430_;
	assign _0704_ = \mchip.index [11] & ~_0703_;
	assign _0705_ = _2200_ | \mchip.index [4];
	assign _0706_ = _0705_ | _1540_;
	assign _0707_ = _0706_ | _1430_;
	assign _0708_ = _1319_ & ~_0707_;
	assign _0709_ = _0065_ | _2161_;
	assign _0710_ = _0709_ | \mchip.index [6];
	assign _0711_ = _1430_ & ~_0710_;
	assign _0712_ = \mchip.index [11] & ~_0495_;
	assign _0714_ = _0878_ | \mchip.index [6];
	assign _0715_ = _0714_ | \mchip.index [7];
	assign _0716_ = _2359_ & ~_0715_;
	assign _0717_ = _0678_ | _1540_;
	assign _0718_ = _1931_ & ~_0717_;
	assign _0719_ = _2222_ | \mchip.index [4];
	assign _0720_ = _0719_ | \mchip.index [6];
	assign _0721_ = _0720_ | _1430_;
	assign _0722_ = _0721_ | _1931_;
	assign _0723_ = _2271_ & ~_0722_;
	assign _0725_ = _0705_ | _2161_;
	assign _0726_ = _0725_ | _1540_;
	assign _0727_ = _1430_ & ~_0726_;
	assign _0728_ = _2491_ | \mchip.index [6];
	assign _0729_ = _0728_ | \mchip.index [8];
	assign _0730_ = \mchip.index [9] & ~_0729_;
	assign _0731_ = \mchip.index [3] | ~\mchip.index [2];
	assign _0732_ = _0731_ | \mchip.index [4];
	assign _0733_ = _0732_ | \mchip.index [5];
	assign _0734_ = _0733_ | _1540_;
	assign _0736_ = _0734_ | _1430_;
	assign _0737_ = \mchip.index [11] & ~_0736_;
	assign _0738_ = _0560_ | _1540_;
	assign _0739_ = _0738_ | \mchip.index [7];
	assign _0740_ = \mchip.index [11] & ~_0739_;
	assign _0741_ = _1958_ | _2161_;
	assign _0742_ = _1430_ & ~_0741_;
	assign _0743_ = _1043_ | \mchip.index [4];
	assign _0744_ = _0743_ | \mchip.index [5];
	assign _0745_ = _0744_ | _1540_;
	assign _0747_ = _0745_ | \mchip.index [7];
	assign _0748_ = \mchip.index [11] & ~_0747_;
	assign _0749_ = _0221_ | \mchip.index [7];
	assign _0750_ = _2359_ & ~_0749_;
	assign _0751_ = _1297_ | _1430_;
	assign _0752_ = _0751_ | \mchip.index [9];
	assign _0753_ = _1931_ & ~_0752_;
	assign _0754_ = _0187_ | \mchip.index [8];
	assign _0755_ = \mchip.index [9] & ~_0754_;
	assign _0756_ = _1430_ & ~_0717_;
	assign _0758_ = _0889_ | _1540_;
	assign _0759_ = _0758_ | _2359_;
	assign _0760_ = _2271_ & ~_0759_;
	assign _0761_ = _0758_ | _1430_;
	assign _0762_ = \mchip.index [8] & ~_0761_;
	assign _0763_ = _2230_ | \mchip.index [4];
	assign _0764_ = _0763_ | _1430_;
	assign _0765_ = _1319_ & ~_0764_;
	assign _0766_ = \mchip.index [11] & ~_2558_;
	assign _0767_ = _0705_ | \mchip.index [5];
	assign _0769_ = _0767_ | \mchip.index [6];
	assign _0770_ = _0769_ | _2359_;
	assign _0771_ = \mchip.index [10] & ~_0770_;
	assign _0772_ = _2458_ | \mchip.index [7];
	assign _0773_ = _1931_ & ~_0772_;
	assign _0774_ = _2593_ | _1430_;
	assign _0775_ = _0774_ | \mchip.index [9];
	assign _0776_ = _1931_ & ~_0775_;
	assign _0777_ = \mchip.index [5] & ~_1098_;
	assign _0778_ = _2496_ | _1540_;
	assign _0780_ = _0778_ | _1430_;
	assign _0781_ = _1319_ & ~_0780_;
	assign _0782_ = _2499_ | _1540_;
	assign _0783_ = _0782_ | _1430_;
	assign _0784_ = _2359_ & ~_0783_;
	assign _0785_ = _0227_ | _1430_;
	assign _0786_ = _2271_ & ~_0785_;
	assign _0787_ = _1431_ | _2161_;
	assign _0788_ = _0787_ | \mchip.index [6];
	assign _0789_ = \mchip.index [7] & ~_0788_;
	assign _0791_ = _0000_ | \mchip.index [4];
	assign _0792_ = _0791_ | _1540_;
	assign _0793_ = _0792_ | \mchip.index [7];
	assign _0794_ = \mchip.index [11] & ~_0793_;
	assign _0795_ = _1959_ | _1430_;
	assign _0796_ = _0795_ | _2359_;
	assign _0797_ = _2271_ & ~_0796_;
	assign _0798_ = _1707_ | \mchip.index [5];
	assign _0799_ = _0798_ | _1540_;
	assign _0800_ = _0799_ | \mchip.index [7];
	assign _0802_ = \mchip.index [11] & ~_0800_;
	assign _0803_ = _1862_ | \mchip.index [8];
	assign _0804_ = _1931_ & ~_0803_;
	assign _0805_ = _0370_ | _1540_;
	assign _0806_ = \mchip.index [11] & ~_0805_;
	assign _0807_ = _2467_ | \mchip.index [9];
	assign _0808_ = _1931_ & ~_0807_;
	assign _0809_ = _1431_ | _1540_;
	assign _0810_ = _0809_ | \mchip.index [7];
	assign _0811_ = _0810_ | _1319_;
	assign _0813_ = _2271_ & ~_0811_;
	assign _0814_ = _2331_ | _1540_;
	assign _0815_ = _0814_ | _1430_;
	assign _0816_ = _0815_ | _2359_;
	assign _0817_ = _1931_ & ~_0816_;
	assign _0818_ = _0481_ | _1430_;
	assign _0819_ = \mchip.index [10] & ~_0818_;
	assign _0820_ = _1927_ | _2161_;
	assign _0821_ = \mchip.index [7] & ~_0820_;
	assign _0822_ = _0068_ | _2359_;
	assign _0824_ = _1931_ & ~_0822_;
	assign _0825_ = _2141_ | _2359_;
	assign _0826_ = _1319_ & ~_0825_;
	assign _0827_ = _0219_ | _2359_;
	assign _0828_ = _1319_ & ~_0827_;
	assign _0829_ = _1518_ | \mchip.index [5];
	assign _0830_ = _0829_ | \mchip.index [7];
	assign _0831_ = \mchip.index [11] & ~_0830_;
	assign _0832_ = _0205_ | \mchip.index [6];
	assign _0833_ = _1319_ & ~_0832_;
	assign _0835_ = _2227_ | \mchip.index [6];
	assign _0836_ = _0835_ | \mchip.index [7];
	assign _0837_ = _1931_ & ~_0836_;
	assign _0838_ = _0351_ | _2359_;
	assign _0839_ = _1319_ & ~_0838_;
	assign _0840_ = _2174_ | \mchip.index [7];
	assign _0841_ = _2271_ & ~_0840_;
	assign _0842_ = _2633_ & ~_2271_;
	assign _0843_ = _2438_ | _2359_;
	assign _0844_ = _2271_ & ~_0843_;
	assign _0846_ = _1430_ & ~_0294_;
	assign _0847_ = _0247_ | \mchip.index [6];
	assign _0848_ = _0847_ | \mchip.index [8];
	assign _0849_ = \mchip.index [9] & ~_0848_;
	assign _0850_ = _0593_ | \mchip.index [6];
	assign _0851_ = _0850_ | _1430_;
	assign _0852_ = \mchip.index [10] & ~_0851_;
	assign _0853_ = _2516_ | \mchip.index [5];
	assign _0854_ = _0853_ | \mchip.index [7];
	assign _0855_ = _0854_ | _2359_;
	assign _0857_ = \mchip.index [10] & ~_0855_;
	assign _0858_ = _0853_ | _1540_;
	assign _0859_ = \mchip.index [11] & ~_0858_;
	assign _0860_ = \mchip.index [5] & ~_2600_;
	assign _0861_ = _2022_ | _1931_;
	assign _0862_ = _2271_ & ~_0861_;
	assign _0863_ = _2359_ & ~_2293_;
	assign _0864_ = _2612_ | _1430_;
	assign _0865_ = _0864_ | \mchip.index [8];
	assign _0866_ = _0865_ | \mchip.index [9];
	assign _0868_ = _0866_ | _1931_;
	assign _0869_ = _2271_ & ~_0868_;
	assign _0870_ = _0092_ | _2359_;
	assign _0871_ = _0870_ | \mchip.index [9];
	assign _0872_ = \mchip.index [10] & ~_0871_;
	assign _0873_ = _0439_ | \mchip.index [6];
	assign _0874_ = _0873_ | _1430_;
	assign _0875_ = _0874_ | \mchip.index [8];
	assign _0876_ = \mchip.index [10] & ~_0875_;
	assign _0877_ = _0187_ | \mchip.index [6];
	assign _0879_ = _0877_ | _1430_;
	assign _0880_ = \mchip.index [10] & ~_0879_;
	assign _0881_ = _2132_ | \mchip.index [6];
	assign _0882_ = _0881_ | _1430_;
	assign _0883_ = _0882_ | _1931_;
	assign _0884_ = _2271_ & ~_0883_;
	assign _0885_ = _0081_ | _1540_;
	assign _0886_ = _1931_ & ~_0885_;
	assign _0887_ = _0682_ | \mchip.index [8];
	assign _0888_ = _1931_ & ~_0887_;
	assign _0890_ = _2684_ | \mchip.index [6];
	assign _0891_ = _0890_ | \mchip.index [8];
	assign _0892_ = \mchip.index [10] & ~_0891_;
	assign _0893_ = _2512_ | \mchip.index [5];
	assign _0894_ = _0893_ | \mchip.index [6];
	assign _0895_ = _0894_ | _2359_;
	assign _0896_ = _0895_ | _1319_;
	assign _0897_ = _0896_ | \mchip.index [10];
	assign _0898_ = _2271_ & ~_0897_;
	assign _0899_ = _2331_ | \mchip.index [5];
	assign _0901_ = _0899_ | \mchip.index [6];
	assign _0902_ = _0901_ | \mchip.index [7];
	assign _0903_ = \mchip.index [11] & ~_0902_;
	assign _0904_ = _2655_ | \mchip.index [9];
	assign _0905_ = _1931_ & ~_0904_;
	assign _0906_ = _2266_ | _2161_;
	assign _0907_ = _1540_ & ~_0906_;
	assign _0908_ = _2551_ | \mchip.index [8];
	assign _0909_ = \mchip.index [9] & ~_0908_;
	assign _0910_ = _0078_ | \mchip.index [7];
	assign _0912_ = _2271_ & ~_0910_;
	assign _0913_ = _1518_ | \mchip.index [7];
	assign _0914_ = _0913_ | \mchip.index [8];
	assign _0915_ = \mchip.index [10] & ~_0914_;
	assign _0916_ = _2041_ | _1540_;
	assign _0917_ = _0916_ | _1430_;
	assign _0918_ = \mchip.index [10] & ~_0917_;
	assign _0919_ = _2300_ | \mchip.index [7];
	assign _0920_ = \mchip.index [11] & ~_0919_;
	assign _0921_ = _1386_ | \mchip.index [6];
	assign _0923_ = _0921_ | \mchip.index [8];
	assign _0924_ = \mchip.index [9] & ~_0923_;
	assign _0925_ = _0604_ | _1540_;
	assign _0926_ = _0925_ | \mchip.index [7];
	assign _0927_ = _2359_ & ~_0926_;
	assign _0928_ = _2436_ | \mchip.index [4];
	assign _0929_ = _0928_ | \mchip.index [6];
	assign _0930_ = _0929_ | \mchip.index [8];
	assign _0931_ = \mchip.index [9] & ~_0930_;
	assign _0932_ = _0344_ | _1319_;
	assign _0934_ = _1931_ & ~_0932_;
	assign _0935_ = _2643_ | _1430_;
	assign _0936_ = \mchip.index [11] & ~_0935_;
	assign _0937_ = _2550_ | _1540_;
	assign _0938_ = _0937_ | \mchip.index [9];
	assign _0939_ = _1931_ & ~_0938_;
	assign _0940_ = _2193_ | \mchip.index [6];
	assign _0941_ = _0940_ | _2359_;
	assign _0942_ = _1931_ & ~_0941_;
	assign _0943_ = _1950_ | _2161_;
	assign _0945_ = \mchip.index [7] & ~_0943_;
	assign _0946_ = _2589_ | \mchip.index [4];
	assign _0947_ = _0946_ | \mchip.index [5];
	assign _0948_ = _0947_ | \mchip.index [6];
	assign _0949_ = _0948_ | \mchip.index [7];
	assign _0950_ = \mchip.index [11] & ~_0949_;
	assign _0951_ = _0744_ | \mchip.index [6];
	assign _0952_ = _0951_ | _1430_;
	assign _0953_ = \mchip.index [10] & ~_0952_;
	assign _0954_ = _0074_ | _1540_;
	assign _0956_ = _0954_ | _1430_;
	assign _0957_ = \mchip.index [8] & ~_0956_;
	assign _0958_ = _2655_ | _1430_;
	assign _0959_ = \mchip.index [11] & ~_0958_;
	assign _0960_ = _0176_ | _2161_;
	assign _0961_ = _0960_ | \mchip.index [6];
	assign _0962_ = _0961_ | _1430_;
	assign _0963_ = \mchip.index [8] & ~_0962_;
	assign _0964_ = _0604_ | \mchip.index [8];
	assign _0965_ = \mchip.index [9] & ~_0964_;
	assign _0967_ = _1930_ | _2030_;
	assign _0968_ = _0967_ | \mchip.index [6];
	assign _0969_ = _0968_ | _1430_;
	assign _0970_ = _0969_ | _2359_;
	assign _0971_ = _2271_ & ~_0970_;
	assign _0972_ = _0971_ | _0965_;
	assign _0973_ = _0972_ | _0963_;
	assign _0974_ = _0973_ | _0959_;
	assign _0975_ = _0974_ | _0957_;
	assign _0976_ = _0975_ | _0953_;
	assign _0978_ = _0976_ | _0950_;
	assign _0979_ = _0978_ | _0945_;
	assign _0980_ = _0979_ | _0942_;
	assign _0981_ = _0980_ | _0939_;
	assign _0982_ = _0981_ | _0936_;
	assign _0983_ = _0982_ | _0934_;
	assign _0984_ = _0983_ | _0931_;
	assign _0985_ = _0984_ | _0484_;
	assign _0986_ = _0985_ | _0480_;
	assign _0987_ = _0986_ | _0927_;
	assign _0989_ = _0987_ | _0924_;
	assign _0990_ = _0989_ | _0920_;
	assign _0991_ = _0990_ | _0918_;
	assign _0992_ = _0991_ | _0915_;
	assign _0993_ = _0992_ | _0912_;
	assign _0994_ = _0993_ | _0909_;
	assign _0995_ = _0994_ | _0907_;
	assign _0996_ = _0995_ | _0905_;
	assign _0997_ = _0996_ | _0903_;
	assign _0998_ = _0997_ | _0898_;
	assign _1000_ = _0998_ | _0892_;
	assign _1001_ = _1000_ | _0888_;
	assign _1002_ = _1001_ | _0886_;
	assign _1003_ = _1002_ | _0884_;
	assign _1004_ = _1003_ | _0880_;
	assign _1005_ = _1004_ | _0876_;
	assign _1006_ = _1005_ | _0872_;
	assign _1007_ = _1006_ | _0869_;
	assign _1008_ = _1007_ | _0441_;
	assign _1009_ = _1008_ | _0863_;
	assign _1011_ = _1009_ | _0862_;
	assign _1012_ = _1011_ | _0860_;
	assign _1013_ = _1012_ | _0859_;
	assign _1014_ = _1013_ | _0857_;
	assign _1015_ = _1014_ | _0852_;
	assign _1016_ = _1015_ | _0849_;
	assign _1017_ = _1016_ | _0846_;
	assign _1018_ = _1017_ | _0844_;
	assign _1019_ = _1018_ | _0842_;
	assign _1020_ = _1019_ | _0841_;
	assign _1022_ = _1020_ | _0839_;
	assign _1023_ = _1022_ | _0837_;
	assign _1024_ = _1023_ | _0833_;
	assign _1025_ = _1024_ | _0831_;
	assign _1026_ = _1025_ | _0415_;
	assign _1027_ = _1026_ | _0828_;
	assign _1028_ = _1027_ | _0826_;
	assign _1029_ = _1028_ | _1021_;
	assign _1030_ = _1029_ | _0824_;
	assign _1031_ = _1030_ | _2657_;
	assign _1033_ = _1031_ | _0821_;
	assign _1034_ = _1033_ | _0819_;
	assign _1035_ = _1034_ | _0817_;
	assign _1036_ = _1035_ | _0813_;
	assign _1037_ = _1036_ | _0808_;
	assign _1038_ = _1037_ | _0806_;
	assign _1039_ = _1038_ | _0804_;
	assign _1040_ = _1039_ | _0802_;
	assign _1041_ = _1040_ | _0797_;
	assign _1042_ = _1041_ | _0794_;
	assign _1044_ = _1042_ | _0789_;
	assign _1045_ = _1044_ | _0786_;
	assign _1046_ = _1045_ | _0784_;
	assign _1047_ = _1046_ | _0781_;
	assign _1048_ = _1047_ | _0777_;
	assign _1049_ = _1048_ | _0776_;
	assign _1050_ = _1049_ | _0389_;
	assign _1051_ = _1050_ | _0773_;
	assign _1052_ = _1051_ | _0771_;
	assign _1053_ = _1052_ | _0766_;
	assign _1055_ = _1053_ | _0765_;
	assign _1056_ = _1055_ | _0762_;
	assign _1057_ = _1056_ | _0760_;
	assign _1058_ = _1057_ | _0756_;
	assign _1059_ = _1058_ | _0755_;
	assign _1060_ = _1059_ | _0753_;
	assign _1061_ = _1060_ | _0750_;
	assign _1062_ = _1061_ | _0748_;
	assign _1063_ = _1062_ | _0742_;
	assign _1064_ = _1063_ | _0740_;
	assign _1066_ = _1064_ | _0737_;
	assign _1067_ = _1066_ | _0730_;
	assign _1068_ = _1067_ | _0727_;
	assign _1069_ = _1068_ | _0723_;
	assign _1070_ = _1069_ | _0718_;
	assign _1071_ = _1070_ | _0716_;
	assign _1072_ = _1071_ | _0712_;
	assign _1073_ = _1072_ | _0711_;
	assign _1074_ = _1073_ | _0708_;
	assign _1075_ = _1074_ | _0704_;
	assign _1077_ = _1075_ | _0700_;
	assign _1078_ = _1077_ | _0695_;
	assign _1079_ = _1078_ | _0692_;
	assign _1080_ = _1079_ | _0687_;
	assign _1081_ = _1080_ | _0684_;
	assign _1082_ = _1081_ | _0681_;
	assign _1083_ = _1082_ | _0677_;
	assign _1084_ = _1083_ | _0676_;
	assign _1085_ = _1084_ | _0226_;
	assign _1086_ = _1085_ | _0674_;
	assign _1088_ = _1086_ | _0672_;
	assign \mchip.val [2] = _1088_ | _0670_;
	assign _1089_ = _2025_ | _1430_;
	assign _1090_ = _1089_ | \mchip.index [9];
	assign _1091_ = _1931_ & ~_1090_;
	assign _1092_ = _1976_ | _2030_;
	assign _1093_ = _1092_ | _2161_;
	assign _1094_ = \mchip.index [6] & ~_1093_;
	assign _1095_ = _0074_ | _1430_;
	assign _1096_ = \mchip.index [11] & ~_1095_;
	assign _1099_ = _1942_ | _2030_;
	assign _1100_ = _1099_ | \mchip.index [6];
	assign _1101_ = _1100_ | \mchip.index [8];
	assign _1102_ = \mchip.index [9] & ~_1101_;
	assign _1103_ = _2029_ | \mchip.index [5];
	assign _1104_ = _1103_ | \mchip.index [6];
	assign _1105_ = _1104_ | \mchip.index [7];
	assign _1106_ = \mchip.index [11] & ~_1105_;
	assign _1107_ = _0492_ | \mchip.index [6];
	assign _1108_ = _1107_ | \mchip.index [7];
	assign _1110_ = \mchip.index [8] & ~_1108_;
	assign _1111_ = _0408_ | \mchip.index [5];
	assign _1112_ = _1111_ | \mchip.index [6];
	assign _1113_ = _1112_ | _1430_;
	assign _1114_ = \mchip.index [8] & ~_1113_;
	assign _1115_ = _2697_ | \mchip.index [8];
	assign _1116_ = \mchip.index [9] & ~_1115_;
	assign _1117_ = _2551_ | \mchip.index [5];
	assign _1118_ = _1117_ | _1540_;
	assign _1119_ = \mchip.index [11] & ~_1118_;
	assign _1121_ = _1931_ & ~_2450_;
	assign _1122_ = _0093_ | \mchip.index [7];
	assign _1123_ = _1122_ | _1319_;
	assign _1124_ = _1931_ & ~_1123_;
	assign _1125_ = _0370_ | \mchip.index [8];
	assign _1126_ = \mchip.index [9] & ~_1125_;
	assign _1127_ = \mchip.index [10] & ~_2448_;
	assign _1128_ = _1941_ | \mchip.index [8];
	assign _1129_ = \mchip.index [10] & ~_1128_;
	assign _1130_ = _2437_ | _1430_;
	assign _1132_ = _1130_ | _2359_;
	assign _1133_ = _1931_ & ~_1132_;
	assign _1134_ = _0370_ | \mchip.index [7];
	assign _1135_ = _1134_ | _1319_;
	assign _1136_ = _2271_ & ~_1135_;
	assign _1137_ = _0288_ | _2359_;
	assign _1138_ = _2271_ & ~_1137_;
	assign _1139_ = _2555_ | \mchip.index [5];
	assign _1140_ = _1139_ | _1540_;
	assign _1141_ = _1140_ | \mchip.index [7];
	assign _1143_ = \mchip.index [11] & ~_1141_;
	assign _1144_ = _2511_ | \mchip.index [7];
	assign _1145_ = _1144_ | _2359_;
	assign _1146_ = _1931_ & ~_1145_;
	assign _1147_ = _2026_ | _2359_;
	assign _1148_ = _1147_ | \mchip.index [9];
	assign _1149_ = \mchip.index [10] & ~_1148_;
	assign _1150_ = \mchip.index [11] & ~_0717_;
	assign _1151_ = _1979_ & ~\mchip.index [11];
	assign _1152_ = _2219_ | _1430_;
	assign _1154_ = _1152_ | \mchip.index [8];
	assign _1155_ = \mchip.index [10] & ~_1154_;
	assign _1156_ = _2392_ | \mchip.index [6];
	assign _1157_ = _1156_ | \mchip.index [7];
	assign _1158_ = \mchip.index [11] & ~_1157_;
	assign _1159_ = \mchip.index [10] & ~_0016_;
	assign _1160_ = _0725_ | \mchip.index [6];
	assign _1161_ = _1160_ | \mchip.index [7];
	assign _1162_ = \mchip.index [10] & ~_1161_;
	assign _1163_ = _2602_ | _1540_;
	assign _1165_ = _1163_ | \mchip.index [7];
	assign _1166_ = _1165_ | _2359_;
	assign _1167_ = _1166_ | _1319_;
	assign _1168_ = _1167_ | \mchip.index [10];
	assign _1169_ = _2271_ & ~_1168_;
	assign _1170_ = _1319_ & ~_2659_;
	assign _1171_ = \mchip.index [11] & ~_0354_;
	assign _1172_ = _2582_ | \mchip.index [8];
	assign _1173_ = _1172_ | \mchip.index [9];
	assign _1174_ = _2271_ & ~_1173_;
	assign _1176_ = \mchip.index [11] & ~_0227_;
	assign _1177_ = _2158_ | \mchip.index [5];
	assign _1178_ = _1177_ | _1540_;
	assign _1179_ = _1178_ | _1430_;
	assign _1180_ = _2359_ & ~_1179_;
	assign _1181_ = _0967_ | _1540_;
	assign _1182_ = _1181_ | _1430_;
	assign _1183_ = _2271_ & ~_1182_;
	assign _1184_ = _0544_ | _1430_;
	assign _1185_ = _1319_ & ~_1184_;
	assign _1187_ = _2026_ | _1430_;
	assign _1188_ = _1319_ & ~_1187_;
	assign _1189_ = _2279_ | \mchip.index [7];
	assign _1190_ = _1189_ | \mchip.index [9];
	assign _1191_ = \mchip.index [10] & ~_1190_;
	assign _1192_ = _2463_ | _1430_;
	assign _1193_ = _1319_ & ~_1192_;
	assign _1194_ = _2685_ | _1319_;
	assign _1195_ = _2271_ & ~_1194_;
	assign _1196_ = _0011_ | _1430_;
	assign _1198_ = _1196_ | \mchip.index [9];
	assign _1199_ = _1931_ & ~_1198_;
	assign _1200_ = _2557_ | \mchip.index [7];
	assign _1201_ = _2359_ & ~_1200_;
	assign _1202_ = \mchip.index [10] & ~_2439_;
	assign _1203_ = _1430_ & ~_0213_;
	assign _1204_ = _1818_ | \mchip.index [8];
	assign _1205_ = \mchip.index [10] & ~_1204_;
	assign _1206_ = _0412_ | \mchip.index [9];
	assign _1207_ = _1931_ & ~_1206_;
	assign _1210_ = _0812_ | \mchip.index [6];
	assign _1211_ = _1210_ | _1430_;
	assign _1212_ = _1211_ | \mchip.index [8];
	assign _1213_ = _1212_ | _1319_;
	assign _1214_ = _1213_ | \mchip.index [10];
	assign _1215_ = _2271_ & ~_1214_;
	assign _1216_ = \mchip.index [9] & ~_0254_;
	assign _1217_ = _0002_ | _1430_;
	assign _1218_ = _1217_ | _2359_;
	assign _1219_ = _1218_ | _1319_;
	assign _1221_ = _1219_ | _1931_;
	assign _1222_ = \mchip.index [11] & ~_1221_;
	assign _1223_ = _1927_ | _2030_;
	assign _1224_ = _1223_ | \mchip.index [7];
	assign _1225_ = _2359_ & ~_1224_;
	assign _1226_ = _2359_ & ~_0925_;
	assign _1227_ = _0092_ | \mchip.index [6];
	assign _1228_ = _1227_ | \mchip.index [7];
	assign _1229_ = _2359_ & ~_1228_;
	assign _1230_ = _2484_ | _2359_;
	assign _1232_ = _1230_ | _1319_;
	assign _1233_ = _1232_ | _1931_;
	assign _1234_ = \mchip.index [11] & ~_1233_;
	assign _1235_ = _1319_ & ~_0264_;
	assign _1236_ = _1319_ & ~_0425_;
	assign _1237_ = _0791_ | _2161_;
	assign _1238_ = _1237_ | \mchip.index [7];
	assign _1239_ = \mchip.index [11] & ~_1238_;
	assign _1240_ = _0782_ | \mchip.index [9];
	assign _1241_ = _1931_ & ~_1240_;
	assign _1243_ = _2512_ | \mchip.index [7];
	assign _1244_ = _1243_ | \mchip.index [8];
	assign _1245_ = _1244_ | \mchip.index [9];
	assign _1246_ = _1245_ | _1931_;
	assign _1247_ = _2271_ & ~_1246_;
	assign _1248_ = _0705_ | \mchip.index [8];
	assign _1249_ = \mchip.index [9] & ~_1248_;
	assign _1250_ = _1935_ | _2030_;
	assign _1251_ = _1250_ | _1540_;
	assign _1252_ = _1251_ | _1430_;
	assign _1254_ = \mchip.index [11] & ~_1252_;
	assign _1255_ = _0221_ | _1319_;
	assign _1256_ = _1931_ & ~_1255_;
	assign _1257_ = _2315_ | _2161_;
	assign _1258_ = \mchip.index [6] & ~_1257_;
	assign _1259_ = _0465_ | _1430_;
	assign _1260_ = \mchip.index [11] & ~_1259_;
	assign _1261_ = _2564_ | \mchip.index [6];
	assign _1262_ = _1319_ & ~_1261_;
	assign _1263_ = _0055_ | \mchip.index [4];
	assign _1265_ = _1263_ | \mchip.index [6];
	assign _1266_ = _1265_ | _1430_;
	assign _1267_ = _1266_ | _2359_;
	assign _1268_ = _2271_ & ~_1267_;
	assign _1269_ = _2525_ | \mchip.index [7];
	assign _1270_ = _2359_ & ~_1269_;
	assign _1271_ = _0944_ | \mchip.index [4];
	assign _1272_ = _1271_ | _1540_;
	assign _1273_ = _1272_ | \mchip.index [7];
	assign _1274_ = _1273_ | \mchip.index [9];
	assign _1276_ = \mchip.index [10] & ~_1274_;
	assign _1277_ = _0308_ | \mchip.index [4];
	assign _1278_ = _1277_ | _1540_;
	assign _1279_ = _1278_ | \mchip.index [7];
	assign _1280_ = _2359_ & ~_1279_;
	assign _1281_ = _2555_ | _2161_;
	assign _1282_ = _1281_ | \mchip.index [6];
	assign _1283_ = _1430_ & ~_1282_;
	assign _1284_ = _0889_ | _2030_;
	assign _1285_ = _1284_ | \mchip.index [7];
	assign _1287_ = \mchip.index [10] & ~_1285_;
	assign _1288_ = _2496_ | \mchip.index [5];
	assign _1289_ = _1288_ | \mchip.index [6];
	assign _1290_ = _1289_ | \mchip.index [7];
	assign _1291_ = \mchip.index [11] & ~_1290_;
	assign _1292_ = _0330_ | \mchip.index [6];
	assign _1293_ = _1292_ | _1430_;
	assign _1294_ = \mchip.index [11] & ~_1293_;
	assign _1295_ = _2551_ | _1430_;
	assign _1296_ = \mchip.index [11] & ~_1295_;
	assign _1298_ = _2230_ | _2161_;
	assign _1299_ = \mchip.index [6] & ~_1298_;
	assign _1300_ = _0758_ | \mchip.index [7];
	assign _1301_ = _1300_ | _1319_;
	assign _1302_ = _2271_ & ~_1301_;
	assign _1303_ = _2611_ | _2359_;
	assign _1304_ = _1319_ & ~_1303_;
	assign _1305_ = _0375_ | _2161_;
	assign _1306_ = \mchip.index [7] & ~_1305_;
	assign _1307_ = _0533_ | \mchip.index [7];
	assign _1309_ = \mchip.index [11] & ~_1307_;
	assign _1310_ = \mchip.index [11] & ~_2454_;
	assign _1311_ = _0860_ & ~_1540_;
	assign _1312_ = \mchip.index [9] & ~_2493_;
	assign _1313_ = _2611_ | _1540_;
	assign _1314_ = _1313_ | _1430_;
	assign _1315_ = _2359_ & ~_1314_;
	assign _1316_ = _0065_ | _1540_;
	assign _1317_ = _1316_ | \mchip.index [8];
	assign _1318_ = _1931_ & ~_1317_;
	assign _1321_ = _1904_ | _2161_;
	assign _1322_ = _1540_ & ~_1321_;
	assign _1323_ = _1092_ | _1540_;
	assign _1324_ = _1323_ | _2359_;
	assign _1325_ = _1324_ | _1319_;
	assign _1326_ = _1931_ & ~_1325_;
	assign _1327_ = _1935_ | _1540_;
	assign _1328_ = _1327_ | \mchip.index [8];
	assign _1329_ = \mchip.index [9] & ~_1328_;
	assign _1330_ = _2459_ | \mchip.index [6];
	assign _1332_ = _1931_ & ~_1330_;
	assign _1333_ = _1253_ | \mchip.index [6];
	assign _1334_ = _1333_ | \mchip.index [7];
	assign _1335_ = _1931_ & ~_1334_;
	assign _1336_ = _2458_ | _1430_;
	assign _1337_ = _1336_ | _2359_;
	assign _1338_ = _1931_ & ~_1337_;
	assign _1339_ = _0081_ | \mchip.index [5];
	assign _1340_ = _1339_ | \mchip.index [7];
	assign _1341_ = \mchip.index [8] & ~_1340_;
	assign _1343_ = _2492_ | \mchip.index [7];
	assign _1344_ = \mchip.index [11] & ~_1343_;
	assign _1345_ = _2541_ | \mchip.index [6];
	assign _1346_ = _1345_ | _1430_;
	assign _1347_ = \mchip.index [10] & ~_1346_;
	assign _1348_ = _0070_ | _1540_;
	assign _1349_ = _1348_ | \mchip.index [7];
	assign _1350_ = \mchip.index [10] & ~_1349_;
	assign _1351_ = _2499_ | \mchip.index [5];
	assign _1352_ = _1351_ | _1430_;
	assign _1354_ = \mchip.index [11] & ~_1352_;
	assign _1355_ = _1982_ | \mchip.index [7];
	assign _1356_ = \mchip.index [9] & ~_1355_;
	assign _1357_ = _0055_ | _1540_;
	assign _1358_ = _1357_ | \mchip.index [7];
	assign _1359_ = _1358_ | \mchip.index [9];
	assign _1360_ = \mchip.index [10] & ~_1359_;
	assign _1361_ = _1360_ | _1356_;
	assign _1362_ = _1361_ | _1354_;
	assign _1363_ = _1362_ | _1350_;
	assign _1365_ = _1363_ | _1347_;
	assign _1366_ = _1365_ | _1344_;
	assign _1367_ = _1366_ | _1341_;
	assign _1368_ = _1367_ | _0957_;
	assign _1369_ = _1368_ | _1338_;
	assign _1370_ = _1369_ | _1335_;
	assign _1371_ = _1370_ | _1332_;
	assign _1372_ = _1371_ | _1329_;
	assign _1373_ = _1372_ | _1326_;
	assign _1374_ = _1373_ | _1322_;
	assign _1376_ = _1374_ | _1318_;
	assign _1377_ = _1376_ | _0491_;
	assign _1378_ = _1377_ | _1315_;
	assign _1379_ = _1378_ | _1312_;
	assign _1380_ = _1379_ | _1311_;
	assign _1381_ = _1380_ | _1310_;
	assign _1382_ = _1381_ | _1309_;
	assign _1383_ = _1382_ | _0396_;
	assign _1384_ = _1383_ | _1306_;
	assign _1385_ = _1384_ | _1304_;
	assign _1387_ = _1385_ | _1302_;
	assign _1388_ = _1387_ | _1299_;
	assign _1389_ = _1388_ | _1296_;
	assign _1390_ = _1389_ | _1294_;
	assign _1391_ = _1390_ | _1291_;
	assign _1392_ = _1391_ | _0459_;
	assign _1393_ = _1392_ | _1287_;
	assign _1394_ = _1393_ | _1283_;
	assign _1395_ = _1394_ | _1280_;
	assign _1396_ = _1395_ | _1276_;
	assign _1398_ = _1396_ | _1270_;
	assign _1399_ = _1398_ | _1268_;
	assign _1400_ = _1399_ | _1262_;
	assign _1401_ = _1400_ | _1260_;
	assign _1402_ = _1401_ | _1258_;
	assign _1403_ = _1402_ | _1256_;
	assign _1404_ = _1403_ | _1254_;
	assign _1405_ = _1404_ | _1249_;
	assign _1406_ = _1405_ | _1247_;
	assign _1407_ = _1406_ | _1241_;
	assign _1409_ = _1407_ | _1239_;
	assign _1410_ = _1409_ | _1236_;
	assign _1411_ = _1410_ | _1235_;
	assign _1412_ = _1411_ | _1234_;
	assign _1413_ = _1412_ | _1229_;
	assign _1414_ = _1413_ | _1226_;
	assign _1415_ = _1414_ | _1225_;
	assign _1416_ = _1415_ | _1222_;
	assign _1417_ = _1416_ | _1216_;
	assign _1418_ = _1417_ | _1215_;
	assign _1420_ = _1418_ | _0821_;
	assign _1421_ = _1420_ | _1207_;
	assign _1422_ = _1421_ | _1205_;
	assign _1423_ = _1422_ | _1203_;
	assign _1424_ = _1423_ | _1202_;
	assign _1425_ = _1424_ | _1201_;
	assign _1426_ = _1425_ | _1199_;
	assign _1427_ = _1426_ | _1195_;
	assign _1428_ = _1427_ | _1193_;
	assign _1429_ = _1428_ | _1191_;
	assign _1432_ = _1429_ | _1188_;
	assign _1433_ = _1432_ | _1185_;
	assign _1434_ = _1433_ | _1183_;
	assign _1435_ = _1434_ | _1180_;
	assign _1436_ = _1435_ | _1176_;
	assign _1437_ = _1436_ | _1174_;
	assign _1438_ = _1437_ | _0342_;
	assign _1439_ = _1438_ | _1171_;
	assign _1440_ = _1439_ | _1170_;
	assign _1441_ = _1440_ | _1169_;
	assign _1443_ = _1441_ | _1162_;
	assign _1444_ = _1443_ | _1159_;
	assign _1445_ = _1444_ | _1158_;
	assign _1446_ = _1445_ | _1155_;
	assign _1447_ = _1446_ | _1151_;
	assign _1448_ = _1447_ | _1150_;
	assign _1449_ = _1448_ | _1149_;
	assign _1450_ = _1449_ | _1146_;
	assign _1451_ = _1450_ | _1143_;
	assign _1452_ = _1451_ | _1138_;
	assign _1454_ = _1452_ | _1136_;
	assign _1455_ = _1454_ | _1133_;
	assign _1456_ = _1455_ | _1129_;
	assign _1457_ = _1456_ | _1127_;
	assign _1458_ = _1457_ | _1126_;
	assign _1459_ = _1458_ | _1124_;
	assign _1460_ = _1459_ | _1121_;
	assign _1461_ = _1460_ | _1119_;
	assign _1462_ = _1461_ | _1116_;
	assign _1463_ = _1462_ | _1114_;
	assign _1465_ = _1463_ | _1110_;
	assign _1466_ = _1465_ | _1106_;
	assign _1467_ = _1466_ | _1102_;
	assign _1468_ = _1467_ | _1096_;
	assign _1469_ = _1468_ | _1094_;
	assign \mchip.val [1] = _1469_ | _1091_;
	assign _1470_ = _2696_ | \mchip.index [6];
	assign _1471_ = _1470_ | \mchip.index [7];
	assign _1472_ = _2359_ & ~_1471_;
	assign _1473_ = _1319_ & ~_2443_;
	assign _1475_ = _2696_ | \mchip.index [9];
	assign _1476_ = _1931_ & ~_1475_;
	assign _1477_ = _0055_ | _2161_;
	assign _1478_ = \mchip.index [7] & ~_1477_;
	assign _1479_ = _1984_ | _2161_;
	assign _1480_ = _1479_ | _1430_;
	assign _1481_ = \mchip.index [8] & ~_1480_;
	assign _1482_ = _1931_ & ~_2118_;
	assign _1483_ = _1263_ | _1430_;
	assign _1484_ = _1483_ | _2359_;
	assign _1486_ = _1931_ & ~_1484_;
	assign _1487_ = _0893_ | \mchip.index [7];
	assign _1488_ = _1487_ | _2359_;
	assign _1489_ = _1488_ | _1319_;
	assign _1490_ = _1489_ | _1931_;
	assign _1491_ = \mchip.index [11] & ~_1490_;
	assign _1492_ = _1319_ & ~_0205_;
	assign _1493_ = _1851_ | \mchip.index [4];
	assign _1494_ = _1493_ | \mchip.index [5];
	assign _1495_ = _1494_ | \mchip.index [6];
	assign _1497_ = _1495_ | \mchip.index [7];
	assign _1498_ = \mchip.index [11] & ~_1497_;
	assign _1499_ = _1976_ | _1540_;
	assign _1500_ = _1499_ | \mchip.index [7];
	assign _1501_ = _1500_ | _1319_;
	assign _1502_ = _1931_ & ~_1501_;
	assign _1503_ = \mchip.index [9] & ~_0238_;
	assign _1504_ = _0282_ | \mchip.index [7];
	assign _1505_ = _2359_ & ~_1504_;
	assign _1506_ = _0682_ | _2359_;
	assign _1508_ = _1931_ & ~_1506_;
	assign _1509_ = _1507_ | \mchip.index [5];
	assign _1510_ = _1509_ | \mchip.index [6];
	assign _1511_ = _1510_ | \mchip.index [7];
	assign _1512_ = \mchip.index [11] & ~_1511_;
	assign _1513_ = _2271_ & ~_1285_;
	assign _1514_ = _0375_ | \mchip.index [5];
	assign _1515_ = _1514_ | _1540_;
	assign _1516_ = _1515_ | \mchip.index [7];
	assign _1517_ = \mchip.index [9] & ~_1516_;
	assign _1519_ = _2611_ | \mchip.index [6];
	assign _1520_ = _1519_ | \mchip.index [8];
	assign _1521_ = \mchip.index [10] & ~_1520_;
	assign _1522_ = _2655_ | \mchip.index [8];
	assign _1523_ = _1931_ & ~_1522_;
	assign _1524_ = _2445_ | _1540_;
	assign _1525_ = _1430_ & ~_1524_;
	assign _1526_ = _0885_ | \mchip.index [7];
	assign _1527_ = \mchip.index [8] & ~_1526_;
	assign _1528_ = _2642_ | \mchip.index [6];
	assign _1530_ = _1528_ | _1430_;
	assign _1531_ = \mchip.index [11] & ~_1530_;
	assign _1532_ = \mchip.index [6] & ~_1321_;
	assign _1533_ = _2516_ | _1540_;
	assign _1534_ = _1533_ | _1430_;
	assign _1535_ = \mchip.index [9] & ~_1534_;
	assign _1536_ = _1043_ | _1430_;
	assign _1537_ = _1536_ | \mchip.index [9];
	assign _1538_ = _1931_ & ~_1537_;
	assign _1539_ = _1936_ | _1540_;
	assign _1542_ = _1539_ | _1430_;
	assign _1543_ = \mchip.index [11] & ~_1542_;
	assign _1544_ = _1552_ | \mchip.index [5];
	assign _1545_ = _1544_ | \mchip.index [6];
	assign _1546_ = _1545_ | _2359_;
	assign _1547_ = \mchip.index [10] & ~_1546_;
	assign _1548_ = _1186_ | _1540_;
	assign _1549_ = _1548_ | _1430_;
	assign _1550_ = _1549_ | _2359_;
	assign _1551_ = _1931_ & ~_1550_;
	assign _1553_ = _0096_ | \mchip.index [5];
	assign _1554_ = _1553_ | _1540_;
	assign _1555_ = \mchip.index [11] & ~_1554_;
	assign _1556_ = _2271_ & ~_0717_;
	assign _1557_ = _1618_ | _1540_;
	assign _1558_ = _1557_ | \mchip.index [7];
	assign _1559_ = _1558_ | _2359_;
	assign _1560_ = _1559_ | _1319_;
	assign _1561_ = _1560_ | \mchip.index [10];
	assign _1562_ = _2271_ & ~_1561_;
	assign _1564_ = _0853_ | _2359_;
	assign _1565_ = \mchip.index [10] & ~_1564_;
	assign _1566_ = _1277_ | \mchip.index [6];
	assign _1567_ = _1566_ | _1430_;
	assign _1568_ = _1567_ | \mchip.index [8];
	assign _1569_ = \mchip.index [10] & ~_1568_;
	assign _1570_ = _0031_ | _1430_;
	assign _1571_ = _1570_ | \mchip.index [9];
	assign _1572_ = _1931_ & ~_1571_;
	assign _1573_ = _1984_ | \mchip.index [6];
	assign _1575_ = _1573_ | _1430_;
	assign _1576_ = _1575_ | \mchip.index [8];
	assign _1577_ = _1576_ | \mchip.index [9];
	assign _1578_ = _1577_ | \mchip.index [10];
	assign _1579_ = _2271_ & ~_1578_;
	assign _1580_ = _0460_ | _2359_;
	assign _1581_ = _1931_ & ~_1580_;
	assign _1582_ = _2175_ & ~\mchip.index [11];
	assign _1583_ = _0763_ | _1540_;
	assign _1584_ = _1583_ | \mchip.index [7];
	assign _1586_ = _1931_ & ~_1584_;
	assign _1587_ = _1087_ | _2161_;
	assign _1588_ = \mchip.index [7] & ~_1587_;
	assign _1589_ = _1607_ | _2030_;
	assign _1590_ = _1589_ | _2161_;
	assign _1591_ = _1590_ | \mchip.index [6];
	assign _1592_ = _1430_ & ~_1591_;
	assign _1593_ = _0648_ | _2161_;
	assign _1594_ = _1593_ | \mchip.index [6];
	assign _1595_ = _1430_ & ~_1594_;
	assign _1597_ = _0015_ | \mchip.index [8];
	assign _1598_ = \mchip.index [10] & ~_1597_;
	assign _1599_ = _2676_ | \mchip.index [5];
	assign _1600_ = _1599_ | _1540_;
	assign _1601_ = _1600_ | \mchip.index [8];
	assign _1602_ = _1601_ | \mchip.index [9];
	assign _1603_ = _1602_ | _1931_;
	assign _1604_ = _2271_ & ~_1603_;
	assign _1605_ = _0889_ | \mchip.index [8];
	assign _1606_ = _1931_ & ~_1605_;
	assign _1608_ = _1947_ | _2359_;
	assign _1609_ = _1608_ | _1319_;
	assign _1610_ = _2271_ & ~_1609_;
	assign _1611_ = _0014_ | _2161_;
	assign _1612_ = _1540_ & ~_1611_;
	assign _1613_ = _0731_ | _2030_;
	assign _1614_ = _1613_ | \mchip.index [5];
	assign _1615_ = _1614_ | _1540_;
	assign _1616_ = _1615_ | \mchip.index [7];
	assign _1617_ = \mchip.index [11] & ~_1616_;
	assign _1619_ = _2501_ | _1540_;
	assign _1620_ = _1619_ | _1430_;
	assign _1621_ = _1620_ | \mchip.index [8];
	assign _1622_ = _1621_ | _1319_;
	assign _1623_ = _1622_ | \mchip.index [10];
	assign _1624_ = _2271_ & ~_1623_;
	assign _1625_ = _2315_ | \mchip.index [4];
	assign _1626_ = _1625_ | _1540_;
	assign _1627_ = _1626_ | _2359_;
	assign _1628_ = _1627_ | _1319_;
	assign _1630_ = _2271_ & ~_1628_;
	assign _1631_ = _2501_ | \mchip.index [6];
	assign _1632_ = _1631_ | \mchip.index [7];
	assign _1633_ = _1632_ | _2359_;
	assign _1634_ = _1633_ | \mchip.index [9];
	assign _1635_ = _1634_ | _1931_;
	assign _1636_ = _2271_ & ~_1635_;
	assign _1637_ = _0002_ | \mchip.index [6];
	assign _1638_ = _1637_ | _1430_;
	assign _1639_ = _1638_ | \mchip.index [8];
	assign _1641_ = _1639_ | \mchip.index [9];
	assign _1642_ = _1641_ | _1931_;
	assign _1643_ = _2271_ & ~_1642_;
	assign _1644_ = _1342_ | _2030_;
	assign _1645_ = _1644_ | \mchip.index [7];
	assign _1646_ = _1931_ & ~_1645_;
	assign _1647_ = _1540_ & ~_1298_;
	assign _1648_ = _0308_ | \mchip.index [7];
	assign _1649_ = _1648_ | \mchip.index [8];
	assign _1650_ = _1931_ & ~_1649_;
	assign _1653_ = _2604_ | _1319_;
	assign _1654_ = _1653_ | \mchip.index [10];
	assign _1655_ = _2271_ & ~_1654_;
	assign _1656_ = _0472_ | _1540_;
	assign _1657_ = _1656_ | \mchip.index [8];
	assign _1658_ = \mchip.index [9] & ~_1657_;
	assign _1659_ = _0009_ | _2161_;
	assign _1660_ = \mchip.index [6] & ~_1659_;
	assign _1661_ = _0366_ | _1540_;
	assign _1662_ = _1661_ | _1430_;
	assign _1664_ = _1319_ & ~_1662_;
	assign _1665_ = _0347_ | _1430_;
	assign _1666_ = \mchip.index [10] & ~_1665_;
	assign _1667_ = _2499_ | \mchip.index [8];
	assign _1668_ = \mchip.index [9] & ~_1667_;
	assign _1669_ = _0691_ | \mchip.index [5];
	assign _1670_ = _1669_ | \mchip.index [6];
	assign _1671_ = _1670_ | \mchip.index [7];
	assign _1672_ = _1931_ & ~_1671_;
	assign _1673_ = _1931_ & ~_0081_;
	assign _1675_ = _1931_ & ~_1200_;
	assign _1676_ = _1284_ | _1540_;
	assign _1677_ = \mchip.index [10] & ~_1676_;
	assign _1678_ = \mchip.index [10] & ~_0495_;
	assign _1679_ = _2085_ | \mchip.index [8];
	assign _1680_ = \mchip.index [9] & ~_1679_;
	assign _1681_ = _1292_ | \mchip.index [8];
	assign _1682_ = \mchip.index [10] & ~_1681_;
	assign _1683_ = _2192_ & ~\mchip.index [10];
	assign _1684_ = _1662_ | _2359_;
	assign _1686_ = _2271_ & ~_1684_;
	assign _1687_ = _0532_ | \mchip.index [6];
	assign _1688_ = _1687_ | _1430_;
	assign _1689_ = _1688_ | _1319_;
	assign _1690_ = _2271_ & ~_1689_;
	assign _1691_ = _0678_ | _2359_;
	assign _1692_ = _2271_ & ~_1691_;
	assign _1693_ = _2002_ | _2359_;
	assign _1694_ = _1319_ & ~_1693_;
	assign _1695_ = _2231_ | \mchip.index [7];
	assign _1697_ = _2359_ & ~_1695_;
	assign _1698_ = _0472_ | _2030_;
	assign _1699_ = _1698_ | \mchip.index [6];
	assign _1700_ = _1699_ | _1430_;
	assign _1701_ = \mchip.index [11] & ~_1700_;
	assign _1702_ = _0809_ | \mchip.index [9];
	assign _1703_ = _1931_ & ~_1702_;
	assign _1704_ = _0728_ | _2359_;
	assign _1705_ = \mchip.index [9] & ~_1704_;
	assign _1706_ = _0705_ | \mchip.index [6];
	assign _1708_ = _1706_ | \mchip.index [7];
	assign _1709_ = _2359_ & ~_1708_;
	assign _1710_ = _2513_ | \mchip.index [6];
	assign _1711_ = \mchip.index [11] & ~_1710_;
	assign _1712_ = _2271_ & ~_0851_;
	assign _1713_ = _2230_ | _1540_;
	assign _1714_ = _1713_ | \mchip.index [8];
	assign _1715_ = \mchip.index [9] & ~_1714_;
	assign _1716_ = _2253_ | \mchip.index [6];
	assign _1717_ = _1716_ | \mchip.index [7];
	assign _1719_ = _1319_ & ~_1717_;
	assign _1720_ = _0439_ | _1540_;
	assign _1721_ = _1720_ | _2359_;
	assign _1722_ = _1319_ & ~_1721_;
	assign _1723_ = \mchip.index [10] & ~_0626_;
	assign _1724_ = \mchip.index [8] & ~_1295_;
	assign _1725_ = _0967_ | \mchip.index [5];
	assign _1726_ = _1725_ | \mchip.index [6];
	assign _1727_ = \mchip.index [11] & ~_1726_;
	assign _1728_ = _1575_ | _2359_;
	assign _1730_ = _1728_ | _1319_;
	assign _1731_ = _1730_ | _1931_;
	assign _1732_ = \mchip.index [11] & ~_1731_;
	assign _1733_ = _1186_ | _2161_;
	assign _1734_ = \mchip.index [6] & ~_1733_;
	assign _1735_ = _1851_ | _1430_;
	assign _1736_ = _1735_ | _2359_;
	assign _1737_ = _1931_ & ~_1736_;
	assign _1738_ = _1319_ & ~_0038_;
	assign _1739_ = _0099_ | _2161_;
	assign _1741_ = _1430_ & ~_1739_;
	assign _1742_ = \mchip.index [7] & ~_0468_;
	assign _1743_ = _1986_ | _1540_;
	assign _1744_ = _1743_ | _2359_;
	assign _1745_ = _1319_ & ~_1744_;
	assign _1746_ = _2516_ | _1430_;
	assign _1747_ = _1746_ | \mchip.index [9];
	assign _1748_ = _1931_ & ~_1747_;
	assign _1749_ = _0782_ | \mchip.index [8];
	assign _1750_ = \mchip.index [10] & ~_1749_;
	assign _1752_ = _2231_ | _1430_;
	assign _1753_ = \mchip.index [11] & ~_1752_;
	assign _1754_ = _2537_ | \mchip.index [8];
	assign _1755_ = \mchip.index [9] & ~_1754_;
	assign _1756_ = _2325_ | \mchip.index [6];
	assign _1757_ = _1756_ | \mchip.index [7];
	assign _1758_ = _1931_ & ~_1757_;
	assign _1759_ = _2208_ | _1540_;
	assign _1760_ = _1759_ | _1430_;
	assign _1761_ = _2271_ & ~_1760_;
	assign _1764_ = \mchip.index [11] & ~_0052_;
	assign _1765_ = _2200_ | _2161_;
	assign _1766_ = _1765_ | \mchip.index [6];
	assign _1767_ = _1766_ | \mchip.index [7];
	assign _1768_ = \mchip.index [10] & ~_1767_;
	assign _1769_ = _2491_ | _1430_;
	assign _1770_ = \mchip.index [10] & ~_1769_;
	assign _1771_ = _0767_ | _1430_;
	assign _1772_ = \mchip.index [11] & ~_1771_;
	assign _1773_ = _1464_ | _2161_;
	assign _1775_ = \mchip.index [7] & ~_1773_;
	assign _1776_ = _0033_ | _1931_;
	assign _1777_ = _2271_ & ~_1776_;
	assign _1778_ = _1777_ | _1775_;
	assign _1779_ = _1778_ | _1772_;
	assign _1780_ = _1779_ | _1770_;
	assign _1781_ = _1780_ | _1768_;
	assign _1782_ = _1781_ | _1764_;
	assign _1783_ = _1782_ | _1761_;
	assign _1784_ = _1783_ | _1758_;
	assign _1786_ = _1784_ | _1755_;
	assign _1787_ = _1786_ | _1753_;
	assign _1788_ = _1787_ | _1750_;
	assign _1789_ = _1788_ | _1748_;
	assign _1790_ = _1789_ | _1745_;
	assign _1791_ = _1790_ | _1742_;
	assign _1792_ = _1791_ | _1741_;
	assign _1793_ = _1792_ | _1738_;
	assign _1794_ = _1793_ | _0502_;
	assign _1795_ = _1794_ | _0086_;
	assign _1797_ = _1795_ | _1737_;
	assign _1798_ = _1797_ | _1734_;
	assign _1799_ = _1798_ | _0484_;
	assign _1800_ = _1799_ | _1732_;
	assign _1801_ = _1800_ | _1727_;
	assign _1802_ = _1801_ | _1724_;
	assign _1803_ = _1802_ | _1723_;
	assign _1804_ = _1803_ | _1722_;
	assign _1805_ = _1804_ | _1719_;
	assign _1806_ = _1805_ | _1715_;
	assign _1808_ = _1806_ | _1712_;
	assign _1809_ = _1808_ | _1711_;
	assign _1810_ = _1809_ | _1709_;
	assign _1811_ = _1810_ | _1705_;
	assign _1812_ = _1811_ | _1703_;
	assign _1813_ = _1812_ | _1701_;
	assign _1814_ = _1813_ | _0445_;
	assign _1815_ = _1814_ | _1697_;
	assign _1816_ = _1815_ | _1694_;
	assign _1817_ = _1816_ | _1692_;
	assign _1819_ = _1817_ | _1690_;
	assign _1820_ = _1819_ | _1686_;
	assign _1821_ = _1820_ | _1683_;
	assign _1822_ = _1821_ | _1682_;
	assign _1823_ = _1822_ | _0839_;
	assign _1824_ = _1823_ | _1680_;
	assign _1825_ = _1824_ | _1678_;
	assign _1826_ = _1825_ | _1677_;
	assign _1827_ = _1826_ | _1675_;
	assign _1828_ = _1827_ | _1673_;
	assign _1830_ = _1828_ | _1672_;
	assign _1831_ = _1830_ | _1668_;
	assign _1832_ = _1831_ | _1666_;
	assign _1833_ = _1832_ | _1664_;
	assign _1834_ = _1833_ | _1660_;
	assign _1835_ = _1834_ | _1658_;
	assign _1836_ = _1835_ | _0977_;
	assign _1837_ = _1836_ | _1655_;
	assign _1838_ = _1837_ | _1650_;
	assign _1839_ = _1838_ | _1647_;
	assign _1841_ = _1839_ | _1646_;
	assign _1842_ = _1841_ | _1643_;
	assign _1843_ = _1842_ | _1636_;
	assign _1844_ = _1843_ | _1630_;
	assign _1845_ = _1844_ | _1624_;
	assign _1846_ = _1845_ | _1617_;
	assign _1847_ = _1846_ | _0802_;
	assign _1848_ = _1847_ | _1612_;
	assign _1849_ = _1848_ | _1610_;
	assign _1850_ = _1849_ | _0369_;
	assign _1852_ = _1850_ | _1606_;
	assign _1853_ = _1852_ | _1604_;
	assign _1854_ = _1853_ | _1598_;
	assign _1855_ = _1854_ | _1595_;
	assign _1856_ = _1855_ | _1592_;
	assign _1857_ = _1856_ | _1588_;
	assign _1858_ = _1857_ | _1586_;
	assign _1859_ = _1858_ | _1582_;
	assign _1860_ = _1859_ | _1581_;
	assign _1861_ = _1860_ | _1579_;
	assign _1863_ = _1861_ | _1572_;
	assign _1864_ = _1863_ | _1569_;
	assign _1865_ = _1864_ | _1565_;
	assign _1866_ = _1865_ | _1562_;
	assign _1867_ = _1866_ | _1556_;
	assign _1868_ = _1867_ | _1555_;
	assign _1869_ = _1868_ | _1551_;
	assign _1870_ = _1869_ | _1547_;
	assign _1871_ = _1870_ | _1543_;
	assign _1872_ = _1871_ | _1538_;
	assign _1875_ = _1872_ | _1535_;
	assign _1876_ = _1875_ | _1532_;
	assign _1877_ = _1876_ | _1531_;
	assign _1878_ = _1877_ | _1527_;
	assign _1879_ = _1878_ | _1525_;
	assign _1880_ = _1879_ | _1523_;
	assign _1881_ = _1880_ | _1129_;
	assign _1882_ = _1881_ | _1521_;
	assign _1883_ = _1882_ | _1517_;
	assign _1884_ = _1883_ | _1513_;
	assign _1886_ = _1884_ | _1512_;
	assign _1887_ = _1886_ | _1508_;
	assign _1888_ = _1887_ | _1505_;
	assign _1889_ = _1888_ | _1503_;
	assign _1890_ = _1889_ | _1502_;
	assign _1891_ = _1890_ | _1498_;
	assign _1892_ = _1891_ | _1492_;
	assign _1893_ = _1892_ | _1491_;
	assign _1894_ = _1893_ | _1486_;
	assign _1895_ = _1894_ | _1482_;
	assign _1897_ = _1895_ | _1481_;
	assign _1898_ = _1897_ | _1478_;
	assign _1899_ = _1898_ | _1476_;
	assign _1900_ = _1899_ | _1473_;
	assign _1901_ = _1900_ | _1472_;
	assign \mchip.val [0] = _1901_ | _0670_;
	always @(posedge io_in[12]) \mchip.index [0] <= io_in[0];
	always @(posedge io_in[12]) \mchip.index [1] <= io_in[1];
	always @(posedge io_in[12]) \mchip.index [2] <= io_in[2];
	always @(posedge io_in[12]) \mchip.index [3] <= io_in[3];
	always @(posedge io_in[12]) \mchip.index [4] <= io_in[4];
	always @(posedge io_in[12]) \mchip.index [5] <= io_in[5];
	always @(posedge io_in[12]) \mchip.index [6] <= io_in[6];
	always @(posedge io_in[12]) \mchip.index [7] <= io_in[7];
	always @(posedge io_in[12]) \mchip.index [8] <= io_in[8];
	always @(posedge io_in[12]) \mchip.index [9] <= io_in[9];
	always @(posedge io_in[12]) \mchip.index [10] <= io_in[10];
	always @(posedge io_in[12]) \mchip.index [11] <= io_in[11];
	reg \mchip.io_out_reg[0] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[0]  <= \mchip.val [0];
	assign \mchip.io_out [0] = \mchip.io_out_reg[0] ;
	reg \mchip.io_out_reg[1] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[1]  <= \mchip.val [1];
	assign \mchip.io_out [1] = \mchip.io_out_reg[1] ;
	reg \mchip.io_out_reg[2] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[2]  <= \mchip.val [2];
	assign \mchip.io_out [2] = \mchip.io_out_reg[2] ;
	reg \mchip.io_out_reg[3] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[3]  <= \mchip.val [3];
	assign \mchip.io_out [3] = \mchip.io_out_reg[3] ;
	reg \mchip.io_out_reg[4] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[4]  <= \mchip.val [4];
	assign \mchip.io_out [4] = \mchip.io_out_reg[4] ;
	reg \mchip.io_out_reg[5] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[5]  <= \mchip.val [5];
	assign \mchip.io_out [5] = \mchip.io_out_reg[5] ;
	reg \mchip.io_out_reg[6] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[6]  <= \mchip.val [6];
	assign \mchip.io_out [6] = \mchip.io_out_reg[6] ;
	assign io_out = {7'h00, \mchip.io_out [6:0]};
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out [11:7] = 5'h00;
	assign \mchip.reset  = io_in[13];
	assign \mchip.val [7] = 1'h0;
endmodule
module d06_demo_vgapong (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire _2025_;
	wire _2026_;
	wire _2027_;
	wire _2028_;
	wire _2029_;
	wire _2030_;
	wire _2031_;
	wire _2032_;
	wire _2033_;
	wire _2034_;
	wire _2035_;
	wire _2036_;
	wire _2037_;
	wire _2038_;
	wire _2039_;
	wire _2040_;
	wire _2041_;
	wire _2042_;
	wire _2043_;
	wire _2044_;
	wire _2045_;
	wire _2046_;
	wire _2047_;
	wire _2048_;
	wire _2049_;
	wire _2050_;
	wire _2051_;
	wire _2052_;
	wire _2053_;
	wire _2054_;
	wire _2055_;
	wire _2056_;
	wire _2057_;
	wire _2058_;
	wire _2059_;
	wire _2060_;
	wire _2061_;
	wire _2062_;
	wire _2063_;
	wire _2064_;
	wire _2065_;
	wire _2066_;
	wire _2067_;
	wire _2068_;
	wire _2069_;
	wire _2070_;
	wire _2071_;
	wire _2072_;
	wire _2073_;
	wire _2074_;
	wire _2075_;
	wire _2076_;
	wire _2077_;
	wire _2078_;
	wire _2079_;
	wire _2080_;
	wire _2081_;
	wire _2082_;
	wire _2083_;
	wire _2084_;
	wire _2085_;
	wire _2086_;
	wire _2087_;
	wire _2088_;
	wire _2089_;
	wire _2090_;
	wire _2091_;
	wire _2092_;
	wire _2093_;
	wire _2094_;
	wire _2095_;
	wire _2096_;
	wire _2097_;
	wire _2098_;
	wire _2099_;
	wire _2100_;
	wire _2101_;
	wire _2102_;
	wire _2103_;
	wire _2104_;
	wire _2105_;
	wire _2106_;
	wire _2107_;
	wire _2108_;
	wire _2109_;
	wire _2110_;
	wire _2111_;
	wire _2112_;
	wire _2113_;
	wire _2114_;
	wire _2115_;
	wire _2116_;
	wire _2117_;
	wire _2118_;
	wire _2119_;
	wire _2120_;
	wire _2121_;
	wire _2122_;
	wire _2123_;
	wire _2124_;
	wire _2125_;
	wire _2126_;
	wire _2127_;
	wire _2128_;
	wire _2129_;
	wire _2130_;
	wire _2131_;
	wire _2132_;
	wire _2133_;
	wire _2134_;
	wire _2135_;
	wire _2136_;
	wire _2137_;
	wire _2138_;
	wire _2139_;
	wire _2140_;
	wire _2141_;
	wire _2142_;
	wire _2143_;
	wire _2144_;
	wire _2145_;
	wire _2146_;
	wire _2147_;
	wire _2148_;
	wire _2149_;
	wire _2150_;
	wire _2151_;
	wire _2152_;
	wire _2153_;
	wire _2154_;
	wire _2155_;
	wire _2156_;
	wire _2157_;
	wire _2158_;
	wire _2159_;
	wire _2160_;
	wire _2161_;
	wire _2162_;
	wire _2163_;
	wire _2164_;
	wire _2165_;
	wire _2166_;
	wire _2167_;
	wire _2168_;
	wire _2169_;
	wire _2170_;
	wire _2171_;
	wire _2172_;
	wire _2173_;
	wire _2174_;
	wire _2175_;
	wire _2176_;
	wire _2177_;
	wire _2178_;
	wire _2179_;
	wire _2180_;
	wire _2181_;
	wire _2182_;
	wire _2183_;
	wire _2184_;
	wire _2185_;
	wire _2186_;
	wire _2187_;
	wire _2188_;
	wire _2189_;
	wire _2190_;
	wire _2191_;
	wire _2192_;
	wire _2193_;
	wire _2194_;
	wire _2195_;
	wire _2196_;
	wire _2197_;
	wire _2198_;
	wire _2199_;
	wire _2200_;
	wire _2201_;
	wire _2202_;
	wire _2203_;
	wire _2204_;
	wire _2205_;
	wire _2206_;
	wire _2207_;
	wire _2208_;
	wire _2209_;
	wire _2210_;
	wire _2211_;
	wire _2212_;
	wire _2213_;
	wire _2214_;
	wire _2215_;
	wire _2216_;
	wire _2217_;
	wire _2218_;
	wire _2219_;
	wire _2220_;
	wire _2221_;
	wire _2222_;
	wire _2223_;
	wire _2224_;
	wire _2225_;
	wire _2226_;
	wire _2227_;
	wire _2228_;
	wire _2229_;
	wire _2230_;
	wire _2231_;
	wire _2232_;
	wire _2233_;
	wire _2234_;
	wire _2235_;
	wire _2236_;
	wire _2237_;
	wire _2238_;
	wire _2239_;
	wire _2240_;
	wire _2241_;
	wire _2242_;
	wire _2243_;
	wire _2244_;
	wire _2245_;
	wire _2246_;
	wire _2247_;
	wire _2248_;
	wire _2249_;
	wire _2250_;
	wire _2251_;
	wire _2252_;
	wire _2253_;
	wire _2254_;
	wire _2255_;
	wire _2256_;
	wire _2257_;
	wire _2258_;
	wire _2259_;
	wire _2260_;
	wire _2261_;
	wire _2262_;
	wire _2263_;
	wire _2264_;
	wire _2265_;
	wire _2266_;
	wire _2267_;
	wire _2268_;
	wire _2269_;
	wire _2270_;
	wire _2271_;
	wire _2272_;
	wire _2273_;
	wire _2274_;
	wire _2275_;
	wire _2276_;
	wire _2277_;
	wire _2278_;
	wire _2279_;
	wire _2280_;
	wire _2281_;
	wire _2282_;
	wire _2283_;
	wire _2284_;
	wire _2285_;
	wire _2286_;
	wire _2287_;
	wire _2288_;
	wire _2289_;
	wire _2290_;
	wire _2291_;
	wire _2292_;
	wire _2293_;
	wire _2294_;
	wire _2295_;
	wire _2296_;
	wire _2297_;
	wire _2298_;
	wire _2299_;
	wire _2300_;
	wire _2301_;
	wire _2302_;
	wire _2303_;
	wire _2304_;
	wire _2305_;
	wire _2306_;
	wire _2307_;
	wire _2308_;
	wire _2309_;
	wire _2310_;
	wire _2311_;
	wire _2312_;
	wire _2313_;
	wire _2314_;
	wire _2315_;
	wire _2316_;
	wire _2317_;
	wire _2318_;
	wire _2319_;
	wire _2320_;
	wire _2321_;
	wire _2322_;
	wire _2323_;
	wire _2324_;
	wire _2325_;
	wire _2326_;
	wire _2327_;
	wire _2328_;
	wire _2329_;
	wire _2330_;
	wire _2331_;
	wire _2332_;
	wire _2333_;
	wire _2334_;
	wire _2335_;
	wire _2336_;
	wire _2337_;
	wire _2338_;
	wire _2339_;
	wire _2340_;
	wire _2341_;
	wire _2342_;
	wire _2343_;
	wire _2344_;
	wire _2345_;
	wire _2346_;
	wire _2347_;
	wire _2348_;
	wire _2349_;
	wire _2350_;
	wire _2351_;
	wire _2352_;
	wire _2353_;
	wire _2354_;
	wire _2355_;
	wire _2356_;
	wire _2357_;
	wire _2358_;
	wire _2359_;
	wire _2360_;
	wire _2361_;
	wire _2362_;
	wire _2363_;
	wire _2364_;
	wire _2365_;
	wire _2366_;
	wire _2367_;
	wire _2368_;
	wire _2369_;
	wire _2370_;
	wire _2371_;
	wire _2372_;
	wire _2373_;
	wire _2374_;
	wire _2375_;
	wire _2376_;
	wire _2377_;
	wire _2378_;
	wire _2379_;
	wire _2380_;
	wire _2381_;
	wire _2382_;
	wire _2383_;
	wire _2384_;
	wire _2385_;
	wire _2386_;
	wire _2387_;
	wire _2388_;
	wire _2389_;
	wire _2390_;
	wire _2391_;
	wire _2392_;
	wire _2393_;
	wire _2394_;
	wire _2395_;
	wire _2396_;
	wire _2397_;
	wire _2398_;
	wire _2399_;
	wire _2400_;
	wire _2401_;
	wire _2402_;
	wire _2403_;
	wire _2404_;
	wire _2405_;
	wire _2406_;
	wire _2407_;
	wire _2408_;
	wire _2409_;
	wire _2410_;
	wire _2411_;
	wire _2412_;
	wire _2413_;
	wire _2414_;
	wire _2415_;
	wire _2416_;
	wire _2417_;
	wire _2418_;
	wire _2419_;
	wire _2420_;
	wire _2421_;
	wire _2422_;
	wire _2423_;
	wire _2424_;
	wire _2425_;
	wire _2426_;
	wire _2427_;
	wire _2428_;
	wire _2429_;
	wire _2430_;
	wire _2431_;
	wire _2432_;
	wire _2433_;
	wire _2434_;
	wire _2435_;
	wire _2436_;
	wire _2437_;
	wire _2438_;
	wire _2439_;
	wire _2440_;
	wire _2441_;
	wire _2442_;
	wire _2443_;
	wire _2444_;
	wire _2445_;
	wire _2446_;
	wire _2447_;
	wire _2448_;
	wire _2449_;
	wire _2450_;
	wire _2451_;
	wire _2452_;
	wire _2453_;
	wire _2454_;
	wire _2455_;
	wire _2456_;
	wire _2457_;
	wire _2458_;
	wire _2459_;
	wire _2460_;
	wire _2461_;
	wire _2462_;
	wire _2463_;
	wire _2464_;
	wire _2465_;
	wire _2466_;
	wire _2467_;
	wire _2468_;
	wire _2469_;
	wire _2470_;
	wire _2471_;
	wire _2472_;
	wire _2473_;
	wire _2474_;
	wire _2475_;
	wire _2476_;
	wire _2477_;
	wire _2478_;
	wire _2479_;
	wire _2480_;
	wire _2481_;
	wire _2482_;
	wire _2483_;
	wire _2484_;
	wire _2485_;
	wire _2486_;
	wire _2487_;
	wire _2488_;
	wire _2489_;
	wire _2490_;
	wire _2491_;
	wire _2492_;
	wire _2493_;
	wire _2494_;
	wire _2495_;
	wire _2496_;
	wire _2497_;
	wire _2498_;
	wire _2499_;
	wire _2500_;
	wire _2501_;
	wire _2502_;
	wire _2503_;
	wire _2504_;
	wire _2505_;
	wire _2506_;
	wire _2507_;
	wire _2508_;
	wire _2509_;
	wire _2510_;
	wire _2511_;
	wire _2512_;
	wire _2513_;
	wire _2514_;
	wire _2515_;
	wire _2516_;
	wire _2517_;
	wire _2518_;
	wire _2519_;
	wire _2520_;
	wire _2521_;
	wire _2522_;
	wire _2523_;
	wire _2524_;
	wire _2525_;
	wire _2526_;
	wire _2527_;
	wire _2528_;
	wire _2529_;
	wire _2530_;
	wire _2531_;
	wire _2532_;
	wire _2533_;
	wire _2534_;
	wire _2535_;
	wire _2536_;
	wire _2537_;
	wire _2538_;
	wire _2539_;
	wire _2540_;
	wire _2541_;
	wire _2542_;
	wire _2543_;
	wire _2544_;
	wire _2545_;
	wire _2546_;
	wire _2547_;
	wire _2548_;
	wire _2549_;
	wire _2550_;
	wire _2551_;
	wire _2552_;
	wire _2553_;
	wire _2554_;
	wire _2555_;
	wire _2556_;
	wire _2557_;
	wire _2558_;
	wire _2559_;
	wire _2560_;
	wire _2561_;
	wire _2562_;
	wire _2563_;
	wire _2564_;
	wire _2565_;
	wire _2566_;
	wire _2567_;
	wire _2568_;
	wire _2569_;
	wire _2570_;
	wire _2571_;
	wire _2572_;
	wire _2573_;
	wire _2574_;
	wire _2575_;
	wire _2576_;
	wire _2577_;
	wire _2578_;
	wire _2579_;
	wire _2580_;
	wire _2581_;
	wire _2582_;
	wire _2583_;
	wire _2584_;
	wire _2585_;
	wire _2586_;
	wire _2587_;
	wire _2588_;
	wire _2589_;
	wire _2590_;
	wire _2591_;
	wire _2592_;
	wire _2593_;
	wire _2594_;
	wire _2595_;
	wire _2596_;
	wire _2597_;
	wire _2598_;
	wire _2599_;
	wire _2600_;
	wire _2601_;
	wire _2602_;
	wire _2603_;
	wire _2604_;
	wire _2605_;
	wire _2606_;
	wire _2607_;
	wire _2608_;
	wire _2609_;
	wire _2610_;
	wire _2611_;
	wire _2612_;
	wire _2613_;
	wire _2614_;
	wire _2615_;
	wire _2616_;
	wire _2617_;
	wire _2618_;
	wire _2619_;
	wire _2620_;
	wire _2621_;
	wire _2622_;
	wire _2623_;
	wire _2624_;
	wire _2625_;
	wire _2626_;
	wire _2627_;
	wire _2628_;
	wire _2629_;
	wire _2630_;
	wire _2631_;
	wire _2632_;
	wire _2633_;
	wire _2634_;
	wire _2635_;
	wire _2636_;
	wire _2637_;
	wire _2638_;
	wire _2639_;
	wire _2640_;
	wire _2641_;
	wire _2642_;
	wire _2643_;
	wire _2644_;
	wire _2645_;
	wire _2646_;
	wire _2647_;
	wire _2648_;
	wire _2649_;
	wire _2650_;
	wire _2651_;
	wire _2652_;
	wire _2653_;
	wire _2654_;
	wire _2655_;
	wire _2656_;
	wire _2657_;
	wire _2658_;
	wire _2659_;
	wire _2660_;
	wire _2661_;
	wire _2662_;
	wire _2663_;
	wire _2664_;
	wire _2665_;
	wire _2666_;
	wire _2667_;
	wire _2668_;
	wire _2669_;
	wire _2670_;
	wire _2671_;
	wire _2672_;
	wire _2673_;
	wire _2674_;
	wire _2675_;
	wire _2676_;
	wire _2677_;
	wire _2678_;
	wire _2679_;
	wire _2680_;
	wire _2681_;
	wire _2682_;
	wire _2683_;
	wire _2684_;
	wire _2685_;
	wire _2686_;
	wire _2687_;
	wire _2688_;
	wire _2689_;
	wire _2690_;
	wire _2691_;
	wire _2692_;
	wire _2693_;
	wire _2694_;
	wire _2695_;
	wire _2696_;
	wire _2697_;
	wire _2698_;
	wire _2699_;
	wire _2700_;
	wire _2701_;
	wire _2702_;
	wire _2703_;
	wire _2704_;
	wire _2705_;
	wire _2706_;
	wire _2707_;
	wire _2708_;
	wire _2709_;
	wire _2710_;
	wire _2711_;
	wire _2712_;
	wire _2713_;
	wire _2714_;
	wire _2715_;
	wire _2716_;
	wire _2717_;
	wire _2718_;
	wire _2719_;
	wire _2720_;
	wire _2721_;
	wire _2722_;
	wire _2723_;
	wire _2724_;
	wire _2725_;
	wire _2726_;
	wire _2727_;
	wire _2728_;
	wire _2729_;
	wire _2730_;
	wire _2731_;
	wire _2732_;
	wire _2733_;
	wire _2734_;
	wire _2735_;
	wire _2736_;
	wire _2737_;
	wire _2738_;
	wire _2739_;
	wire _2740_;
	wire _2741_;
	wire _2742_;
	wire _2743_;
	wire _2744_;
	wire _2745_;
	wire _2746_;
	wire _2747_;
	wire _2748_;
	wire _2749_;
	wire _2750_;
	wire _2751_;
	wire _2752_;
	wire _2753_;
	wire _2754_;
	wire _2755_;
	wire _2756_;
	wire _2757_;
	wire _2758_;
	wire _2759_;
	wire _2760_;
	wire _2761_;
	wire _2762_;
	wire _2763_;
	wire _2764_;
	wire _2765_;
	wire _2766_;
	wire _2767_;
	wire _2768_;
	wire _2769_;
	wire _2770_;
	wire _2771_;
	wire _2772_;
	wire _2773_;
	wire _2774_;
	wire _2775_;
	wire _2776_;
	wire _2777_;
	wire _2778_;
	wire _2779_;
	wire _2780_;
	wire _2781_;
	wire _2782_;
	wire _2783_;
	wire _2784_;
	wire _2785_;
	wire _2786_;
	wire _2787_;
	wire _2788_;
	wire _2789_;
	wire _2790_;
	wire _2791_;
	wire _2792_;
	wire _2793_;
	wire _2794_;
	wire _2795_;
	wire _2796_;
	wire _2797_;
	wire _2798_;
	wire _2799_;
	wire _2800_;
	wire _2801_;
	wire _2802_;
	wire _2803_;
	wire _2804_;
	wire _2805_;
	wire _2806_;
	wire _2807_;
	wire _2808_;
	wire _2809_;
	wire _2810_;
	wire _2811_;
	wire _2812_;
	wire _2813_;
	wire _2814_;
	wire _2815_;
	wire _2816_;
	wire _2817_;
	wire _2818_;
	wire _2819_;
	wire _2820_;
	wire _2821_;
	wire _2822_;
	wire _2823_;
	wire _2824_;
	wire _2825_;
	wire _2826_;
	wire _2827_;
	wire _2828_;
	wire _2829_;
	wire _2830_;
	wire _2831_;
	wire _2832_;
	wire _2833_;
	wire _2834_;
	wire _2835_;
	wire _2836_;
	wire _2837_;
	wire _2838_;
	wire _2839_;
	wire _2840_;
	wire _2841_;
	wire _2842_;
	wire _2843_;
	wire _2844_;
	wire _2845_;
	wire _2846_;
	wire _2847_;
	wire _2848_;
	wire _2849_;
	wire _2850_;
	wire _2851_;
	wire _2852_;
	wire _2853_;
	wire _2854_;
	wire _2855_;
	wire _2856_;
	wire _2857_;
	wire _2858_;
	wire _2859_;
	wire _2860_;
	wire _2861_;
	wire _2862_;
	wire _2863_;
	wire _2864_;
	wire _2865_;
	wire _2866_;
	wire _2867_;
	wire _2868_;
	wire _2869_;
	wire _2870_;
	wire _2871_;
	wire _2872_;
	wire _2873_;
	wire _2874_;
	wire _2875_;
	wire _2876_;
	wire _2877_;
	wire _2878_;
	wire _2879_;
	wire _2880_;
	wire _2881_;
	wire _2882_;
	wire _2883_;
	wire _2884_;
	wire _2885_;
	wire _2886_;
	wire _2887_;
	wire _2888_;
	wire _2889_;
	wire _2890_;
	wire _2891_;
	wire _2892_;
	wire _2893_;
	wire _2894_;
	wire _2895_;
	wire _2896_;
	wire _2897_;
	wire _2898_;
	wire _2899_;
	wire _2900_;
	wire _2901_;
	wire _2902_;
	wire _2903_;
	wire _2904_;
	wire _2905_;
	wire _2906_;
	wire _2907_;
	wire _2908_;
	wire _2909_;
	wire _2910_;
	wire _2911_;
	wire _2912_;
	wire _2913_;
	wire _2914_;
	wire _2915_;
	wire _2916_;
	wire _2917_;
	wire _2918_;
	wire _2919_;
	wire _2920_;
	wire _2921_;
	wire _2922_;
	wire _2923_;
	wire _2924_;
	wire _2925_;
	wire _2926_;
	wire _2927_;
	wire _2928_;
	wire _2929_;
	wire _2930_;
	wire _2931_;
	wire _2932_;
	wire _2933_;
	wire _2934_;
	wire _2935_;
	wire _2936_;
	wire _2937_;
	wire _2938_;
	wire _2939_;
	wire _2940_;
	wire _2941_;
	wire _2942_;
	wire _2943_;
	wire _2944_;
	wire _2945_;
	wire _2946_;
	wire _2947_;
	wire _2948_;
	wire _2949_;
	wire _2950_;
	wire _2951_;
	wire _2952_;
	wire _2953_;
	wire _2954_;
	wire _2955_;
	wire _2956_;
	wire _2957_;
	wire _2958_;
	wire _2959_;
	wire _2960_;
	wire _2961_;
	wire _2962_;
	wire _2963_;
	wire _2964_;
	wire _2965_;
	wire _2966_;
	wire _2967_;
	wire _2968_;
	wire _2969_;
	wire _2970_;
	wire _2971_;
	wire _2972_;
	wire _2973_;
	wire _2974_;
	wire _2975_;
	wire _2976_;
	wire _2977_;
	wire _2978_;
	wire _2979_;
	wire _2980_;
	wire _2981_;
	wire _2982_;
	wire _2983_;
	wire _2984_;
	wire _2985_;
	wire _2986_;
	wire _2987_;
	wire _2988_;
	wire _2989_;
	wire _2990_;
	wire _2991_;
	wire _2992_;
	wire _2993_;
	wire _2994_;
	wire _2995_;
	wire _2996_;
	wire _2997_;
	wire _2998_;
	wire _2999_;
	wire _3000_;
	wire _3001_;
	wire _3002_;
	wire _3003_;
	wire _3004_;
	wire _3005_;
	wire _3006_;
	wire _3007_;
	wire _3008_;
	wire _3009_;
	wire _3010_;
	wire _3011_;
	wire _3012_;
	wire _3013_;
	wire _3014_;
	wire _3015_;
	wire _3016_;
	wire _3017_;
	wire _3018_;
	wire _3019_;
	wire _3020_;
	wire _3021_;
	wire _3022_;
	wire _3023_;
	wire _3024_;
	wire _3025_;
	wire _3026_;
	wire _3027_;
	wire _3028_;
	wire _3029_;
	wire _3030_;
	wire _3031_;
	wire _3032_;
	wire _3033_;
	wire _3034_;
	wire _3035_;
	wire _3036_;
	wire _3037_;
	wire _3038_;
	wire _3039_;
	wire _3040_;
	wire _3041_;
	wire _3042_;
	wire _3043_;
	wire _3044_;
	wire _3045_;
	wire _3046_;
	wire _3047_;
	wire _3048_;
	wire _3049_;
	wire _3050_;
	wire _3051_;
	wire _3052_;
	wire _3053_;
	wire _3054_;
	wire _3055_;
	wire _3056_;
	wire _3057_;
	wire _3058_;
	wire _3059_;
	wire _3060_;
	wire _3061_;
	wire _3062_;
	wire _3063_;
	wire _3064_;
	wire _3065_;
	wire _3066_;
	wire _3067_;
	wire _3068_;
	wire _3069_;
	wire _3070_;
	wire _3071_;
	wire _3072_;
	wire _3073_;
	wire _3074_;
	wire _3075_;
	wire _3076_;
	wire _3077_;
	wire _3078_;
	wire _3079_;
	wire _3080_;
	wire _3081_;
	wire _3082_;
	wire _3083_;
	wire _3084_;
	wire _3085_;
	wire _3086_;
	wire _3087_;
	wire _3088_;
	wire _3089_;
	wire _3090_;
	wire _3091_;
	wire _3092_;
	wire _3093_;
	wire _3094_;
	wire _3095_;
	wire _3096_;
	wire _3097_;
	wire _3098_;
	wire _3099_;
	wire _3100_;
	wire _3101_;
	wire _3102_;
	wire _3103_;
	wire _3104_;
	wire _3105_;
	wire _3106_;
	wire _3107_;
	wire _3108_;
	wire _3109_;
	wire _3110_;
	wire _3111_;
	wire _3112_;
	wire _3113_;
	wire _3114_;
	wire _3115_;
	wire _3116_;
	wire _3117_;
	wire _3118_;
	wire _3119_;
	wire _3120_;
	wire _3121_;
	wire _3122_;
	wire _3123_;
	wire _3124_;
	wire _3125_;
	wire _3126_;
	wire _3127_;
	wire _3128_;
	wire _3129_;
	wire _3130_;
	wire _3131_;
	wire _3132_;
	wire _3133_;
	wire _3134_;
	wire _3135_;
	wire _3136_;
	wire _3137_;
	wire _3138_;
	wire _3139_;
	wire _3140_;
	wire _3141_;
	wire _3142_;
	wire _3143_;
	wire _3144_;
	wire _3145_;
	wire _3146_;
	wire _3147_;
	wire _3148_;
	wire _3149_;
	wire _3150_;
	wire _3151_;
	wire _3152_;
	wire _3153_;
	wire _3154_;
	wire _3155_;
	wire _3156_;
	wire _3157_;
	wire _3158_;
	wire _3159_;
	wire _3160_;
	wire _3161_;
	wire _3162_;
	wire _3163_;
	wire _3164_;
	wire _3165_;
	wire _3166_;
	wire _3167_;
	wire _3168_;
	wire _3169_;
	wire _3170_;
	wire _3171_;
	wire _3172_;
	wire _3173_;
	wire _3174_;
	wire _3175_;
	wire _3176_;
	wire _3177_;
	wire _3178_;
	wire _3179_;
	wire _3180_;
	wire _3181_;
	wire _3182_;
	wire _3183_;
	wire _3184_;
	wire _3185_;
	wire _3186_;
	wire _3187_;
	wire _3188_;
	wire _3189_;
	wire _3190_;
	wire _3191_;
	wire _3192_;
	wire _3193_;
	wire _3194_;
	wire _3195_;
	wire _3196_;
	wire _3197_;
	wire _3198_;
	wire _3199_;
	wire _3200_;
	wire _3201_;
	wire _3202_;
	wire _3203_;
	wire _3204_;
	wire _3205_;
	wire _3206_;
	wire _3207_;
	wire _3208_;
	wire _3209_;
	wire _3210_;
	wire _3211_;
	wire _3212_;
	wire _3213_;
	wire _3214_;
	wire _3215_;
	wire _3216_;
	wire _3217_;
	wire _3218_;
	wire _3219_;
	wire _3220_;
	wire _3221_;
	wire _3222_;
	wire _3223_;
	wire _3224_;
	wire _3225_;
	wire _3226_;
	wire _3227_;
	wire _3228_;
	wire _3229_;
	wire _3230_;
	wire _3231_;
	wire _3232_;
	wire _3233_;
	wire _3234_;
	wire _3235_;
	wire _3236_;
	wire _3237_;
	wire _3238_;
	wire _3239_;
	wire _3240_;
	wire _3241_;
	wire _3242_;
	wire _3243_;
	wire _3244_;
	wire _3245_;
	wire _3246_;
	wire _3247_;
	wire _3248_;
	wire _3249_;
	wire _3250_;
	wire _3251_;
	wire _3252_;
	wire _3253_;
	wire _3254_;
	wire _3255_;
	wire _3256_;
	wire _3257_;
	wire _3258_;
	wire _3259_;
	wire _3260_;
	wire _3261_;
	wire _3262_;
	wire _3263_;
	wire _3264_;
	wire _3265_;
	wire _3266_;
	wire _3267_;
	wire _3268_;
	wire _3269_;
	wire _3270_;
	wire _3271_;
	wire _3272_;
	wire _3273_;
	wire _3274_;
	wire _3275_;
	wire _3276_;
	wire _3277_;
	wire _3278_;
	wire _3279_;
	wire _3280_;
	wire _3281_;
	wire _3282_;
	wire _3283_;
	wire _3284_;
	wire _3285_;
	wire _3286_;
	wire _3287_;
	wire _3288_;
	wire _3289_;
	wire _3290_;
	wire _3291_;
	wire _3292_;
	wire _3293_;
	wire _3294_;
	wire _3295_;
	wire _3296_;
	wire _3297_;
	wire _3298_;
	wire _3299_;
	wire _3300_;
	wire _3301_;
	wire _3302_;
	wire _3303_;
	wire _3304_;
	wire _3305_;
	wire _3306_;
	wire _3307_;
	wire _3308_;
	wire _3309_;
	wire _3310_;
	wire _3311_;
	wire _3312_;
	wire _3313_;
	wire _3314_;
	wire _3315_;
	wire _3316_;
	wire _3317_;
	wire _3318_;
	wire _3319_;
	wire _3320_;
	wire _3321_;
	wire _3322_;
	wire _3323_;
	wire _3324_;
	wire _3325_;
	wire _3326_;
	wire _3327_;
	wire _3328_;
	wire _3329_;
	wire _3330_;
	wire _3331_;
	wire _3332_;
	wire _3333_;
	wire _3334_;
	wire _3335_;
	wire _3336_;
	wire _3337_;
	wire _3338_;
	wire _3339_;
	wire _3340_;
	wire _3341_;
	wire _3342_;
	wire _3343_;
	wire _3344_;
	wire _3345_;
	wire _3346_;
	wire _3347_;
	wire _3348_;
	wire _3349_;
	wire _3350_;
	wire _3351_;
	wire _3352_;
	wire _3353_;
	wire _3354_;
	wire _3355_;
	wire _3356_;
	wire _3357_;
	wire _3358_;
	wire _3359_;
	wire _3360_;
	wire _3361_;
	wire _3362_;
	wire _3363_;
	wire _3364_;
	wire _3365_;
	wire _3366_;
	wire _3367_;
	wire _3368_;
	wire _3369_;
	wire _3370_;
	wire _3371_;
	wire _3372_;
	wire _3373_;
	wire _3374_;
	wire _3375_;
	wire _3376_;
	wire _3377_;
	wire _3378_;
	wire _3379_;
	wire _3380_;
	wire _3381_;
	wire _3382_;
	wire _3383_;
	wire _3384_;
	wire _3385_;
	wire _3386_;
	wire _3387_;
	wire _3388_;
	wire _3389_;
	wire _3390_;
	wire _3391_;
	wire _3392_;
	wire _3393_;
	wire _3394_;
	wire _3395_;
	wire _3396_;
	wire _3397_;
	wire _3398_;
	wire _3399_;
	wire _3400_;
	wire _3401_;
	wire _3402_;
	wire _3403_;
	wire _3404_;
	wire _3405_;
	wire _3406_;
	wire _3407_;
	wire _3408_;
	wire _3409_;
	wire _3410_;
	wire _3411_;
	wire _3412_;
	wire _3413_;
	wire _3414_;
	wire _3415_;
	wire _3416_;
	wire _3417_;
	wire _3418_;
	wire _3419_;
	wire _3420_;
	wire _3421_;
	wire _3422_;
	wire _3423_;
	wire _3424_;
	wire _3425_;
	wire _3426_;
	wire _3427_;
	wire _3428_;
	wire _3429_;
	wire _3430_;
	wire _3431_;
	wire _3432_;
	wire _3433_;
	wire _3434_;
	wire _3435_;
	wire _3436_;
	wire _3437_;
	wire _3438_;
	wire _3439_;
	wire _3440_;
	wire _3441_;
	wire _3442_;
	wire _3443_;
	wire _3444_;
	wire _3445_;
	wire _3446_;
	wire _3447_;
	wire _3448_;
	wire _3449_;
	wire _3450_;
	wire _3451_;
	wire _3452_;
	wire _3453_;
	wire _3454_;
	wire _3455_;
	wire _3456_;
	wire _3457_;
	wire _3458_;
	wire _3459_;
	wire _3460_;
	wire _3461_;
	wire _3462_;
	wire _3463_;
	wire _3464_;
	wire _3465_;
	wire _3466_;
	wire _3467_;
	wire _3468_;
	wire _3469_;
	wire _3470_;
	wire _3471_;
	wire _3472_;
	wire _3473_;
	wire _3474_;
	wire _3475_;
	wire _3476_;
	wire _3477_;
	wire _3478_;
	wire _3479_;
	wire _3480_;
	wire _3481_;
	wire _3482_;
	wire _3483_;
	wire _3484_;
	wire _3485_;
	wire _3486_;
	wire _3487_;
	wire _3488_;
	wire _3489_;
	wire _3490_;
	wire _3491_;
	wire _3492_;
	wire _3493_;
	wire _3494_;
	wire _3495_;
	wire _3496_;
	wire _3497_;
	wire _3498_;
	wire _3499_;
	wire _3500_;
	wire _3501_;
	wire _3502_;
	wire _3503_;
	wire _3504_;
	wire _3505_;
	wire _3506_;
	wire _3507_;
	wire _3508_;
	wire _3509_;
	wire _3510_;
	wire _3511_;
	wire _3512_;
	wire _3513_;
	wire _3514_;
	wire _3515_;
	wire _3516_;
	wire _3517_;
	wire _3518_;
	wire _3519_;
	wire _3520_;
	wire _3521_;
	wire _3522_;
	wire _3523_;
	wire _3524_;
	wire _3525_;
	wire _3526_;
	wire _3527_;
	wire _3528_;
	wire _3529_;
	wire _3530_;
	wire _3531_;
	wire _3532_;
	wire _3533_;
	wire _3534_;
	wire _3535_;
	wire _3536_;
	wire _3537_;
	wire _3538_;
	wire _3539_;
	wire _3540_;
	wire _3541_;
	wire _3542_;
	wire _3543_;
	wire _3544_;
	wire _3545_;
	wire _3546_;
	wire _3547_;
	wire _3548_;
	wire _3549_;
	wire _3550_;
	wire _3551_;
	wire _3552_;
	wire _3553_;
	wire _3554_;
	wire _3555_;
	wire _3556_;
	wire _3557_;
	wire _3558_;
	wire _3559_;
	wire _3560_;
	wire _3561_;
	wire _3562_;
	wire _3563_;
	wire _3564_;
	wire _3565_;
	wire _3566_;
	wire _3567_;
	wire _3568_;
	wire _3569_;
	wire _3570_;
	wire _3571_;
	wire _3572_;
	wire _3573_;
	wire _3574_;
	wire _3575_;
	wire _3576_;
	wire _3577_;
	wire _3578_;
	wire _3579_;
	wire _3580_;
	wire _3581_;
	wire _3582_;
	wire _3583_;
	wire _3584_;
	wire _3585_;
	wire _3586_;
	wire _3587_;
	wire _3588_;
	wire _3589_;
	wire _3590_;
	wire _3591_;
	wire _3592_;
	wire _3593_;
	wire _3594_;
	wire _3595_;
	wire _3596_;
	wire _3597_;
	wire _3598_;
	wire _3599_;
	wire _3600_;
	wire _3601_;
	wire _3602_;
	wire _3603_;
	wire _3604_;
	wire _3605_;
	wire _3606_;
	wire _3607_;
	wire _3608_;
	wire _3609_;
	wire _3610_;
	wire _3611_;
	wire _3612_;
	wire _3613_;
	wire _3614_;
	wire _3615_;
	wire _3616_;
	wire _3617_;
	wire _3618_;
	wire _3619_;
	wire _3620_;
	wire _3621_;
	wire _3622_;
	wire _3623_;
	wire _3624_;
	wire _3625_;
	wire _3626_;
	wire _3627_;
	wire _3628_;
	wire _3629_;
	wire _3630_;
	wire _3631_;
	wire _3632_;
	wire _3633_;
	wire _3634_;
	wire _3635_;
	wire _3636_;
	wire _3637_;
	wire _3638_;
	wire _3639_;
	wire _3640_;
	wire _3641_;
	wire _3642_;
	wire _3643_;
	wire _3644_;
	wire _3645_;
	wire _3646_;
	wire _3647_;
	wire _3648_;
	wire _3649_;
	wire _3650_;
	wire _3651_;
	wire _3652_;
	wire _3653_;
	wire _3654_;
	wire _3655_;
	wire _3656_;
	wire _3657_;
	wire _3658_;
	wire _3659_;
	wire _3660_;
	wire _3661_;
	wire _3662_;
	wire _3663_;
	wire _3664_;
	wire _3665_;
	wire _3666_;
	wire _3667_;
	wire _3668_;
	wire _3669_;
	wire _3670_;
	wire _3671_;
	wire _3672_;
	wire _3673_;
	wire _3674_;
	wire _3675_;
	wire _3676_;
	wire _3677_;
	wire _3678_;
	wire _3679_;
	wire _3680_;
	wire _3681_;
	wire _3682_;
	wire _3683_;
	wire _3684_;
	wire _3685_;
	wire _3686_;
	wire _3687_;
	wire _3688_;
	wire _3689_;
	wire _3690_;
	wire _3691_;
	wire _3692_;
	wire _3693_;
	wire _3694_;
	wire _3695_;
	wire _3696_;
	wire _3697_;
	wire _3698_;
	wire _3699_;
	wire _3700_;
	wire _3701_;
	wire _3702_;
	wire _3703_;
	wire _3704_;
	wire _3705_;
	wire _3706_;
	wire _3707_;
	wire _3708_;
	wire _3709_;
	wire _3710_;
	wire _3711_;
	wire _3712_;
	wire _3713_;
	wire _3714_;
	wire _3715_;
	wire _3716_;
	wire _3717_;
	wire _3718_;
	wire _3719_;
	wire _3720_;
	wire _3721_;
	wire _3722_;
	wire _3723_;
	wire _3724_;
	wire _3725_;
	wire _3726_;
	wire _3727_;
	wire _3728_;
	wire _3729_;
	wire _3730_;
	wire _3731_;
	wire _3732_;
	wire _3733_;
	wire _3734_;
	wire _3735_;
	wire _3736_;
	wire _3737_;
	wire _3738_;
	wire _3739_;
	wire _3740_;
	wire _3741_;
	wire _3742_;
	wire _3743_;
	wire _3744_;
	wire _3745_;
	wire _3746_;
	wire _3747_;
	wire _3748_;
	wire _3749_;
	wire _3750_;
	wire _3751_;
	wire _3752_;
	wire _3753_;
	wire _3754_;
	wire _3755_;
	wire _3756_;
	wire _3757_;
	wire _3758_;
	wire _3759_;
	wire _3760_;
	wire _3761_;
	wire _3762_;
	wire _3763_;
	wire _3764_;
	wire _3765_;
	wire _3766_;
	wire _3767_;
	wire _3768_;
	wire _3769_;
	wire _3770_;
	wire _3771_;
	wire _3772_;
	wire _3773_;
	wire _3774_;
	wire _3775_;
	wire _3776_;
	wire _3777_;
	wire _3778_;
	wire _3779_;
	wire _3780_;
	wire _3781_;
	wire _3782_;
	wire _3783_;
	wire _3784_;
	wire _3785_;
	wire _3786_;
	wire _3787_;
	wire _3788_;
	wire _3789_;
	wire _3790_;
	wire _3791_;
	wire _3792_;
	wire _3793_;
	wire _3794_;
	wire _3795_;
	wire _3796_;
	wire _3797_;
	wire _3798_;
	wire _3799_;
	wire _3800_;
	wire _3801_;
	wire _3802_;
	wire _3803_;
	wire _3804_;
	wire _3805_;
	wire _3806_;
	wire _3807_;
	wire _3808_;
	wire _3809_;
	wire _3810_;
	wire _3811_;
	wire _3812_;
	wire _3813_;
	wire _3814_;
	wire _3815_;
	wire _3816_;
	wire _3817_;
	wire _3818_;
	wire _3819_;
	wire _3820_;
	wire _3821_;
	wire _3822_;
	wire _3823_;
	wire _3824_;
	wire _3825_;
	wire _3826_;
	wire _3827_;
	wire _3828_;
	wire _3829_;
	wire _3830_;
	wire _3831_;
	wire _3832_;
	wire _3833_;
	wire _3834_;
	wire _3835_;
	wire _3836_;
	wire _3837_;
	wire _3838_;
	wire _3839_;
	wire _3840_;
	wire _3841_;
	wire _3842_;
	wire _3843_;
	wire _3844_;
	wire _3845_;
	wire _3846_;
	wire _3847_;
	wire _3848_;
	wire _3849_;
	wire _3850_;
	wire _3851_;
	wire _3852_;
	wire _3853_;
	wire _3854_;
	wire _3855_;
	wire _3856_;
	wire _3857_;
	wire _3858_;
	wire _3859_;
	wire _3860_;
	wire _3861_;
	wire _3862_;
	wire _3863_;
	wire _3864_;
	wire _3865_;
	wire _3866_;
	wire _3867_;
	wire _3868_;
	wire _3869_;
	wire _3870_;
	wire _3871_;
	wire _3872_;
	wire _3873_;
	wire _3874_;
	wire _3875_;
	wire _3876_;
	wire _3877_;
	wire _3878_;
	wire _3879_;
	wire _3880_;
	wire _3881_;
	wire _3882_;
	wire _3883_;
	wire _3884_;
	wire _3885_;
	wire _3886_;
	wire _3887_;
	wire _3888_;
	wire _3889_;
	wire _3890_;
	wire _3891_;
	wire _3892_;
	wire _3893_;
	wire _3894_;
	wire _3895_;
	wire _3896_;
	wire _3897_;
	wire _3898_;
	wire _3899_;
	wire _3900_;
	wire _3901_;
	wire _3902_;
	wire _3903_;
	wire _3904_;
	wire _3905_;
	wire _3906_;
	wire _3907_;
	wire _3908_;
	wire _3909_;
	wire _3910_;
	wire _3911_;
	wire _3912_;
	wire _3913_;
	wire _3914_;
	wire _3915_;
	wire _3916_;
	wire _3917_;
	wire _3918_;
	wire _3919_;
	wire _3920_;
	wire _3921_;
	wire _3922_;
	wire _3923_;
	wire _3924_;
	wire _3925_;
	wire _3926_;
	wire _3927_;
	wire _3928_;
	wire _3929_;
	wire _3930_;
	wire _3931_;
	wire _3932_;
	wire _3933_;
	wire _3934_;
	wire _3935_;
	wire _3936_;
	wire _3937_;
	wire _3938_;
	wire _3939_;
	wire _3940_;
	wire _3941_;
	wire _3942_;
	wire _3943_;
	wire _3944_;
	wire _3945_;
	wire _3946_;
	wire _3947_;
	wire _3948_;
	wire _3949_;
	wire _3950_;
	wire _3951_;
	wire _3952_;
	wire _3953_;
	wire _3954_;
	wire _3955_;
	wire _3956_;
	wire _3957_;
	wire _3958_;
	wire _3959_;
	wire _3960_;
	wire _3961_;
	wire _3962_;
	wire _3963_;
	wire _3964_;
	wire _3965_;
	wire _3966_;
	wire _3967_;
	wire _3968_;
	wire _3969_;
	wire _3970_;
	wire _3971_;
	wire _3972_;
	wire _3973_;
	wire _3974_;
	wire _3975_;
	wire _3976_;
	wire _3977_;
	wire _3978_;
	wire _3979_;
	wire _3980_;
	wire _3981_;
	wire _3982_;
	wire _3983_;
	wire _3984_;
	wire _3985_;
	wire _3986_;
	wire _3987_;
	wire _3988_;
	wire _3989_;
	wire _3990_;
	wire _3991_;
	wire _3992_;
	wire _3993_;
	wire _3994_;
	wire _3995_;
	wire _3996_;
	wire _3997_;
	wire _3998_;
	wire _3999_;
	wire _4000_;
	wire _4001_;
	wire _4002_;
	wire _4003_;
	wire _4004_;
	wire _4005_;
	wire _4006_;
	wire _4007_;
	wire _4008_;
	wire _4009_;
	wire _4010_;
	wire _4011_;
	wire _4012_;
	wire _4013_;
	wire _4014_;
	wire _4015_;
	wire _4016_;
	wire _4017_;
	wire _4018_;
	wire _4019_;
	wire _4020_;
	wire _4021_;
	wire _4022_;
	wire _4023_;
	wire _4024_;
	wire _4025_;
	wire _4026_;
	wire _4027_;
	wire _4028_;
	wire _4029_;
	wire _4030_;
	wire _4031_;
	wire _4032_;
	wire _4033_;
	wire _4034_;
	wire _4035_;
	wire _4036_;
	wire _4037_;
	wire _4038_;
	wire _4039_;
	wire _4040_;
	wire _4041_;
	wire _4042_;
	wire _4043_;
	wire _4044_;
	wire _4045_;
	wire _4046_;
	wire _4047_;
	wire _4048_;
	wire _4049_;
	wire _4050_;
	wire _4051_;
	wire _4052_;
	wire _4053_;
	wire _4054_;
	wire _4055_;
	wire _4056_;
	wire _4057_;
	wire _4058_;
	wire _4059_;
	wire _4060_;
	wire _4061_;
	wire _4062_;
	wire _4063_;
	wire _4064_;
	wire _4065_;
	wire _4066_;
	wire _4067_;
	wire _4068_;
	wire _4069_;
	wire _4070_;
	wire _4071_;
	wire _4072_;
	wire _4073_;
	wire _4074_;
	wire _4075_;
	wire _4076_;
	wire _4077_;
	wire _4078_;
	wire _4079_;
	wire _4080_;
	wire _4081_;
	wire _4082_;
	wire _4083_;
	wire _4084_;
	wire _4085_;
	wire _4086_;
	wire _4087_;
	wire _4088_;
	wire _4089_;
	wire _4090_;
	wire _4091_;
	wire _4092_;
	wire _4093_;
	wire _4094_;
	wire _4095_;
	wire _4096_;
	wire _4097_;
	wire _4098_;
	wire _4099_;
	wire _4100_;
	wire _4101_;
	wire _4102_;
	wire _4103_;
	wire _4104_;
	wire _4105_;
	wire _4106_;
	wire _4107_;
	wire _4108_;
	wire _4109_;
	wire _4110_;
	wire _4111_;
	wire _4112_;
	wire _4113_;
	wire _4114_;
	wire _4115_;
	wire _4116_;
	wire _4117_;
	wire _4118_;
	wire _4119_;
	wire _4120_;
	wire _4121_;
	wire _4122_;
	wire _4123_;
	wire _4124_;
	wire _4125_;
	wire _4126_;
	wire _4127_;
	wire _4128_;
	wire _4129_;
	wire _4130_;
	wire _4131_;
	wire _4132_;
	wire _4133_;
	wire _4134_;
	wire _4135_;
	wire _4136_;
	wire _4137_;
	wire _4138_;
	wire _4139_;
	wire _4140_;
	wire _4141_;
	wire _4142_;
	wire _4143_;
	wire _4144_;
	wire _4145_;
	wire _4146_;
	wire _4147_;
	wire _4148_;
	wire _4149_;
	wire _4150_;
	wire _4151_;
	wire _4152_;
	wire _4153_;
	wire _4154_;
	wire _4155_;
	wire _4156_;
	wire _4157_;
	wire _4158_;
	wire _4159_;
	wire _4160_;
	wire _4161_;
	wire _4162_;
	wire _4163_;
	wire _4164_;
	wire _4165_;
	wire _4166_;
	wire _4167_;
	wire _4168_;
	wire _4169_;
	wire _4170_;
	wire _4171_;
	wire _4172_;
	wire _4173_;
	wire _4174_;
	wire _4175_;
	wire _4176_;
	wire _4177_;
	wire _4178_;
	wire _4179_;
	wire _4180_;
	wire _4181_;
	wire _4182_;
	wire _4183_;
	wire _4184_;
	wire _4185_;
	wire _4186_;
	wire _4187_;
	wire _4188_;
	wire _4189_;
	wire _4190_;
	wire _4191_;
	wire _4192_;
	wire _4193_;
	wire _4194_;
	wire _4195_;
	wire _4196_;
	wire _4197_;
	wire _4198_;
	wire _4199_;
	wire _4200_;
	wire _4201_;
	wire _4202_;
	wire _4203_;
	wire _4204_;
	wire _4205_;
	wire _4206_;
	wire _4207_;
	wire _4208_;
	wire _4209_;
	wire _4210_;
	wire _4211_;
	wire _4212_;
	wire _4213_;
	wire _4214_;
	wire _4215_;
	wire _4216_;
	wire _4217_;
	wire _4218_;
	wire _4219_;
	wire _4220_;
	wire _4221_;
	wire _4222_;
	wire _4223_;
	wire _4224_;
	wire _4225_;
	wire _4226_;
	wire _4227_;
	wire _4228_;
	wire _4229_;
	wire _4230_;
	wire _4231_;
	wire _4232_;
	wire _4233_;
	wire _4234_;
	wire _4235_;
	wire _4236_;
	wire _4237_;
	wire _4238_;
	wire _4239_;
	wire _4240_;
	wire _4241_;
	wire _4242_;
	wire _4243_;
	wire _4244_;
	wire _4245_;
	wire _4246_;
	wire _4247_;
	wire _4248_;
	wire _4249_;
	wire _4250_;
	wire _4251_;
	wire _4252_;
	wire _4253_;
	wire _4254_;
	wire _4255_;
	wire _4256_;
	wire _4257_;
	wire _4258_;
	wire _4259_;
	wire _4260_;
	wire _4261_;
	wire _4262_;
	wire _4263_;
	wire _4264_;
	wire _4265_;
	wire _4266_;
	wire _4267_;
	wire _4268_;
	wire _4269_;
	wire _4270_;
	wire _4271_;
	wire _4272_;
	wire _4273_;
	wire _4274_;
	wire _4275_;
	wire _4276_;
	wire _4277_;
	wire _4278_;
	wire _4279_;
	wire _4280_;
	wire _4281_;
	wire _4282_;
	wire _4283_;
	wire _4284_;
	wire _4285_;
	wire _4286_;
	wire _4287_;
	wire _4288_;
	wire _4289_;
	wire _4290_;
	wire _4291_;
	wire _4292_;
	wire _4293_;
	wire _4294_;
	wire _4295_;
	wire _4296_;
	wire _4297_;
	wire _4298_;
	wire _4299_;
	wire _4300_;
	wire _4301_;
	wire _4302_;
	wire _4303_;
	wire _4304_;
	wire _4305_;
	wire _4306_;
	wire _4307_;
	wire _4308_;
	wire _4309_;
	wire _4310_;
	wire _4311_;
	wire _4312_;
	wire _4313_;
	wire _4314_;
	wire _4315_;
	wire _4316_;
	wire _4317_;
	wire _4318_;
	wire _4319_;
	wire _4320_;
	wire _4321_;
	wire _4322_;
	wire _4323_;
	wire _4324_;
	wire _4325_;
	wire _4326_;
	wire _4327_;
	wire _4328_;
	wire _4329_;
	wire _4330_;
	wire _4331_;
	wire _4332_;
	wire _4333_;
	wire _4334_;
	wire _4335_;
	wire _4336_;
	wire _4337_;
	wire _4338_;
	wire _4339_;
	wire _4340_;
	wire _4341_;
	wire _4342_;
	wire _4343_;
	wire _4344_;
	wire _4345_;
	wire _4346_;
	wire _4347_;
	wire _4348_;
	wire _4349_;
	wire _4350_;
	wire _4351_;
	wire _4352_;
	wire _4353_;
	wire _4354_;
	wire _4355_;
	wire _4356_;
	wire _4357_;
	wire _4358_;
	wire _4359_;
	wire _4360_;
	wire _4361_;
	wire _4362_;
	wire _4363_;
	wire _4364_;
	wire _4365_;
	wire _4366_;
	wire _4367_;
	wire _4368_;
	wire _4369_;
	wire _4370_;
	wire _4371_;
	wire _4372_;
	wire _4373_;
	wire _4374_;
	wire _4375_;
	wire _4376_;
	wire _4377_;
	wire _4378_;
	wire _4379_;
	wire _4380_;
	wire _4381_;
	wire _4382_;
	wire _4383_;
	wire _4384_;
	wire _4385_;
	wire _4386_;
	wire _4387_;
	wire _4388_;
	wire _4389_;
	wire _4390_;
	wire _4391_;
	wire _4392_;
	wire _4393_;
	wire _4394_;
	wire _4395_;
	wire _4396_;
	wire _4397_;
	wire _4398_;
	wire _4399_;
	wire _4400_;
	wire _4401_;
	wire _4402_;
	wire _4403_;
	wire _4404_;
	wire _4405_;
	wire _4406_;
	wire _4407_;
	wire _4408_;
	wire _4409_;
	wire _4410_;
	wire _4411_;
	wire _4412_;
	wire _4413_;
	wire _4414_;
	wire _4415_;
	wire _4416_;
	wire _4417_;
	wire _4418_;
	wire _4419_;
	wire _4420_;
	wire _4421_;
	wire _4422_;
	wire _4423_;
	wire _4424_;
	wire _4425_;
	wire _4426_;
	wire _4427_;
	wire _4428_;
	wire _4429_;
	wire _4430_;
	wire _4431_;
	wire _4432_;
	wire _4433_;
	wire _4434_;
	wire _4435_;
	wire _4436_;
	wire _4437_;
	wire _4438_;
	wire _4439_;
	wire _4440_;
	wire _4441_;
	wire _4442_;
	wire _4443_;
	wire _4444_;
	wire _4445_;
	wire _4446_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire [7:0] \mchip.pong.VGA_B ;
	wire \mchip.pong.VGA_B0 ;
	wire \mchip.pong.VGA_B1 ;
	wire \mchip.pong.VGA_B2 ;
	wire \mchip.pong.VGA_B3 ;
	wire [7:0] \mchip.pong.VGA_G ;
	wire \mchip.pong.VGA_G0 ;
	wire \mchip.pong.VGA_G1 ;
	wire \mchip.pong.VGA_G2 ;
	wire \mchip.pong.VGA_G3 ;
	wire \mchip.pong.VGA_HS ;
	wire [7:0] \mchip.pong.VGA_R ;
	wire \mchip.pong.VGA_R0 ;
	wire \mchip.pong.VGA_R1 ;
	wire \mchip.pong.VGA_R2 ;
	wire \mchip.pong.VGA_R3 ;
	wire \mchip.pong.VGA_VS ;
	wire \mchip.pong.btn_rst ;
	wire \mchip.pong.btn_serve ;
	wire \mchip.pong.cfg1 ;
	wire \mchip.pong.cfg1_o ;
	wire \mchip.pong.cfg2 ;
	wire \mchip.pong.cfg2_o ;
	wire \mchip.pong.clk_25mhz ;
	wire \mchip.pong.game.Cnewgame ;
	wire [7:0] \mchip.pong.game.VGA_B ;
	wire [7:0] \mchip.pong.game.VGA_G ;
	wire \mchip.pong.game.VGA_HS ;
	wire [7:0] \mchip.pong.game.VGA_R ;
	wire \mchip.pong.game.VGA_VS ;
	wire \mchip.pong.game.ball.Cnewgame ;
	wire [9:0] \mchip.pong.game.ball.ballX ;
	wire [8:0] \mchip.pong.game.ball.ballY ;
	wire \mchip.pong.game.ball.clock ;
	wire \mchip.pong.game.ball.cpath.Cnewgame ;
	wire \mchip.pong.game.ball.cpath.clock ;
	wire \mchip.pong.game.ball.cpath.reset ;
	wire \mchip.pong.game.ball.cpath.serve_input ;
	reg [8:0] \mchip.pong.game.ball.cpath.state ;
	wire \mchip.pong.game.ball.dpath.Cnewgame ;
	wire [9:0] \mchip.pong.game.ball.dpath.ballX ;
	reg [8:0] \mchip.pong.game.ball.dpath.ballY ;
	wire \mchip.pong.game.ball.dpath.clock ;
	wire \mchip.pong.game.ball.dpath.en_pos_reg ;
	wire [9:0] \mchip.pong.game.ball.dpath.nextX ;
	wire [8:0] \mchip.pong.game.ball.dpath.nextY ;
	wire [8:0] \mchip.pong.game.ball.dpath.paddleLY ;
	wire [8:0] \mchip.pong.game.ball.dpath.paddleRY ;
	wire [8:0] \mchip.pong.game.ball.paddleLY ;
	wire [8:0] \mchip.pong.game.ball.paddleRY ;
	wire \mchip.pong.game.ball.reset ;
	wire \mchip.pong.game.ball.serve_input ;
	wire [9:0] \mchip.pong.game.ballX ;
	wire [8:0] \mchip.pong.game.ballY ;
	wire \mchip.pong.game.cfg1 ;
	wire \mchip.pong.game.cfg2 ;
	wire \mchip.pong.game.clock ;
	wire \mchip.pong.game.left_movedir ;
	wire \mchip.pong.game.left_paddle.Cnewgame ;
	wire \mchip.pong.game.left_paddle.clock ;
	reg [8:0] \mchip.pong.game.left_paddle.coord ;
	wire \mchip.pong.game.left_paddle.movedir_input ;
	wire [8:0] \mchip.pong.game.left_paddle.next_coord ;
	wire [8:0] \mchip.pong.game.paddleLY ;
	wire [8:0] \mchip.pong.game.paddleRY ;
	wire [23:0] \mchip.pong.game.renderer.ball.color ;
	wire [23:0] \mchip.pong.game.renderer.ball1.color ;
	wire [23:0] \mchip.pong.game.renderer.ball2.color ;
	wire [9:0] \mchip.pong.game.renderer.ballX ;
	wire [8:0] \mchip.pong.game.renderer.ballY ;
	wire [23:0] \mchip.pong.game.renderer.ballrom_out ;
	wire [23:0] \mchip.pong.game.renderer.ballrom_out0 ;
	wire [23:0] \mchip.pong.game.renderer.ballrom_out1 ;
	wire [23:0] \mchip.pong.game.renderer.ballrom_out2 ;
	wire \mchip.pong.game.renderer.cfg1 ;
	wire \mchip.pong.game.renderer.cfg2 ;
	wire [8:0] \mchip.pong.game.renderer.paddleLY ;
	wire [8:0] \mchip.pong.game.renderer.paddleRY ;
	wire [7:0] \mchip.pong.game.renderer.vga_b ;
	wire [9:0] \mchip.pong.game.renderer.vga_col ;
	wire [7:0] \mchip.pong.game.renderer.vga_g ;
	wire [7:0] \mchip.pong.game.renderer.vga_r ;
	wire \mchip.pong.game.reset ;
	wire \mchip.pong.game.right_movedir ;
	wire \mchip.pong.game.right_paddle.Cnewgame ;
	wire \mchip.pong.game.right_paddle.clock ;
	reg [8:0] \mchip.pong.game.right_paddle.coord ;
	wire \mchip.pong.game.right_paddle.movedir_input ;
	wire [8:0] \mchip.pong.game.right_paddle.next_coord ;
	wire \mchip.pong.game.score.Cnewgame ;
	wire \mchip.pong.game.score.clock ;
	wire [15:0] \mchip.pong.game.score.lscore_adder.B ;
	wire [3:0] \mchip.pong.game.score.lscore_adder.add0.B ;
	wire \mchip.pong.game.score.lscore_adder.add0.Cin ;
	wire [3:0] \mchip.pong.game.score.lscore_adder.add1.B ;
	wire [3:0] \mchip.pong.game.score.lscore_adder.add2.B ;
	wire [3:0] \mchip.pong.game.score.lscore_adder.add3.B ;
	wire [15:0] \mchip.pong.game.score.rscore_adder.B ;
	wire [3:0] \mchip.pong.game.score.rscore_adder.add0.B ;
	wire \mchip.pong.game.score.rscore_adder.add0.Cin ;
	wire [3:0] \mchip.pong.game.score.rscore_adder.add1.B ;
	wire [3:0] \mchip.pong.game.score.rscore_adder.add2.B ;
	wire [3:0] \mchip.pong.game.score.rscore_adder.add3.B ;
	wire \mchip.pong.game.serve_input ;
	wire \mchip.pong.game.tick.clock ;
	wire [9:0] \mchip.pong.game.tick.col ;
	wire \mchip.pong.game.vga.HS ;
	wire \mchip.pong.game.vga.VS ;
	wire \mchip.pong.game.vga.clock ;
	wire [9:0] \mchip.pong.game.vga.col ;
	reg [9:0] \mchip.pong.game.vga.line_ind ;
	reg \mchip.pong.game.vga.pclk_ctr ;
	reg [9:0] \mchip.pong.game.vga.pix_ind ;
	wire \mchip.pong.game.vga.reset ;
	wire [9:0] \mchip.pong.game.vga_col ;
	wire \mchip.pong.left_down ;
	wire \mchip.pong.left_up ;
	wire \mchip.pong.right_down ;
	wire \mchip.pong.right_up ;
	wire \mchip.pong.rst ;
	wire \mchip.pong.serve ;
	wire \mchip.pong.sync.i_clk ;
	wire [7:0] \mchip.pong.sync.i_in ;
	wire \mchip.pong.sync.i_rst ;
	reg [7:0] \mchip.pong.sync.o_out  = 8'h00;
	reg [7:0] \mchip.pong.sync.sync  = 8'h00;
	wire \mchip.reset ;
	assign \mchip.pong.game.left_paddle.next_coord [0] = ~\mchip.pong.game.left_paddle.coord [0];
	assign _0589_ = \mchip.pong.game.left_paddle.coord [3] & \mchip.pong.sync.o_out [7];
	assign _0600_ = \mchip.pong.game.left_paddle.coord [2] & ~\mchip.pong.sync.o_out [7];
	assign _0611_ = \mchip.pong.game.left_paddle.coord [3] ^ \mchip.pong.sync.o_out [7];
	assign _0622_ = _0611_ & _0600_;
	assign _0633_ = _0622_ | _0589_;
	assign _0644_ = ~(\mchip.pong.game.left_paddle.coord [2] ^ \mchip.pong.sync.o_out [7]);
	assign _0655_ = _0644_ & _0611_;
	assign _0666_ = ~(\mchip.pong.game.left_paddle.coord [1] & \mchip.pong.sync.o_out [7]);
	assign _0677_ = \mchip.pong.game.left_paddle.coord [1] ^ \mchip.pong.sync.o_out [7];
	assign _0688_ = _0677_ & ~\mchip.pong.game.left_paddle.next_coord [0];
	assign _0699_ = _0666_ & ~_0688_;
	assign _0710_ = _0655_ & ~_0699_;
	assign _0721_ = _0710_ | _0633_;
	assign _0732_ = \mchip.pong.game.left_paddle.coord [4] ^ \mchip.pong.sync.o_out [7];
	assign \mchip.pong.game.left_paddle.next_coord [4] = _0732_ ^ _0721_;
	assign _0753_ = \mchip.pong.game.left_paddle.coord [4] & \mchip.pong.sync.o_out [7];
	assign _0764_ = _0732_ & _0721_;
	assign _0775_ = ~(_0764_ | _0753_);
	assign _0786_ = \mchip.pong.game.left_paddle.coord [5] ^ \mchip.pong.sync.o_out [7];
	assign \mchip.pong.game.left_paddle.next_coord [5] = ~(_0786_ ^ _0775_);
	assign _0807_ = \mchip.pong.game.right_paddle.coord [4] & \mchip.pong.sync.o_out [5];
	assign _0818_ = \mchip.pong.game.right_paddle.coord [4] ^ \mchip.pong.sync.o_out [5];
	assign _0829_ = ~(\mchip.pong.game.right_paddle.coord [3] & \mchip.pong.sync.o_out [5]);
	assign _0840_ = \mchip.pong.game.right_paddle.coord [2] & ~\mchip.pong.sync.o_out [5];
	assign _0851_ = \mchip.pong.game.right_paddle.coord [3] ^ \mchip.pong.sync.o_out [5];
	assign _0862_ = _0851_ & _0840_;
	assign _0873_ = _0829_ & ~_0862_;
	assign _0884_ = ~(\mchip.pong.game.right_paddle.coord [2] ^ \mchip.pong.sync.o_out [5]);
	assign _0895_ = _0884_ & _0851_;
	assign _0906_ = ~(\mchip.pong.game.right_paddle.coord [1] & \mchip.pong.sync.o_out [5]);
	assign \mchip.pong.game.right_paddle.next_coord [0] = ~\mchip.pong.game.right_paddle.coord [0];
	assign _0927_ = \mchip.pong.game.right_paddle.coord [1] ^ \mchip.pong.sync.o_out [5];
	assign _0938_ = _0927_ & ~\mchip.pong.game.right_paddle.next_coord [0];
	assign _0949_ = _0906_ & ~_0938_;
	assign _0960_ = _0895_ & ~_0949_;
	assign _0971_ = _0873_ & ~_0960_;
	assign _0982_ = _0818_ & ~_0971_;
	assign _0993_ = ~(_0982_ | _0807_);
	assign _1004_ = \mchip.pong.sync.o_out [5] ^ \mchip.pong.game.right_paddle.coord [5];
	assign \mchip.pong.game.right_paddle.next_coord [5] = ~(_1004_ ^ _0993_);
	assign \mchip.pong.game.right_paddle.next_coord [4] = ~(_0971_ ^ _0818_);
	assign _4446_ = ~\mchip.pong.game.vga.pclk_ctr ;
	assign _1045_ = \mchip.pong.game.vga.line_ind [0] & \mchip.pong.game.vga.line_ind [1];
	assign _1056_ = \mchip.pong.game.vga.line_ind [2] | \mchip.pong.game.vga.line_ind [3];
	assign _1067_ = _1056_ | _1045_;
	assign _1078_ = \mchip.pong.game.vga.line_ind [4] | \mchip.pong.game.vga.line_ind [5];
	assign _1089_ = \mchip.pong.game.vga.line_ind [6] | \mchip.pong.game.vga.line_ind [7];
	assign _1100_ = _1089_ | _1078_;
	assign _1111_ = ~(_1100_ | _1067_);
	assign _1122_ = ~(\mchip.pong.game.vga.line_ind [9] | \mchip.pong.game.vga.line_ind [8]);
	assign _1133_ = ~(_1122_ & _1111_);
	assign _1144_ = \mchip.pong.game.vga.line_ind [1] & ~\mchip.pong.game.vga.line_ind [0];
	assign _1155_ = _1056_ | ~_1144_;
	assign _1166_ = _1155_ | _1100_;
	assign _1177_ = _1122_ & ~_1166_;
	assign \mchip.pong.VGA_VS  = _1177_ | _1133_;
	assign \mchip.pong.game.ball.dpath.nextY [0] = ~\mchip.pong.game.ball.dpath.ballY [0];
	assign _1208_ = ~\mchip.pong.sync.o_out [2];
	assign _1219_ = \mchip.pong.game.ball.dpath.ballX [9] & ~\mchip.pong.game.ball.dpath.ballX [8];
	assign _1230_ = ~(\mchip.pong.game.ball.dpath.ballX [7] | \mchip.pong.game.ball.dpath.ballX [6]);
	assign _1241_ = ~(\mchip.pong.game.ball.dpath.ballX [5] | \mchip.pong.game.ball.dpath.ballX [4]);
	assign _1252_ = _1241_ & _1230_;
	assign \mchip.pong.game.ball.dpath.nextX [1] = ~\mchip.pong.game.ball.dpath.ballX [1];
	assign _1283_ = \mchip.pong.game.ball.dpath.ballX [2] | \mchip.pong.game.ball.dpath.ballX [3];
	assign _1294_ = \mchip.pong.game.ball.dpath.nextX [1] & ~_1283_;
	assign _1305_ = _1252_ & ~_1294_;
	assign _1316_ = _1252_ & ~_1305_;
	assign _1327_ = _1219_ & ~_1316_;
	assign _1338_ = \mchip.pong.game.ball.dpath.ballX [8] & \mchip.pong.game.ball.dpath.ballX [9];
	assign _1349_ = _1338_ | _1327_;
	assign _1360_ = \mchip.pong.game.ball.dpath.ballX [1] | ~\mchip.pong.game.ball.dpath.ballX [9];
	assign _1371_ = \mchip.pong.game.ball.dpath.ballX [5] | ~\mchip.pong.game.ball.dpath.ballX [6];
	assign _1382_ = \mchip.pong.game.ball.dpath.ballX [8] | \mchip.pong.game.ball.dpath.ballX [7];
	assign _1393_ = _1382_ | _1371_;
	assign _1404_ = \mchip.pong.game.ball.dpath.ballX [4] | \mchip.pong.game.ball.dpath.ballX [3];
	assign _1415_ = _1404_ | \mchip.pong.game.ball.dpath.ballX [2];
	assign _1426_ = _1415_ | _1393_;
	assign _1437_ = _1426_ | _1360_;
	assign _1448_ = _1230_ | ~_1219_;
	assign _1459_ = _1448_ & ~_1338_;
	assign _1470_ = _1437_ & ~_1459_;
	assign _1481_ = _1349_ & ~_1470_;
	assign _1492_ = \mchip.pong.game.ball.dpath.ballY [7] & \mchip.pong.game.ball.dpath.ballY [6];
	assign _1503_ = ~(\mchip.pong.game.ball.dpath.ballY [5] | \mchip.pong.game.ball.dpath.ballY [4]);
	assign _1514_ = _1503_ | ~_1492_;
	assign _1523_ = _1503_ & _1492_;
	assign _1534_ = ~(\mchip.pong.game.ball.dpath.ballY [3] | \mchip.pong.game.ball.dpath.ballY [2]);
	assign _1545_ = ~(\mchip.pong.game.ball.dpath.ballY [1] | \mchip.pong.game.ball.dpath.ballY [0]);
	assign _1556_ = _1545_ & _1534_;
	assign _1567_ = _1523_ & ~_1556_;
	assign _1578_ = _1514_ & ~_1567_;
	assign _1589_ = \mchip.pong.game.ball.dpath.ballY [8] & ~_1578_;
	assign _1600_ = ~_1589_;
	assign _1611_ = ~\mchip.pong.game.ball.dpath.ballY [8];
	assign _1622_ = _1578_ ^ _1611_;
	assign _1633_ = _1622_ ^ \mchip.pong.game.right_paddle.coord [8];
	assign _1643_ = _1600_ & ~_1633_;
	assign _1654_ = ~\mchip.pong.game.right_paddle.coord [5];
	assign _1665_ = _1556_ & ~\mchip.pong.game.ball.dpath.ballY [4];
	assign _1675_ = _1665_ ^ \mchip.pong.game.ball.dpath.ballY [5];
	assign _1686_ = _1675_ ^ _1654_;
	assign _1697_ = _1556_ ^ \mchip.pong.game.ball.dpath.ballY [4];
	assign _1707_ = _1697_ ^ \mchip.pong.game.right_paddle.coord [4];
	assign _1718_ = _1686_ & ~_1707_;
	assign _1728_ = ~\mchip.pong.game.right_paddle.coord [6];
	assign _1739_ = ~\mchip.pong.game.ball.dpath.ballY [6];
	assign _1750_ = _1556_ & _1503_;
	assign _1761_ = _1750_ ^ _1739_;
	assign _1772_ = _1761_ ^ _1728_;
	assign _1783_ = ~\mchip.pong.game.right_paddle.coord [7];
	assign _1794_ = \mchip.pong.game.ball.dpath.ballY [6] & ~_1750_;
	assign _1805_ = _1794_ ^ \mchip.pong.game.ball.dpath.ballY [7];
	assign _1816_ = _1805_ ^ _1783_;
	assign _1827_ = _1816_ & _1772_;
	assign _1838_ = _1827_ & _1718_;
	assign _1849_ = ~\mchip.pong.game.right_paddle.coord [3];
	assign _1860_ = _1545_ & ~\mchip.pong.game.ball.dpath.ballY [2];
	assign _1871_ = _1860_ ^ \mchip.pong.game.ball.dpath.ballY [3];
	assign _1882_ = _1871_ ^ _1849_;
	assign _1893_ = _1545_ ^ \mchip.pong.game.ball.dpath.ballY [2];
	assign _1904_ = _1893_ ^ \mchip.pong.game.right_paddle.coord [2];
	assign _1915_ = _1882_ & ~_1904_;
	assign _1926_ = ~\mchip.pong.game.right_paddle.coord [1];
	assign _1937_ = ~(\mchip.pong.game.ball.dpath.ballY [1] ^ \mchip.pong.game.ball.dpath.ballY [0]);
	assign _1948_ = _1937_ ^ _1926_;
	assign _1958_ = ~(\mchip.pong.game.ball.dpath.ballY [0] ^ \mchip.pong.game.right_paddle.coord [0]);
	assign _1969_ = _1948_ & ~_1958_;
	assign _1980_ = _1969_ & _1915_;
	assign _1991_ = _1980_ & _1838_;
	assign _2002_ = ~(_1991_ & _1643_);
	assign _2013_ = ~\mchip.pong.game.right_paddle.coord [8];
	assign _2024_ = _1622_ | _2013_;
	assign _2035_ = _2024_ | _1589_;
	assign _2046_ = _1805_ | _1783_;
	assign _2067_ = _1761_ | _1728_;
	assign _2078_ = _1816_ & ~_2067_;
	assign _2089_ = _2046_ & ~_2078_;
	assign _2100_ = _1675_ | _1654_;
	assign _2111_ = ~\mchip.pong.game.right_paddle.coord [4];
	assign _2122_ = _1697_ | _2111_;
	assign _2133_ = _1686_ & ~_2122_;
	assign _2144_ = _2100_ & ~_2133_;
	assign _2155_ = _1827_ & ~_2144_;
	assign _2166_ = _2089_ & ~_2155_;
	assign _2177_ = _1871_ | _1849_;
	assign _2188_ = ~\mchip.pong.game.right_paddle.coord [2];
	assign _2199_ = _1893_ | _2188_;
	assign _2210_ = _1882_ & ~_2199_;
	assign _2221_ = _2177_ & ~_2210_;
	assign _2232_ = _1937_ | _1926_;
	assign _2243_ = ~(\mchip.pong.game.ball.dpath.ballY [0] | \mchip.pong.game.right_paddle.coord [0]);
	assign _2253_ = _1948_ & ~_2243_;
	assign _2264_ = _2232_ & ~_2253_;
	assign _2275_ = _1915_ & ~_2264_;
	assign _2286_ = _2221_ & ~_2275_;
	assign _2297_ = _1838_ & ~_2286_;
	assign _2308_ = _2166_ & ~_2297_;
	assign _2319_ = _1643_ & ~_2308_;
	assign _2330_ = _2035_ & ~_2319_;
	assign _2341_ = _2002_ & ~_2330_;
	assign _2352_ = \mchip.pong.game.right_paddle.coord [7] & \mchip.pong.game.right_paddle.coord [6];
	assign _2363_ = ~(\mchip.pong.game.right_paddle.coord [4] & \mchip.pong.game.right_paddle.coord [5]);
	assign _2374_ = _2363_ | ~_2352_;
	assign _2384_ = \mchip.pong.game.right_paddle.coord [5] & ~\mchip.pong.game.right_paddle.coord [4];
	assign _2395_ = _2384_ & _2352_;
	assign _2405_ = ~(\mchip.pong.game.right_paddle.coord [2] & \mchip.pong.game.right_paddle.coord [3]);
	assign _2416_ = \mchip.pong.game.right_paddle.coord [0] | \mchip.pong.game.right_paddle.coord [1];
	assign _2427_ = \mchip.pong.game.right_paddle.coord [2] | ~\mchip.pong.game.right_paddle.coord [3];
	assign _2438_ = _2416_ & ~_2427_;
	assign _2449_ = _2405_ & ~_2438_;
	assign _2460_ = _2395_ & ~_2449_;
	assign _2471_ = _2374_ & ~_2460_;
	assign _2482_ = \mchip.pong.game.right_paddle.coord [8] & ~_2471_;
	assign _2493_ = ~_2482_;
	assign _2504_ = _2471_ ^ _2013_;
	assign _2515_ = _2504_ ^ \mchip.pong.game.ball.dpath.ballY [8];
	assign _2526_ = _2493_ & ~_2515_;
	assign _2537_ = _2384_ & ~_2449_;
	assign _2548_ = _2363_ & ~_2537_;
	assign _2559_ = \mchip.pong.game.right_paddle.coord [6] & ~_2548_;
	assign _2570_ = _2559_ ^ _1783_;
	assign _2581_ = _2570_ ^ \mchip.pong.game.ball.dpath.ballY [7];
	assign _2592_ = _2548_ ^ _1728_;
	assign _2603_ = _2592_ ^ \mchip.pong.game.ball.dpath.ballY [6];
	assign _2614_ = _2581_ & ~_2603_;
	assign _2625_ = ~\mchip.pong.game.ball.dpath.ballY [4];
	assign _2636_ = _2449_ ^ \mchip.pong.game.right_paddle.coord [4];
	assign _2647_ = _2636_ ^ _2625_;
	assign _2658_ = ~\mchip.pong.game.ball.dpath.ballY [5];
	assign _2669_ = _2449_ & ~\mchip.pong.game.right_paddle.coord [4];
	assign _2680_ = _2669_ ^ _1654_;
	assign _2691_ = _2680_ ^ _2658_;
	assign _2701_ = ~(_2691_ & _2647_);
	assign _2712_ = _2614_ & ~_2701_;
	assign _2723_ = _2188_ & ~_2416_;
	assign _2734_ = _2723_ ^ \mchip.pong.game.right_paddle.coord [3];
	assign _2745_ = _2734_ ^ \mchip.pong.game.ball.dpath.ballY [3];
	assign _2756_ = _2416_ ^ _2188_;
	assign _2767_ = _2756_ ^ \mchip.pong.game.ball.dpath.ballY [2];
	assign _2778_ = _2745_ & ~_2767_;
	assign _2789_ = ~(\mchip.pong.game.right_paddle.coord [0] ^ \mchip.pong.game.right_paddle.coord [1]);
	assign _2800_ = _2789_ ^ \mchip.pong.game.ball.dpath.ballY [1];
	assign _2811_ = ~(_2800_ | _1958_);
	assign _2822_ = _2811_ & _2778_;
	assign _2833_ = _2822_ & _2712_;
	assign _2844_ = ~(_2833_ & _2526_);
	assign _2855_ = _2504_ | _1611_;
	assign _2866_ = _2855_ | _2482_;
	assign _2877_ = ~\mchip.pong.game.ball.dpath.ballY [7];
	assign _2888_ = _2559_ ^ \mchip.pong.game.right_paddle.coord [7];
	assign _2899_ = _2888_ | _2877_;
	assign _2920_ = _2592_ | _1739_;
	assign _2931_ = _2581_ & ~_2920_;
	assign _2942_ = _2899_ & ~_2931_;
	assign _2953_ = _2680_ | _2658_;
	assign _2963_ = _2636_ | _2625_;
	assign _2974_ = _2691_ & ~_2963_;
	assign _2985_ = _2953_ & ~_2974_;
	assign _2996_ = _2614_ & ~_2985_;
	assign _3007_ = _2942_ & ~_2996_;
	assign _3018_ = ~(_2734_ & \mchip.pong.game.ball.dpath.ballY [3]);
	assign _3029_ = ~\mchip.pong.game.ball.dpath.ballY [2];
	assign _3040_ = _2756_ | _3029_;
	assign _3051_ = _2745_ & ~_3040_;
	assign _3062_ = _3018_ & ~_3051_;
	assign _3073_ = ~\mchip.pong.game.ball.dpath.ballY [1];
	assign _3084_ = _2789_ | _3073_;
	assign _3095_ = ~(_2800_ | _2243_);
	assign _3106_ = _3084_ & ~_3095_;
	assign _3117_ = _2778_ & ~_3106_;
	assign _3128_ = _3062_ & ~_3117_;
	assign _3139_ = _2712_ & ~_3128_;
	assign _3150_ = _3007_ & ~_3139_;
	assign _3161_ = _2526_ & ~_3150_;
	assign _3172_ = _2866_ & ~_3161_;
	assign _3183_ = _2844_ & ~_3172_;
	assign _3194_ = _3183_ | _2341_;
	assign _3205_ = _1481_ & ~_3194_;
	assign _3216_ = ~(_3205_ & _1208_);
	assign _3227_ = \mchip.pong.game.ball.cpath.state [5] & ~_3216_;
	assign _3238_ = \mchip.pong.sync.o_out [3] & ~\mchip.pong.sync.o_out [2];
	assign _3249_ = _3238_ & \mchip.pong.game.ball.cpath.state [4];
	assign _3260_ = _3249_ | _3227_;
	assign _3271_ = ~\mchip.pong.game.ball.dpath.ballX [7];
	assign _3282_ = \mchip.pong.game.ball.dpath.ballX [6] & ~\mchip.pong.game.ball.dpath.ballX [7];
	assign _3293_ = \mchip.pong.game.ball.dpath.ballX [5] & \mchip.pong.game.ball.dpath.ballX [4];
	assign _3304_ = _3293_ & _3282_;
	assign _3315_ = ~(\mchip.pong.game.ball.dpath.ballX [2] & \mchip.pong.game.ball.dpath.ballX [3]);
	assign _3326_ = _3304_ & ~_3315_;
	assign _3337_ = _3271_ & ~_3326_;
	assign _3348_ = _1219_ & ~_3337_;
	assign _3359_ = ~(_3348_ | _1338_);
	assign _3370_ = ~\mchip.pong.game.ball.dpath.ballX [9];
	assign _3381_ = ~(\mchip.pong.game.ball.dpath.ballX [1] | \mchip.pong.game.ball.dpath.ballX [2]);
	assign _3392_ = _1404_ | ~_3381_;
	assign _3403_ = \mchip.pong.game.ball.dpath.ballX [5] | \mchip.pong.game.ball.dpath.ballX [6];
	assign _3414_ = _3403_ | _1382_;
	assign _3425_ = _3414_ | _3392_;
	assign _3436_ = _3370_ & ~_3425_;
	assign _3447_ = _3359_ & ~_3436_;
	assign _3458_ = ~_3447_;
	assign _3469_ = _3293_ | ~_1230_;
	assign _3480_ = _3315_ | \mchip.pong.game.ball.dpath.nextX [1];
	assign _3491_ = ~(_3293_ & _1230_);
	assign _3501_ = _3480_ & ~_3491_;
	assign _3512_ = _3501_ | ~_3469_;
	assign _3523_ = ~(\mchip.pong.game.ball.dpath.ballX [8] | \mchip.pong.game.ball.dpath.ballX [9]);
	assign _3534_ = ~(_3523_ & _3512_);
	assign _3545_ = _3315_ | \mchip.pong.game.ball.dpath.ballX [1];
	assign _3556_ = _3491_ | _3545_;
	assign _3567_ = _3523_ & ~_3556_;
	assign _3578_ = _3567_ | _3534_;
	assign _3588_ = ~(_3523_ & _1230_);
	assign _3599_ = _3523_ & _3282_;
	assign _3610_ = _1283_ | ~_1241_;
	assign _3621_ = _3599_ & ~_3610_;
	assign _3632_ = _3588_ & ~_3621_;
	assign _3643_ = _3578_ & ~_3632_;
	assign _3654_ = _1622_ ^ \mchip.pong.game.left_paddle.coord [8];
	assign _3665_ = _1600_ & ~_3654_;
	assign _3676_ = ~\mchip.pong.game.left_paddle.coord [7];
	assign _3687_ = _1805_ ^ _3676_;
	assign _3698_ = _1761_ ^ \mchip.pong.game.left_paddle.coord [6];
	assign _3709_ = _3687_ & ~_3698_;
	assign _3720_ = ~\mchip.pong.game.left_paddle.coord [4];
	assign _3731_ = _1697_ ^ _3720_;
	assign _3742_ = ~\mchip.pong.game.left_paddle.coord [5];
	assign _3753_ = _1675_ ^ _3742_;
	assign _3764_ = ~(_3753_ & _3731_);
	assign _3775_ = _3709_ & ~_3764_;
	assign _3786_ = ~\mchip.pong.game.left_paddle.coord [3];
	assign _3797_ = _1871_ ^ _3786_;
	assign _3808_ = _1893_ ^ \mchip.pong.game.left_paddle.coord [2];
	assign _3819_ = _3797_ & ~_3808_;
	assign _3830_ = ~\mchip.pong.game.left_paddle.coord [1];
	assign _3841_ = _1937_ ^ _3830_;
	assign _3852_ = ~(\mchip.pong.game.ball.dpath.ballY [0] ^ \mchip.pong.game.left_paddle.coord [0]);
	assign _3863_ = _3841_ & ~_3852_;
	assign _3873_ = _3863_ & _3819_;
	assign _3880_ = _3873_ & _3775_;
	assign _3890_ = ~(_3880_ & _3665_);
	assign _3899_ = ~\mchip.pong.game.left_paddle.coord [8];
	assign _3909_ = _1622_ | _3899_;
	assign _3919_ = _3909_ | _1589_;
	assign _3936_ = _1805_ | _3676_;
	assign _3945_ = ~\mchip.pong.game.left_paddle.coord [6];
	assign _3954_ = _1761_ | _3945_;
	assign _3965_ = _3687_ & ~_3954_;
	assign _3966_ = _3936_ & ~_3965_;
	assign _3967_ = _1675_ | _3742_;
	assign _3968_ = _1697_ | _3720_;
	assign _3969_ = _3753_ & ~_3968_;
	assign _3970_ = _3967_ & ~_3969_;
	assign _3971_ = _3709_ & ~_3970_;
	assign _3972_ = _3966_ & ~_3971_;
	assign _3973_ = _1871_ | _3786_;
	assign _3974_ = ~\mchip.pong.game.left_paddle.coord [2];
	assign _3975_ = _1893_ | _3974_;
	assign _3976_ = _3797_ & ~_3975_;
	assign _3977_ = _3973_ & ~_3976_;
	assign _3978_ = _1937_ | _3830_;
	assign _3979_ = ~(\mchip.pong.game.ball.dpath.ballY [0] | \mchip.pong.game.left_paddle.coord [0]);
	assign _3980_ = _3841_ & ~_3979_;
	assign _3981_ = _3978_ & ~_3980_;
	assign _3982_ = _3819_ & ~_3981_;
	assign _3983_ = _3977_ & ~_3982_;
	assign _3984_ = _3775_ & ~_3983_;
	assign _3985_ = _3972_ & ~_3984_;
	assign _3986_ = _3665_ & ~_3985_;
	assign _3987_ = _3919_ & ~_3986_;
	assign _3988_ = _3890_ & ~_3987_;
	assign _3989_ = \mchip.pong.game.left_paddle.coord [7] & \mchip.pong.game.left_paddle.coord [6];
	assign _3990_ = ~(\mchip.pong.game.left_paddle.coord [5] & \mchip.pong.game.left_paddle.coord [4]);
	assign _3991_ = _3990_ | ~_3989_;
	assign _3992_ = \mchip.pong.game.left_paddle.coord [5] & ~\mchip.pong.game.left_paddle.coord [4];
	assign _3993_ = _3992_ & _3989_;
	assign _3994_ = ~(\mchip.pong.game.left_paddle.coord [2] & \mchip.pong.game.left_paddle.coord [3]);
	assign _3995_ = \mchip.pong.game.left_paddle.coord [1] | \mchip.pong.game.left_paddle.coord [0];
	assign _3996_ = \mchip.pong.game.left_paddle.coord [2] | ~\mchip.pong.game.left_paddle.coord [3];
	assign _3997_ = _3995_ & ~_3996_;
	assign _3998_ = _3994_ & ~_3997_;
	assign _3999_ = _3993_ & ~_3998_;
	assign _4000_ = _3991_ & ~_3999_;
	assign _4001_ = \mchip.pong.game.left_paddle.coord [8] & ~_4000_;
	assign _4002_ = ~_4001_;
	assign _4003_ = _4000_ ^ _3899_;
	assign _4004_ = _4003_ ^ \mchip.pong.game.ball.dpath.ballY [8];
	assign _4005_ = _4002_ & ~_4004_;
	assign _4006_ = _3992_ & ~_3998_;
	assign _4007_ = _3990_ & ~_4006_;
	assign _4008_ = \mchip.pong.game.left_paddle.coord [6] & ~_4007_;
	assign _4009_ = _4008_ ^ _3676_;
	assign _4010_ = _4009_ ^ \mchip.pong.game.ball.dpath.ballY [7];
	assign _4011_ = _4007_ ^ _3945_;
	assign _4012_ = _4011_ ^ \mchip.pong.game.ball.dpath.ballY [6];
	assign _4013_ = _4010_ & ~_4012_;
	assign _4014_ = _3998_ ^ \mchip.pong.game.left_paddle.coord [4];
	assign _4015_ = _4014_ ^ _2625_;
	assign _4016_ = _3998_ & ~\mchip.pong.game.left_paddle.coord [4];
	assign _4017_ = _4016_ ^ _3742_;
	assign _4018_ = _4017_ ^ _2658_;
	assign _4019_ = ~(_4018_ & _4015_);
	assign _4020_ = _4013_ & ~_4019_;
	assign _4021_ = _3974_ & ~_3995_;
	assign _4022_ = _4021_ ^ \mchip.pong.game.left_paddle.coord [3];
	assign _4023_ = _4022_ ^ \mchip.pong.game.ball.dpath.ballY [3];
	assign _4024_ = _3995_ ^ _3974_;
	assign _4025_ = _4024_ ^ \mchip.pong.game.ball.dpath.ballY [2];
	assign _4026_ = _4023_ & ~_4025_;
	assign _4027_ = ~(\mchip.pong.game.left_paddle.coord [1] ^ \mchip.pong.game.left_paddle.coord [0]);
	assign _4028_ = _4027_ ^ \mchip.pong.game.ball.dpath.ballY [1];
	assign _4029_ = ~(_4028_ | _3852_);
	assign _4030_ = _4029_ & _4026_;
	assign _4031_ = _4030_ & _4020_;
	assign _4032_ = ~(_4031_ & _4005_);
	assign _4033_ = _4003_ | _1611_;
	assign _4034_ = _4033_ | _4001_;
	assign _4035_ = _4008_ ^ \mchip.pong.game.left_paddle.coord [7];
	assign _4036_ = _4035_ | _2877_;
	assign _4037_ = _4011_ | _1739_;
	assign _4038_ = _4010_ & ~_4037_;
	assign _4039_ = _4036_ & ~_4038_;
	assign _4040_ = _4017_ | _2658_;
	assign _4041_ = _4014_ | _2625_;
	assign _4042_ = _4018_ & ~_4041_;
	assign _4043_ = _4040_ & ~_4042_;
	assign _4044_ = _4013_ & ~_4043_;
	assign _4045_ = _4039_ & ~_4044_;
	assign _4046_ = ~(_4022_ & \mchip.pong.game.ball.dpath.ballY [3]);
	assign _4047_ = _4024_ | _3029_;
	assign _4048_ = _4023_ & ~_4047_;
	assign _4049_ = _4046_ & ~_4048_;
	assign _4050_ = _4027_ | _3073_;
	assign _4051_ = ~(_4028_ | _3979_);
	assign _4052_ = _4050_ & ~_4051_;
	assign _4053_ = _4026_ & ~_4052_;
	assign _4054_ = _4049_ & ~_4053_;
	assign _4055_ = _4020_ & ~_4054_;
	assign _4056_ = _4045_ & ~_4055_;
	assign _4057_ = _4005_ & ~_4056_;
	assign _4058_ = _4034_ & ~_4057_;
	assign _4059_ = _4032_ & ~_4058_;
	assign _4060_ = _4059_ | _3988_;
	assign _4061_ = _3643_ & ~_4060_;
	assign _4062_ = _4061_ | _3458_;
	assign _4063_ = \mchip.pong.game.ball.dpath.ballY [6] | ~\mchip.pong.game.ball.dpath.ballY [7];
	assign _4064_ = _4063_ | _2658_;
	assign _4065_ = _4064_ & ~_1492_;
	assign _4066_ = \mchip.pong.game.ball.dpath.ballY [5] | ~\mchip.pong.game.ball.dpath.ballY [4];
	assign _4067_ = ~(_4066_ | _4063_);
	assign _4068_ = ~(\mchip.pong.game.ball.dpath.ballY [3] & \mchip.pong.game.ball.dpath.ballY [2]);
	assign _4069_ = ~(\mchip.pong.game.ball.dpath.ballY [1] & \mchip.pong.game.ball.dpath.ballY [0]);
	assign _4070_ = _4069_ | _4068_;
	assign _4071_ = _4067_ & ~_4070_;
	assign _4072_ = _4065_ & ~_4071_;
	assign _4073_ = \mchip.pong.game.ball.dpath.ballY [8] & ~_4072_;
	assign _4074_ = _4071_ & ~_1611_;
	assign _4075_ = _4073_ & ~_4074_;
	assign _4076_ = _4075_ | \mchip.pong.sync.o_out [2];
	assign _4077_ = _4076_ | _4062_;
	assign _4078_ = \mchip.pong.game.ball.cpath.state [7] & ~_4077_;
	assign _4079_ = \mchip.pong.game.ball.dpath.ballY [8] | \mchip.pong.game.ball.dpath.ballY [7];
	assign _4080_ = \mchip.pong.game.ball.dpath.ballY [5] | \mchip.pong.game.ball.dpath.ballY [6];
	assign _4081_ = _4080_ | _4079_;
	assign _4082_ = \mchip.pong.game.ball.dpath.ballY [3] | \mchip.pong.game.ball.dpath.ballY [4];
	assign _4083_ = \mchip.pong.game.ball.dpath.ballY [1] | \mchip.pong.game.ball.dpath.ballY [2];
	assign _4084_ = _4083_ | _4082_;
	assign _4085_ = _4084_ | _4081_;
	assign _4086_ = \mchip.pong.game.ball.dpath.nextY [0] & ~_4085_;
	assign _4087_ = ~(_4086_ & _1208_);
	assign _4088_ = _4087_ | _4061_;
	assign _4089_ = \mchip.pong.game.ball.cpath.state [2] & ~_4088_;
	assign _4090_ = _4089_ | _4078_;
	assign _0007_ = _4090_ | _3260_;
	assign _4091_ = _4086_ | \mchip.pong.sync.o_out [2];
	assign _4092_ = _3447_ | _3205_;
	assign _4093_ = _4092_ | _4091_;
	assign _4094_ = \mchip.pong.game.ball.cpath.state [3] & ~_4093_;
	assign _4095_ = _4092_ | _4076_;
	assign _4096_ = \mchip.pong.game.ball.cpath.state [5] & ~_4095_;
	assign _0008_ = _4096_ | _4094_;
	assign _4097_ = \mchip.pong.game.vga.pix_ind [9] & \mchip.pong.game.vga.pix_ind [8];
	assign _4098_ = ~(\mchip.pong.game.vga.pix_ind [6] | \mchip.pong.game.vga.pix_ind [7]);
	assign _4099_ = \mchip.pong.game.vga.pix_ind [4] & ~\mchip.pong.game.vga.pix_ind [5];
	assign _4100_ = _4099_ & _4098_;
	assign _4101_ = \mchip.pong.game.vga.pix_ind [3] & \mchip.pong.game.vga.pix_ind [2];
	assign _4102_ = \mchip.pong.game.vga.pix_ind [0] & \mchip.pong.game.vga.pix_ind [1];
	assign _4103_ = _4102_ & _4101_;
	assign _4104_ = ~(_4103_ & _4100_);
	assign _4105_ = _4104_ | ~_4097_;
	assign _0009_ = _4446_ & ~_4105_;
	assign _4106_ = _4061_ | _3447_;
	assign _4107_ = _4106_ | _4076_;
	assign _4108_ = \mchip.pong.game.ball.cpath.state [7] & ~_4107_;
	assign _4109_ = _4106_ | _4091_;
	assign _4110_ = \mchip.pong.game.ball.cpath.state [2] & ~_4109_;
	assign _0006_ = _4110_ | _4108_;
	assign _4111_ = ~(\mchip.pong.game.ball.cpath.state [0] | \mchip.pong.game.ball.cpath.state [1]);
	assign _4112_ = _3238_ & ~_4111_;
	assign _4113_ = _3458_ | _3205_;
	assign _4114_ = _4113_ | _4076_;
	assign _4115_ = \mchip.pong.game.ball.cpath.state [5] & ~_4114_;
	assign _4116_ = _4115_ | _4112_;
	assign _4117_ = _4087_ | _3205_;
	assign _4118_ = \mchip.pong.game.ball.cpath.state [3] & ~_4117_;
	assign _4119_ = ~(_4061_ & _1208_);
	assign _4120_ = \mchip.pong.game.ball.cpath.state [7] & ~_4119_;
	assign _4121_ = _4120_ | _4118_;
	assign _0005_ = _4121_ | _4116_;
	assign _4122_ = \mchip.pong.sync.o_out [3] | \mchip.pong.sync.o_out [2];
	assign _4123_ = \mchip.pong.game.ball.cpath.state [4] & ~_4122_;
	assign _4124_ = \mchip.pong.game.ball.cpath.state [6] & ~\mchip.pong.sync.o_out [2];
	assign _0004_ = _4124_ | _4123_;
	assign _4125_ = _0644_ & ~_0699_;
	assign _4126_ = _4125_ | _0600_;
	assign \mchip.pong.game.left_paddle.next_coord [3] = _4126_ ^ _0611_;
	assign _4127_ = \mchip.pong.game.left_paddle.coord [5] & \mchip.pong.sync.o_out [7];
	assign _4128_ = _0786_ & _0753_;
	assign _4129_ = _4128_ | _4127_;
	assign _4130_ = ~(_0786_ & _0732_);
	assign _4131_ = _0721_ & ~_4130_;
	assign _4132_ = _4131_ | _4129_;
	assign _4133_ = \mchip.pong.game.left_paddle.coord [6] ^ \mchip.pong.sync.o_out [7];
	assign \mchip.pong.game.left_paddle.next_coord [6] = _4133_ ^ _4132_;
	assign _4134_ = \mchip.pong.game.left_paddle.coord [6] & \mchip.pong.sync.o_out [7];
	assign _4135_ = _4133_ & _4132_;
	assign _4136_ = ~(_4135_ | _4134_);
	assign _4137_ = \mchip.pong.game.left_paddle.coord [7] ^ \mchip.pong.sync.o_out [7];
	assign \mchip.pong.game.left_paddle.next_coord [7] = ~(_4137_ ^ _4136_);
	assign _4138_ = \mchip.pong.game.left_paddle.coord [7] & \mchip.pong.sync.o_out [7];
	assign _4139_ = _4137_ & _4134_;
	assign _4140_ = ~(_4139_ | _4138_);
	assign _4141_ = ~(_4137_ & _4133_);
	assign _4142_ = _4129_ & ~_4141_;
	assign _4143_ = _4140_ & ~_4142_;
	assign _4144_ = _4141_ | _4130_;
	assign _4145_ = _0721_ & ~_4144_;
	assign _4146_ = _4143_ & ~_4145_;
	assign _4147_ = \mchip.pong.game.left_paddle.coord [8] ^ \mchip.pong.sync.o_out [7];
	assign \mchip.pong.game.left_paddle.next_coord [8] = ~(_4147_ ^ _4146_);
	assign _4148_ = \mchip.pong.game.ball.cpath.state [0] & ~_4122_;
	assign _0000_ = _4148_ | \mchip.pong.sync.o_out [2];
	assign _4149_ = \mchip.pong.game.ball.cpath.state [8] & ~\mchip.pong.sync.o_out [2];
	assign _4150_ = \mchip.pong.game.ball.cpath.state [1] & ~_4122_;
	assign _0001_ = _4150_ | _4149_;
	assign _4151_ = ~\mchip.pong.game.vga.pix_ind [5];
	assign _4152_ = \mchip.pong.game.vga.pix_ind [6] & ~\mchip.pong.game.vga.pix_ind [7];
	assign _4153_ = ~(_4152_ & _4151_);
	assign _4154_ = _4153_ & ~_4098_;
	assign _4155_ = \mchip.pong.game.vga.pix_ind [4] | ~\mchip.pong.game.vga.pix_ind [5];
	assign _4156_ = _4152_ & ~_4155_;
	assign _4157_ = ~(\mchip.pong.game.vga.pix_ind [0] | \mchip.pong.game.vga.pix_ind [1]);
	assign _4158_ = \mchip.pong.game.vga.pix_ind [3] | \mchip.pong.game.vga.pix_ind [2];
	assign _4159_ = _4158_ | ~_4157_;
	assign _4160_ = _4156_ & ~_4159_;
	assign _4161_ = _4154_ & ~_4160_;
	assign _4162_ = \mchip.pong.game.vga.pix_ind [9] | \mchip.pong.game.vga.pix_ind [8];
	assign _4163_ = _4162_ | _4161_;
	assign _4164_ = _4160_ & ~_4162_;
	assign \mchip.pong.VGA_HS  = _4164_ | _4163_;
	assign _4165_ = ~(\mchip.pong.game.ball.cpath.state [5] | \mchip.pong.game.ball.cpath.state [7]);
	assign _4166_ = \mchip.pong.game.ball.cpath.state [3] | \mchip.pong.game.ball.cpath.state [2];
	assign _0033_ = _4165_ & ~_4166_;
	assign _4167_ = _0884_ & ~_0949_;
	assign _4168_ = _4167_ | _0840_;
	assign \mchip.pong.game.right_paddle.next_coord [3] = _4168_ ^ _0851_;
	assign _4169_ = \mchip.pong.sync.o_out [5] & \mchip.pong.game.right_paddle.coord [5];
	assign _4170_ = _1004_ & _0807_;
	assign _4171_ = _4170_ | _4169_;
	assign _4172_ = ~(_1004_ & _0818_);
	assign _4173_ = ~(_4172_ | _0971_);
	assign _4174_ = _4173_ | _4171_;
	assign _4175_ = \mchip.pong.game.right_paddle.coord [6] ^ \mchip.pong.sync.o_out [5];
	assign \mchip.pong.game.right_paddle.next_coord [6] = _4175_ ^ _4174_;
	assign _4176_ = \mchip.pong.game.right_paddle.coord [6] & \mchip.pong.sync.o_out [5];
	assign _4177_ = _4175_ & _4174_;
	assign _4178_ = _4177_ | _4176_;
	assign _4179_ = \mchip.pong.game.right_paddle.coord [7] ^ \mchip.pong.sync.o_out [5];
	assign \mchip.pong.game.right_paddle.next_coord [7] = _4179_ ^ _4178_;
	assign _4180_ = \mchip.pong.game.right_paddle.coord [7] & \mchip.pong.sync.o_out [5];
	assign _4181_ = _4179_ & _4176_;
	assign _4182_ = _4181_ | _4180_;
	assign _4183_ = ~(_4179_ & _4175_);
	assign _4184_ = _4171_ & ~_4183_;
	assign _4185_ = _4184_ | _4182_;
	assign _4186_ = _4183_ | _4172_;
	assign _4187_ = ~(_4186_ | _0971_);
	assign _4188_ = _4187_ | _4185_;
	assign _4189_ = \mchip.pong.game.right_paddle.coord [8] ^ \mchip.pong.sync.o_out [5];
	assign \mchip.pong.game.right_paddle.next_coord [8] = _4189_ ^ _4188_;
	assign _4190_ = ~(_4075_ & _1208_);
	assign _4191_ = _4190_ | _3205_;
	assign _4192_ = \mchip.pong.game.ball.cpath.state [5] & ~_4191_;
	assign _4193_ = _4113_ | _4091_;
	assign _4194_ = \mchip.pong.game.ball.cpath.state [3] & ~_4193_;
	assign _4195_ = \mchip.pong.game.ball.cpath.state [2] & ~_4119_;
	assign _4196_ = _4195_ | _4194_;
	assign _0003_ = _4196_ | _4192_;
	assign _0010_ = \mchip.pong.sync.o_out [2] | ~\mchip.pong.game.vga.pclk_ctr ;
	assign _4197_ = _4091_ | _4062_;
	assign _4198_ = \mchip.pong.game.ball.cpath.state [2] & ~_4197_;
	assign _4199_ = \mchip.pong.game.ball.cpath.state [3] & ~_3216_;
	assign _4200_ = _4190_ | _4061_;
	assign _4201_ = \mchip.pong.game.ball.cpath.state [7] & ~_4200_;
	assign _4202_ = _4201_ | _4199_;
	assign _0002_ = _4202_ | _4198_;
	assign \mchip.pong.game.right_paddle.next_coord [2] = ~(_0949_ ^ _0884_);
	assign _4203_ = ~\mchip.pong.game.vga.line_ind [2];
	assign _4204_ = _1045_ & ~_4203_;
	assign _4205_ = ~(_4204_ ^ \mchip.pong.game.vga.line_ind [3]);
	assign _4206_ = _1045_ ^ _4203_;
	assign _4207_ = _4206_ | _4205_;
	assign _4208_ = _1144_ & ~_4207_;
	assign _4209_ = ~\mchip.pong.game.vga.line_ind [5];
	assign _4210_ = \mchip.pong.game.vga.line_ind [4] & ~\mchip.pong.game.vga.line_ind [5];
	assign _4211_ = ~(\mchip.pong.game.vga.line_ind [2] & \mchip.pong.game.vga.line_ind [3]);
	assign _4212_ = _1045_ & ~_4211_;
	assign _4213_ = _4212_ & _4210_;
	assign _4214_ = _4209_ & ~_4213_;
	assign _4215_ = _4214_ & ~\mchip.pong.game.vga.line_ind [6];
	assign _4216_ = _4215_ ^ \mchip.pong.game.vga.line_ind [7];
	assign _4217_ = _4214_ ^ \mchip.pong.game.vga.line_ind [6];
	assign _4218_ = ~(_4217_ & _4216_);
	assign _4219_ = _4212_ & \mchip.pong.game.vga.line_ind [4];
	assign _4220_ = _4219_ ^ _4209_;
	assign _4221_ = _4212_ ^ \mchip.pong.game.vga.line_ind [4];
	assign _4222_ = ~_4221_;
	assign _4223_ = _4222_ | _4220_;
	assign _4224_ = _4223_ | _4218_;
	assign _4225_ = _4224_ | ~_4208_;
	assign _4226_ = _4209_ & ~_1089_;
	assign _4227_ = _1089_ | ~_4210_;
	assign _4228_ = _4212_ & ~_4227_;
	assign _4229_ = _4226_ & ~_4228_;
	assign _4230_ = _4229_ ^ \mchip.pong.game.vga.line_ind [8];
	assign _4231_ = _4230_ & ~_4225_;
	assign _4232_ = ~(\mchip.pong.game.vga.pix_ind [6] & \mchip.pong.game.vga.pix_ind [7]);
	assign _4233_ = \mchip.pong.game.vga.pix_ind [7] & ~\mchip.pong.game.vga.pix_ind [6];
	assign _4234_ = ~(\mchip.pong.game.vga.pix_ind [4] | \mchip.pong.game.vga.pix_ind [5]);
	assign _4235_ = _4233_ & ~_4234_;
	assign _4236_ = _4232_ & ~_4235_;
	assign _4237_ = _4236_ ^ \mchip.pong.game.vga.pix_ind [8];
	assign _4238_ = _4236_ & ~\mchip.pong.game.vga.pix_ind [8];
	assign _4239_ = _4238_ ^ \mchip.pong.game.vga.pix_ind [9];
	assign _4240_ = _4239_ & ~_4237_;
	assign _4241_ = ~\mchip.pong.game.vga.pix_ind [7];
	assign _4242_ = _4234_ & ~\mchip.pong.game.vga.pix_ind [6];
	assign _4243_ = _4242_ ^ _4241_;
	assign _4244_ = _4234_ ^ \mchip.pong.game.vga.pix_ind [6];
	assign _4245_ = _4244_ & ~_4243_;
	assign _4246_ = ~(_4245_ & _4234_);
	assign _4247_ = _4103_ & ~_4246_;
	assign _4248_ = ~(_4247_ & _4240_);
	assign _4249_ = _4231_ & ~_4248_;
	assign _4250_ = ~(\mchip.pong.game.vga.line_ind [6] & \mchip.pong.game.vga.line_ind [7]);
	assign _4251_ = ~(\mchip.pong.game.vga.line_ind [4] & \mchip.pong.game.vga.line_ind [5]);
	assign _4252_ = _4251_ | _4250_;
	assign _4253_ = _4212_ & ~_4252_;
	assign _4254_ = \mchip.pong.game.vga.line_ind [9] | ~\mchip.pong.game.vga.line_ind [8];
	assign _4255_ = _4253_ & ~_4254_;
	assign _4256_ = _4255_ | \mchip.pong.game.vga.line_ind [9];
	assign _4257_ = ~(_4228_ & _1122_);
	assign _4258_ = \mchip.pong.game.vga.line_ind [5] | \mchip.pong.game.vga.line_ind [6];
	assign _4259_ = \mchip.pong.game.vga.line_ind [8] | \mchip.pong.game.vga.line_ind [7];
	assign _4260_ = _4259_ | _4258_;
	assign _4261_ = _4260_ | \mchip.pong.game.vga.line_ind [9];
	assign _4262_ = _4257_ & ~_4261_;
	assign _4263_ = _4262_ | _4256_;
	assign _4264_ = _4234_ & _4098_;
	assign _4265_ = _4097_ & ~_4264_;
	assign _4266_ = ~(_4233_ & _4099_);
	assign _4267_ = _4266_ | _4159_;
	assign _4268_ = _4267_ | _4162_;
	assign _4269_ = _4234_ & _4233_;
	assign _4270_ = _4269_ | _4241_;
	assign _4271_ = _4267_ & ~_4270_;
	assign _4272_ = _4271_ | _4162_;
	assign _4273_ = _4268_ & ~_4272_;
	assign _4274_ = _4273_ | _4265_;
	assign _4275_ = _4274_ | _4263_;
	assign _4276_ = _4249_ & ~_4275_;
	assign _4277_ = ~(\mchip.pong.sync.o_out [4] | \mchip.pong.sync.o_out [5]);
	assign _4278_ = _4276_ & ~_4277_;
	assign _4279_ = \mchip.pong.game.right_paddle.next_coord [8] & \mchip.pong.game.right_paddle.next_coord [7];
	assign _4280_ = ~(\mchip.pong.game.right_paddle.next_coord [6] & \mchip.pong.game.right_paddle.next_coord [5]);
	assign _4281_ = \mchip.pong.game.right_paddle.next_coord [6] & ~\mchip.pong.game.right_paddle.next_coord [5];
	assign _4282_ = ~(\mchip.pong.game.right_paddle.next_coord [3] | \mchip.pong.game.right_paddle.next_coord [4]);
	assign _4283_ = _4281_ & ~_4282_;
	assign _4284_ = _4280_ & ~_4283_;
	assign _4285_ = _4279_ & ~_4284_;
	assign _4286_ = ~(\mchip.pong.game.right_paddle.next_coord [7] & \mchip.pong.game.right_paddle.next_coord [6]);
	assign _4287_ = \mchip.pong.game.right_paddle.next_coord [4] | \mchip.pong.game.right_paddle.next_coord [5];
	assign _4288_ = _4287_ | _4286_;
	assign _4289_ = \mchip.pong.game.right_paddle.next_coord [3] & ~\mchip.pong.game.right_paddle.next_coord [2];
	assign _4290_ = ~(_4289_ & _0938_);
	assign _4291_ = _4290_ | _4288_;
	assign _4292_ = \mchip.pong.game.right_paddle.next_coord [8] & ~_4291_;
	assign _4293_ = _4285_ & ~_4292_;
	assign _0012_ = _4278_ & ~_4293_;
	assign \mchip.pong.game.left_paddle.next_coord [2] = ~(_0699_ ^ _0644_);
	assign _4294_ = ~(\mchip.pong.sync.o_out [6] | \mchip.pong.sync.o_out [7]);
	assign _4295_ = _4276_ & ~_4294_;
	assign _4296_ = ~(\mchip.pong.game.left_paddle.next_coord [7] & \mchip.pong.game.left_paddle.next_coord [6]);
	assign _4297_ = \mchip.pong.game.left_paddle.next_coord [5] | \mchip.pong.game.left_paddle.next_coord [4];
	assign _4298_ = _4297_ | _4296_;
	assign _4299_ = \mchip.pong.game.left_paddle.next_coord [3] & ~\mchip.pong.game.left_paddle.next_coord [2];
	assign _4300_ = ~(_4299_ & _0688_);
	assign _4301_ = ~(_4300_ | _4298_);
	assign _4302_ = ~(_4301_ & \mchip.pong.game.left_paddle.next_coord [8]);
	assign _4303_ = ~(\mchip.pong.game.left_paddle.next_coord [6] & \mchip.pong.game.left_paddle.next_coord [5]);
	assign _4304_ = \mchip.pong.game.left_paddle.next_coord [6] & ~\mchip.pong.game.left_paddle.next_coord [5];
	assign _4305_ = ~(\mchip.pong.game.left_paddle.next_coord [3] | \mchip.pong.game.left_paddle.next_coord [4]);
	assign _4306_ = _4304_ & ~_4305_;
	assign _4307_ = _4303_ & ~_4306_;
	assign _4308_ = ~(\mchip.pong.game.left_paddle.next_coord [8] & \mchip.pong.game.left_paddle.next_coord [7]);
	assign _4309_ = _4308_ | _4307_;
	assign _4310_ = _4302_ & ~_4309_;
	assign _0011_ = _4295_ & ~_4310_;
	assign \mchip.pong.game.ball.dpath.en_pos_reg  = _4276_ | _0033_;
	assign _4311_ = \mchip.pong.game.vga.line_ind [2] | ~\mchip.pong.game.vga.line_ind [3];
	assign _4312_ = \mchip.pong.game.vga.line_ind [0] | \mchip.pong.game.vga.line_ind [1];
	assign _4313_ = _4312_ | _4311_;
	assign _4314_ = ~(_4313_ | _1100_);
	assign _4315_ = \mchip.pong.game.vga.line_ind [8] | ~\mchip.pong.game.vga.line_ind [9];
	assign _4316_ = _4314_ & ~_4315_;
	assign _0013_ = ~(_4316_ | \mchip.pong.game.vga.line_ind [0]);
	assign _4317_ = \mchip.pong.game.vga.line_ind [0] ^ \mchip.pong.game.vga.line_ind [1];
	assign _0014_ = _4317_ & ~_4316_;
	assign _4318_ = _1045_ ^ \mchip.pong.game.vga.line_ind [2];
	assign _0015_ = _4318_ & ~_4316_;
	assign _4319_ = _4204_ ^ \mchip.pong.game.vga.line_ind [3];
	assign _0016_ = _4319_ & ~_4316_;
	assign _0017_ = _4221_ & ~_4316_;
	assign _0018_ = ~(_4316_ | _4220_);
	assign _4320_ = _4212_ & ~_4251_;
	assign _4321_ = _4320_ ^ \mchip.pong.game.vga.line_ind [6];
	assign _0019_ = _4321_ & ~_4316_;
	assign _4322_ = ~_4316_;
	assign _4323_ = ~(_4320_ & \mchip.pong.game.vga.line_ind [6]);
	assign _4324_ = _4323_ ^ \mchip.pong.game.vga.line_ind [7];
	assign _0020_ = _4322_ & ~_4324_;
	assign _4325_ = ~(_4253_ ^ \mchip.pong.game.vga.line_ind [8]);
	assign _0021_ = ~(_4325_ | _4316_);
	assign _4326_ = ~(_4253_ & \mchip.pong.game.vga.line_ind [8]);
	assign _4327_ = _4326_ ^ \mchip.pong.game.vga.line_ind [9];
	assign _0022_ = _4322_ & ~_4327_;
	assign _0023_ = _4105_ & ~\mchip.pong.game.vga.pix_ind [0];
	assign _0024_ = \mchip.pong.game.vga.pix_ind [0] ^ \mchip.pong.game.vga.pix_ind [1];
	assign _4328_ = ~\mchip.pong.game.vga.pix_ind [2];
	assign _4329_ = _4102_ ^ _4328_;
	assign _0025_ = _4105_ & ~_4329_;
	assign _4330_ = ~\mchip.pong.game.vga.pix_ind [3];
	assign _4331_ = _4102_ & ~_4328_;
	assign _4332_ = _4331_ ^ _4330_;
	assign _0026_ = _4105_ & ~_4332_;
	assign _4333_ = ~\mchip.pong.game.vga.pix_ind [4];
	assign _4334_ = _4103_ ^ _4333_;
	assign _0027_ = _4105_ & ~_4334_;
	assign _4335_ = _4103_ & ~_4333_;
	assign _4336_ = _4335_ ^ _4151_;
	assign _0028_ = _4105_ & ~_4336_;
	assign _4337_ = ~\mchip.pong.game.vga.pix_ind [6];
	assign _4338_ = ~(\mchip.pong.game.vga.pix_ind [4] & \mchip.pong.game.vga.pix_ind [5]);
	assign _4339_ = _4103_ & ~_4338_;
	assign _4340_ = _4339_ ^ _4337_;
	assign _0029_ = _4105_ & ~_4340_;
	assign _4341_ = _4339_ & ~_4337_;
	assign _4342_ = _4341_ ^ _4241_;
	assign _0030_ = _4105_ & ~_4342_;
	assign _4343_ = _4338_ | _4232_;
	assign _4344_ = _4103_ & ~_4343_;
	assign _4345_ = ~(_4344_ ^ \mchip.pong.game.vga.pix_ind [8]);
	assign _0031_ = _4105_ & ~_4345_;
	assign _4346_ = ~(_4344_ & \mchip.pong.game.vga.pix_ind [8]);
	assign _4347_ = _4346_ ^ \mchip.pong.game.vga.pix_ind [9];
	assign _0032_ = _4105_ & ~_4347_;
	assign _4348_ = ~(\mchip.pong.game.vga.pix_ind [4] | \mchip.pong.game.ball.dpath.ballX [4]);
	assign _4349_ = \mchip.pong.game.vga.pix_ind [3] & ~\mchip.pong.game.ball.dpath.ballX [3];
	assign _4350_ = \mchip.pong.game.vga.pix_ind [2] & ~\mchip.pong.game.ball.dpath.ballX [2];
	assign _4351_ = \mchip.pong.game.vga.pix_ind [3] | ~\mchip.pong.game.ball.dpath.ballX [3];
	assign _4352_ = _4351_ & ~_4349_;
	assign _4353_ = _4352_ & _4350_;
	assign _4354_ = _4353_ | _4349_;
	assign _4355_ = \mchip.pong.game.ball.dpath.ballX [1] & ~\mchip.pong.game.vga.pix_ind [1];
	assign _4356_ = \mchip.pong.game.ball.dpath.ballX [2] & ~\mchip.pong.game.vga.pix_ind [2];
	assign _4357_ = ~(_4350_ | _4356_);
	assign _4358_ = _4352_ & _4357_;
	assign _4359_ = _4358_ & ~_4355_;
	assign _4360_ = _4359_ | _4354_;
	assign _4361_ = \mchip.pong.game.vga.pix_ind [4] & \mchip.pong.game.ball.dpath.ballX [4];
	assign _4362_ = ~(_4361_ | _4348_);
	assign _4363_ = _4362_ & _4360_;
	assign _4364_ = _4363_ | _4348_;
	assign _4365_ = _4338_ & ~_4234_;
	assign _4366_ = _4365_ ^ \mchip.pong.game.ball.dpath.ballX [5];
	assign _4367_ = _4366_ ^ _4364_;
	assign _4368_ = _4362_ ^ _4360_;
	assign _4369_ = ~(\mchip.pong.game.ball.dpath.ballY [0] & \mchip.pong.game.vga.line_ind [0]);
	assign _4370_ = _4317_ ^ \mchip.pong.game.ball.dpath.ballY [1];
	assign _4371_ = ~(_4370_ ^ _4369_);
	assign _4372_ = ~_4371_;
	assign _4373_ = \mchip.pong.game.ball.dpath.ballY [0] | \mchip.pong.game.vga.line_ind [0];
	assign _4374_ = ~(_4369_ & _4373_);
	assign _4375_ = _4371_ & _4374_;
	assign _4376_ = ~(_4317_ & _3073_);
	assign _4377_ = _4369_ & ~_4370_;
	assign _4378_ = _4376_ & ~_4377_;
	assign _4379_ = _4318_ ^ \mchip.pong.game.ball.dpath.ballY [2];
	assign _4380_ = _4379_ ^ _4378_;
	assign _4381_ = (_4380_ ? _4372_ : _4375_);
	assign _4382_ = _4379_ | _4378_;
	assign _4383_ = _3029_ & ~_4206_;
	assign _4384_ = _4383_ | ~_4382_;
	assign _4385_ = _4319_ ^ \mchip.pong.game.ball.dpath.ballY [3];
	assign _4386_ = ~_4385_;
	assign _4387_ = _4386_ ^ _4384_;
	assign _4388_ = _4377_ | ~_4376_;
	assign _4389_ = _4379_ ^ _4388_;
	assign _4390_ = _4374_ & ~_4389_;
	assign _4391_ = ~_4390_;
	assign _4392_ = (_4387_ ? _4391_ : _4381_);
	assign _4393_ = ~\mchip.pong.game.ball.dpath.ballY [3];
	assign _4394_ = _4393_ & ~_4205_;
	assign _4395_ = _4383_ & ~_4385_;
	assign _4396_ = _4395_ | _4394_;
	assign _4397_ = _4385_ | _4379_;
	assign _4398_ = _4388_ & ~_4397_;
	assign _4399_ = _4398_ | _4396_;
	assign _4400_ = ~(_4221_ & _2625_);
	assign _4401_ = \mchip.pong.game.ball.dpath.ballY [4] & ~_4221_;
	assign _4402_ = _4400_ & ~_4401_;
	assign _0127_ = _4402_ ^ _4399_;
	assign _4403_ = _4392_ & ~_0127_;
	assign _4404_ = _4402_ & _4399_;
	assign _4405_ = _4404_ | ~_4400_;
	assign _4406_ = _4220_ ^ _2658_;
	assign _0146_ = _4406_ ^ _4405_;
	assign _4407_ = ~(_4371_ | _4374_);
	assign _4408_ = ~_4407_;
	assign _4409_ = _4408_ & _4389_;
	assign _4410_ = ~_4409_;
	assign _4411_ = _4382_ & ~_4383_;
	assign _4412_ = _4385_ ^ _4411_;
	assign _4413_ = _4389_ & ~_4374_;
	assign _4414_ = (_4412_ ? _4410_ : _4413_);
	assign _4415_ = _0127_ & ~_4414_;
	assign _4416_ = (_0146_ ? _4403_ : _4415_);
	assign _4417_ = _4389_ & ~_4408_;
	assign _4418_ = _4417_ & ~_4387_;
	assign _4419_ = _4371_ & ~_4374_;
	assign _4420_ = (_4389_ ? _4419_ : _4375_);
	assign _4421_ = _4387_ & ~_4420_;
	assign _4422_ = (_0127_ ? _4418_ : _4421_);
	assign _4423_ = _4385_ ^ _4384_;
	assign _4424_ = _4374_ & ~_4371_;
	assign _4425_ = (_4389_ ? _4407_ : _4424_);
	assign _4426_ = _4423_ & ~_4425_;
	assign _4427_ = ~_4375_;
	assign _4428_ = ~(_4389_ | _4427_);
	assign _4429_ = _4428_ & ~_4423_;
	assign _4430_ = (_0127_ ? _4426_ : _4429_);
	assign _4431_ = (_0146_ ? _4422_ : _4430_);
	assign _4432_ = (\mchip.pong.game.vga.pix_ind [0] ? _4416_ : _4431_);
	assign _1103_ = ~(\mchip.pong.game.vga.pix_ind [1] ^ \mchip.pong.game.ball.dpath.ballX [1]);
	assign _4433_ = ~(_4424_ | _4419_);
	assign _4434_ = _4389_ & ~_4433_;
	assign _4435_ = _4387_ & ~_4434_;
	assign _4436_ = _4435_ | _0127_;
	assign _0056_ = ~(_4402_ ^ _4399_);
	assign _4437_ = _4424_ & ~_4389_;
	assign _4438_ = _4423_ & ~_4437_;
	assign _4439_ = _4438_ | _0056_;
	assign _4440_ = (_0146_ ? _4436_ : _4439_);
	assign _4441_ = \mchip.pong.game.vga.pix_ind [0] & ~_4440_;
	assign _4442_ = ~\mchip.pong.game.vga.pix_ind [0];
	assign _4443_ = _4389_ & _4427_;
	assign _4444_ = (_4389_ ? _4375_ : _4408_);
	assign _4445_ = (_4387_ ? _4444_ : _4443_);
	assign _0034_ = _4445_ | _0127_;
	assign _0035_ = _4408_ & ~_4389_;
	assign _0036_ = (_4380_ ? _4407_ : _4427_);
	assign _0037_ = (_4423_ ? _0036_ : _0035_);
	assign _0038_ = _0037_ | _0056_;
	assign _0039_ = (_0146_ ? _0034_ : _0038_);
	assign _0040_ = _4442_ & ~_0039_;
	assign _0041_ = _0040_ | _4441_;
	assign _0042_ = (_1103_ ? _4432_ : _0041_);
	assign _0043_ = ~_4355_;
	assign _0044_ = _4357_ ^ _0043_;
	assign _0045_ = (_4380_ ? _4371_ : _4424_);
	assign _0046_ = _0045_ | _4387_;
	assign _0047_ = _0046_ | _0056_;
	assign _0048_ = _4381_ & ~_4423_;
	assign _0049_ = ~(_0048_ & _0056_);
	assign _0050_ = (_0146_ ? _0047_ : _0049_);
	assign _0051_ = _0035_ | ~_4423_;
	assign _0052_ = ~(_4428_ & _4387_);
	assign _0053_ = (_0127_ ? _0051_ : _0052_);
	assign _0054_ = _4427_ & ~_4389_;
	assign _0055_ = ~(_0054_ & _4387_);
	assign _0057_ = _4417_ & _4423_;
	assign _0058_ = ~_0057_;
	assign _0059_ = (_0056_ ? _0055_ : _0058_);
	assign _0060_ = (_0146_ ? _0053_ : _0059_);
	assign _0061_ = (\mchip.pong.game.vga.pix_ind [0] ? _0060_ : _0050_);
	assign _0062_ = _1103_ & ~_0061_;
	assign _0063_ = ~_1103_;
	assign _0064_ = _4391_ | ~_4387_;
	assign _0065_ = ~_4419_;
	assign _0066_ = _0065_ & _4389_;
	assign _0067_ = ~_0066_;
	assign _0068_ = _0067_ | _4387_;
	assign _0069_ = (_0056_ ? _0064_ : _0068_);
	assign _0070_ = ~_4413_;
	assign _0071_ = _0070_ | _4412_;
	assign _0072_ = _4389_ | ~_4387_;
	assign _0073_ = (_0127_ ? _0071_ : _0072_);
	assign _0074_ = (_0146_ ? _0069_ : _0073_);
	assign _0075_ = _4387_ | ~_4417_;
	assign _0076_ = _0036_ | ~_4387_;
	assign _0077_ = (_0127_ ? _0075_ : _0076_);
	assign _0078_ = _4444_ | ~_4423_;
	assign _0079_ = (_0056_ ? _0064_ : _0078_);
	assign _0080_ = (_0146_ ? _0077_ : _0079_);
	assign _0081_ = (\mchip.pong.game.vga.pix_ind [0] ? _0080_ : _0074_);
	assign _0082_ = _0063_ & ~_0081_;
	assign _0083_ = _0082_ | _0062_;
	assign _0084_ = (_0044_ ? _0042_ : _0083_);
	assign _0085_ = _4357_ & ~_4355_;
	assign _0086_ = ~(_0085_ | _4350_);
	assign _0087_ = ~_4352_;
	assign _0088_ = _0087_ ^ _0086_;
	assign _0089_ = _4427_ & ~_4380_;
	assign _0090_ = ~_0089_;
	assign _0091_ = ~(_4423_ & _0090_);
	assign _0092_ = _0127_ & ~_0091_;
	assign _0093_ = _4408_ | _4389_;
	assign _0094_ = _0093_ & ~_4409_;
	assign _0095_ = _0094_ | _4423_;
	assign _0096_ = _0056_ & ~_0095_;
	assign _0097_ = (_0146_ ? _0092_ : _0096_);
	assign _0098_ = ~(_4423_ & _4381_);
	assign _0099_ = _0127_ & ~_0098_;
	assign _0100_ = _4389_ & _4371_;
	assign _0101_ = _4389_ | _4371_;
	assign _0102_ = _0101_ & ~_0100_;
	assign _0103_ = _0102_ | _4423_;
	assign _0104_ = _0056_ & ~_0103_;
	assign _0105_ = (_0146_ ? _0099_ : _0104_);
	assign _0106_ = (\mchip.pong.game.vga.pix_ind [0] ? _0105_ : _0097_);
	assign _0107_ = ~_4417_;
	assign _0108_ = (_4423_ ? _4389_ : _0107_);
	assign _0109_ = _0127_ & ~_0108_;
	assign _0110_ = ~(_4389_ & _4387_);
	assign _0111_ = _0056_ & ~_0110_;
	assign _0112_ = (_0146_ ? _0109_ : _0111_);
	assign _0113_ = ~_4443_;
	assign _0114_ = _4389_ | ~_4371_;
	assign _0115_ = (_4387_ ? _0113_ : _0114_);
	assign _0116_ = _0056_ & ~_0115_;
	assign _0117_ = ~_0035_;
	assign _0118_ = _4389_ & ~_4371_;
	assign _0119_ = ~_0118_;
	assign _0120_ = (_4387_ ? _0119_ : _0117_);
	assign _0121_ = _0127_ & ~_0120_;
	assign _0122_ = (_0146_ ? _0121_ : _0116_);
	assign _0123_ = (\mchip.pong.game.vga.pix_ind [0] ? _0112_ : _0122_);
	assign _0124_ = (_1103_ ? _0123_ : _0106_);
	assign _0125_ = ~(_0035_ & _4423_);
	assign _0126_ = _0056_ & ~_0125_;
	assign _0128_ = ~(_4443_ & _4387_);
	assign _0129_ = _0127_ & ~_0128_;
	assign _0130_ = (_0146_ ? _0129_ : _0126_);
	assign _0131_ = ~_4428_;
	assign _0132_ = (_4387_ ? _4380_ : _0131_);
	assign _0133_ = _0127_ & ~_0132_;
	assign _0134_ = ~(_0054_ & _4423_);
	assign _0135_ = _0056_ & ~_0134_;
	assign _0136_ = (_0146_ ? _0133_ : _0135_);
	assign _0137_ = (\mchip.pong.game.vga.pix_ind [0] ? _0136_ : _0130_);
	assign _0138_ = _0119_ | ~_4387_;
	assign _0139_ = _0127_ & ~_0138_;
	assign _0140_ = _0114_ | ~_4423_;
	assign _0141_ = ~(_0140_ | _0127_);
	assign _0142_ = (_0146_ ? _0139_ : _0141_);
	assign _0143_ = (_4387_ ? _0107_ : _0131_);
	assign _0144_ = _0127_ & ~_0143_;
	assign _0145_ = _0056_ & ~_0120_;
	assign _0147_ = (_0146_ ? _0144_ : _0145_);
	assign _0148_ = (\mchip.pong.game.vga.pix_ind [0] ? _0147_ : _0142_);
	assign _0149_ = (_1103_ ? _0137_ : _0148_);
	assign _0150_ = (_0044_ ? _0124_ : _0149_);
	assign _0151_ = (_0088_ ? _0084_ : _0150_);
	assign _0152_ = ~_0088_;
	assign _0153_ = (_4389_ ? _4371_ : _4407_);
	assign _0154_ = _0153_ & ~_4423_;
	assign _0155_ = _0154_ & ~_0056_;
	assign _0156_ = _0056_ & ~_0098_;
	assign _0157_ = (_0146_ ? _0155_ : _0156_);
	assign _0158_ = _4400_ & ~_4404_;
	assign _0159_ = _4406_ ^ _0158_;
	assign _0160_ = _0153_ & ~_4387_;
	assign _0161_ = _0160_ & ~_0127_;
	assign _0162_ = ~(_4387_ & _4381_);
	assign _0163_ = _0127_ & ~_0162_;
	assign _0164_ = (_0159_ ? _0161_ : _0163_);
	assign _0165_ = (\mchip.pong.game.vga.pix_ind [0] ? _0164_ : _0157_);
	assign _0166_ = ~(_4409_ & _4387_);
	assign _0167_ = _0127_ & ~_0166_;
	assign _0168_ = (_0146_ ? _0167_ : _0135_);
	assign _0169_ = (\mchip.pong.game.vga.pix_ind [0] ? _0157_ : _0168_);
	assign _0170_ = (_1103_ ? _0165_ : _0169_);
	assign _0171_ = _4423_ | ~_4437_;
	assign _0172_ = _0127_ & ~_0171_;
	assign _0173_ = ~(_4443_ & _4423_);
	assign _0174_ = _0056_ & ~_0173_;
	assign _0175_ = (_0146_ ? _0172_ : _0174_);
	assign _0176_ = (\mchip.pong.game.vga.pix_ind [0] ? _0164_ : _0175_);
	assign _0177_ = _0127_ & ~_0055_;
	assign _0178_ = (_0159_ ? _0161_ : _0177_);
	assign _0179_ = ~(_0101_ | _4423_);
	assign _0180_ = _0179_ & ~_0056_;
	assign _0181_ = ~(_4423_ & _4409_);
	assign _0182_ = _0056_ & ~_0181_;
	assign _0183_ = (_0146_ ? _0180_ : _0182_);
	assign _0184_ = (\mchip.pong.game.vga.pix_ind [0] ? _0183_ : _0178_);
	assign _0185_ = (_1103_ ? _0176_ : _0184_);
	assign _0186_ = (_0044_ ? _0170_ : _0185_);
	assign _0187_ = _0186_ & ~_0152_;
	assign _0188_ = _0055_ | _0056_;
	assign _0189_ = ~(_4434_ & _4423_);
	assign _0190_ = _0189_ | _0127_;
	assign _0191_ = (_0146_ ? _0188_ : _0190_);
	assign _0192_ = _0181_ | _0127_;
	assign _0193_ = _4423_ | _4389_;
	assign _0194_ = _0193_ | _0056_;
	assign _0195_ = (_0146_ ? _0194_ : _0192_);
	assign _0196_ = (\mchip.pong.game.vga.pix_ind [0] ? _0195_ : _0191_);
	assign _0197_ = ~(_4423_ & _4389_);
	assign _0198_ = _0197_ | _0127_;
	assign _0199_ = ~(_0035_ & _4387_);
	assign _0200_ = _0199_ | _0056_;
	assign _0201_ = (_0159_ ? _0198_ : _0200_);
	assign _0202_ = (_1103_ ? _0196_ : _0201_);
	assign _0203_ = ~(_0065_ | _4389_);
	assign _0204_ = ~(_0203_ & _4387_);
	assign _0205_ = _0204_ | _0056_;
	assign _0206_ = _4424_ & _4389_;
	assign _0207_ = ~_0206_;
	assign _0208_ = ~(_0207_ | _4387_);
	assign _0209_ = _0208_ & ~_0127_;
	assign _0210_ = ~_0209_;
	assign _0211_ = (_0146_ ? _0205_ : _0210_);
	assign _0212_ = (_0146_ ? _0188_ : _0210_);
	assign _0213_ = (_1103_ ? _0211_ : _0212_);
	assign _0214_ = (_0044_ ? _0202_ : _0213_);
	assign _0215_ = _0152_ & ~_0214_;
	assign _0216_ = _0215_ | _0187_;
	assign _0217_ = (_4368_ ? _0151_ : _0216_);
	assign _0218_ = (_0146_ ? _0188_ : _0192_);
	assign _0219_ = (\mchip.pong.game.vga.pix_ind [0] ? _0218_ : _0195_);
	assign _0220_ = (_1103_ ? _0219_ : _0212_);
	assign _0221_ = _0044_ & ~_0220_;
	assign _0222_ = ~(_0189_ | _0127_);
	assign _0223_ = (_0146_ ? _0172_ : _0222_);
	assign _0224_ = (\mchip.pong.game.vga.pix_ind [0] ? _0223_ : _0164_);
	assign _0225_ = _0056_ & ~_0197_;
	assign _0226_ = _0127_ & ~_0199_;
	assign _0227_ = (_0159_ ? _0225_ : _0226_);
	assign _0228_ = (_0146_ ? _0226_ : _0174_);
	assign _0229_ = (\mchip.pong.game.vga.pix_ind [0] ? _0227_ : _0228_);
	assign _0230_ = (_1103_ ? _0224_ : _0229_);
	assign _0231_ = _0230_ & ~_0044_;
	assign _0232_ = _0231_ | _0221_;
	assign _0233_ = (\mchip.pong.game.vga.pix_ind [0] ? _0157_ : _0164_);
	assign _0234_ = _0093_ | _4423_;
	assign _0235_ = _0127_ & ~_0234_;
	assign _0236_ = (_0146_ ? _0235_ : _0182_);
	assign _0237_ = _0094_ | _4387_;
	assign _0238_ = _0056_ & ~_0237_;
	assign _0239_ = (_0146_ ? _0177_ : _0238_);
	assign _0240_ = (\mchip.pong.game.vga.pix_ind [0] ? _0239_ : _0236_);
	assign _0241_ = (_1103_ ? _0233_ : _0240_);
	assign _0242_ = _0056_ & ~_0108_;
	assign _0243_ = (_0146_ ? _0133_ : _0242_);
	assign _0244_ = ~(_4434_ & _4387_);
	assign _0245_ = _0127_ & ~_0244_;
	assign _0246_ = (_0146_ ? _0245_ : _0126_);
	assign _0247_ = (\mchip.pong.game.vga.pix_ind [0] ? _0246_ : _0243_);
	assign _0248_ = (\mchip.pong.game.vga.pix_ind [0] ? _0168_ : _0157_);
	assign _0249_ = (_1103_ ? _0247_ : _0248_);
	assign _0250_ = (_0044_ ? _0241_ : _0249_);
	assign _0251_ = (_0088_ ? _0232_ : _0250_);
	assign _0252_ = (_4423_ ? _0094_ : _4390_);
	assign _0253_ = _0056_ & ~_0252_;
	assign _0254_ = _4427_ | ~_4389_;
	assign _0255_ = _0254_ & ~_0054_;
	assign _0256_ = (_4423_ ? _4413_ : _0255_);
	assign _0257_ = _0127_ & ~_0256_;
	assign _0258_ = (_0146_ ? _0253_ : _0257_);
	assign _0259_ = ~(_4407_ | _4375_);
	assign _0260_ = (_4389_ ? _0259_ : _4375_);
	assign _0261_ = _4387_ & ~_0260_;
	assign _0262_ = (_0127_ ? _4418_ : _0261_);
	assign _0263_ = (_4389_ ? _4407_ : _0259_);
	assign _0264_ = ~_0263_;
	assign _0265_ = _0264_ & _4423_;
	assign _0266_ = (_0056_ ? _4429_ : _0265_);
	assign _0267_ = (_0146_ ? _0262_ : _0266_);
	assign _0268_ = (\mchip.pong.game.vga.pix_ind [0] ? _0267_ : _0258_);
	assign _0269_ = _4387_ & ~_0036_;
	assign _0270_ = ~(_0119_ | _4387_);
	assign _0271_ = (_0056_ ? _0269_ : _0270_);
	assign _0272_ = _4423_ & ~_4444_;
	assign _0273_ = (_0056_ ? _4429_ : _0272_);
	assign _0274_ = (_0146_ ? _0271_ : _0273_);
	assign _0275_ = _4387_ & ~_4391_;
	assign _0276_ = _4386_ ^ _4411_;
	assign _0277_ = _0276_ & ~_0067_;
	assign _0278_ = (_0056_ ? _0275_ : _0277_);
	assign _0279_ = _4423_ & ~_0070_;
	assign _0280_ = ~(_4424_ | _4389_);
	assign _0281_ = ~_0280_;
	assign _0282_ = _4387_ & ~_0281_;
	assign _0283_ = (_0127_ ? _0279_ : _0282_);
	assign _0284_ = (_0146_ ? _0278_ : _0283_);
	assign _0285_ = (\mchip.pong.game.vga.pix_ind [0] ? _0284_ : _0274_);
	assign _0286_ = (_1103_ ? _0268_ : _0285_);
	assign _0287_ = _0134_ | _0127_;
	assign _0288_ = _4423_ | ~_4409_;
	assign _0289_ = _0288_ | _0056_;
	assign _0290_ = (_0146_ ? _0287_ : _0289_);
	assign _0291_ = \mchip.pong.game.vga.pix_ind [0] & ~_0290_;
	assign _0292_ = _4380_ & ~_4427_;
	assign _0293_ = (_4423_ ? _0292_ : _0207_);
	assign _0294_ = _0056_ & ~_0293_;
	assign _0295_ = ~_0203_;
	assign _0296_ = (_4423_ ? _0295_ : _4417_);
	assign _0297_ = _0127_ & ~_0296_;
	assign _0298_ = (_0146_ ? _0294_ : _0297_);
	assign _0299_ = (_4389_ ? _4371_ : _4408_);
	assign _0300_ = (_4423_ ? _4417_ : _0299_);
	assign _0301_ = _0056_ & ~_0300_;
	assign _0302_ = (_4387_ ? _0292_ : _0036_);
	assign _0303_ = _0127_ & ~_0302_;
	assign _0304_ = (_0146_ ? _0301_ : _0303_);
	assign _0305_ = (\mchip.pong.game.vga.pix_ind [0] ? _0304_ : _0298_);
	assign _0306_ = (_1103_ ? _0291_ : _0305_);
	assign _0307_ = (_0044_ ? _0286_ : _0306_);
	assign _0308_ = ~_0044_;
	assign _0309_ = _0127_ & ~_0051_;
	assign _0310_ = _0090_ & ~_4423_;
	assign _0311_ = (_0127_ ? _4418_ : _0310_);
	assign _0312_ = (_0146_ ? _0309_ : _0311_);
	assign _0313_ = _0127_ & ~_0046_;
	assign _0314_ = (_4389_ ? _4371_ : _0065_);
	assign _0315_ = ~(_0314_ & _4387_);
	assign _0316_ = _0056_ & ~_0315_;
	assign _0317_ = (_0146_ ? _0313_ : _0316_);
	assign _0318_ = (\mchip.pong.game.vga.pix_ind [0] ? _0317_ : _0312_);
	assign _0319_ = _0154_ & ~_0127_;
	assign _0320_ = _0255_ | _4387_;
	assign _0321_ = _0127_ & ~_0320_;
	assign _0322_ = (_0159_ ? _0319_ : _0321_);
	assign _0323_ = _4389_ | _4387_;
	assign _0324_ = _0127_ & ~_0323_;
	assign _0325_ = _0035_ | ~_4387_;
	assign _0326_ = _0056_ & ~_0325_;
	assign _0327_ = (_0146_ ? _0324_ : _0326_);
	assign _0328_ = (\mchip.pong.game.vga.pix_ind [0] ? _0327_ : _0322_);
	assign _0329_ = (_1103_ ? _0318_ : _0328_);
	assign _0330_ = (_4387_ ? _0107_ : _0117_);
	assign _0331_ = _0127_ & ~_0330_;
	assign _0332_ = _0056_ & ~_0132_;
	assign _0333_ = (_0146_ ? _0331_ : _0332_);
	assign _0334_ = (_4387_ ? _0119_ : _0114_);
	assign _0335_ = _0127_ & ~_0334_;
	assign _0336_ = (_0146_ ? _0335_ : _0116_);
	assign _0337_ = (\mchip.pong.game.vga.pix_ind [0] ? _0336_ : _0333_);
	assign _0338_ = _0056_ & ~_0143_;
	assign _0339_ = (_0146_ ? _0144_ : _0338_);
	assign _0340_ = _0056_ & ~_0140_;
	assign _0341_ = (_0146_ ? _0129_ : _0340_);
	assign _0342_ = (\mchip.pong.game.vga.pix_ind [0] ? _0341_ : _0339_);
	assign _0343_ = (_1103_ ? _0337_ : _0342_);
	assign _0344_ = (_0044_ ? _0343_ : _0329_);
	assign _0345_ = (_0088_ ? _0344_ : _0307_);
	assign _0346_ = (_4368_ ? _0251_ : _0345_);
	assign _0347_ = (_4367_ ? _0217_ : _0346_);
	assign _0348_ = (_0127_ ? _0120_ : _0173_);
	assign _0349_ = ~_0348_;
	assign _0350_ = ~(_0114_ & _4423_);
	assign _0351_ = _0127_ & ~_0350_;
	assign _0352_ = _0116_ | _0351_;
	assign _0353_ = (_0146_ ? _0349_ : _0352_);
	assign _0354_ = (\mchip.pong.game.vga.pix_ind [0] ? _0112_ : _0353_);
	assign _0355_ = (_1103_ ? _0354_ : _0106_);
	assign _0356_ = ~_0128_;
	assign _0357_ = (_4387_ ? _0118_ : _0114_);
	assign _0358_ = (_0127_ ? _0356_ : _0357_);
	assign _0359_ = (_4389_ ? _4427_ : _4374_);
	assign _0360_ = (_4423_ ? _0090_ : _0359_);
	assign _0361_ = ~(_4433_ | _4389_);
	assign _0362_ = (_4423_ ? _0035_ : _0361_);
	assign _0363_ = (_0127_ ? _0360_ : _0362_);
	assign _0364_ = (_0146_ ? _0358_ : _0363_);
	assign _0365_ = ~_0132_;
	assign _0366_ = ~(_0259_ | _4389_);
	assign _0367_ = _4389_ & _4374_;
	assign _0368_ = _0367_ | _0366_;
	assign _0369_ = (_4387_ ? _4417_ : _0368_);
	assign _0370_ = (_0127_ ? _0365_ : _0369_);
	assign _0371_ = _4380_ & ~_0065_;
	assign _0372_ = ~_0371_;
	assign _0373_ = (_4423_ ? _0090_ : _0372_);
	assign _0374_ = (_4423_ ? _0054_ : _0361_);
	assign _0375_ = (_0127_ ? _0373_ : _0374_);
	assign _0376_ = (_0146_ ? _0370_ : _0375_);
	assign _0377_ = (\mchip.pong.game.vga.pix_ind [0] ? _0376_ : _0364_);
	assign _0378_ = ~_0138_;
	assign _0379_ = _0359_ & ~_4387_;
	assign _0380_ = (_0127_ ? _0378_ : _0379_);
	assign _0381_ = (_4380_ ? _4371_ : _0065_);
	assign _0382_ = (_4423_ ? _4428_ : _0381_);
	assign _0383_ = ~(_0114_ | _4387_);
	assign _0384_ = (_0127_ ? _0382_ : _0383_);
	assign _0385_ = (_0146_ ? _0380_ : _0384_);
	assign _0386_ = ~_0143_;
	assign _0387_ = _4424_ ^ _4380_;
	assign _0388_ = _4423_ & ~_0387_;
	assign _0389_ = (_0127_ ? _0386_ : _0388_);
	assign _0390_ = ~_0120_;
	assign _0391_ = ~_4381_;
	assign _0392_ = (_4423_ ? _4417_ : _0391_);
	assign _0393_ = (_0056_ ? _0390_ : _0392_);
	assign _0394_ = (_0146_ ? _0389_ : _0393_);
	assign _0395_ = (\mchip.pong.game.vga.pix_ind [0] ? _0394_ : _0385_);
	assign _0396_ = (_1103_ ? _0377_ : _0395_);
	assign _0397_ = (_0044_ ? _0355_ : _0396_);
	assign _0398_ = (_0088_ ? _0084_ : _0397_);
	assign _0399_ = ~_0166_;
	assign _0400_ = (_0127_ ? _0154_ : _0399_);
	assign _0401_ = (_4380_ ? _4371_ : _4407_);
	assign _0402_ = _0401_ | ~_4387_;
	assign _0403_ = _4389_ & ~_4424_;
	assign _0404_ = ~_0403_;
	assign _0405_ = (_4423_ ? _4381_ : _0404_);
	assign _0406_ = (_0127_ ? _0402_ : _0405_);
	assign _0407_ = (_0146_ ? _0400_ : _0406_);
	assign _0408_ = _4387_ & ~_0070_;
	assign _0409_ = (_0127_ ? _0048_ : _0408_);
	assign _0410_ = (_4389_ ? _4372_ : _4375_);
	assign _0411_ = ~(_0410_ & _4387_);
	assign _0412_ = _0065_ & ~_4389_;
	assign _0413_ = (_4423_ ? _0153_ : _0412_);
	assign _0414_ = (_0127_ ? _0411_ : _0413_);
	assign _0415_ = (_0146_ ? _0409_ : _0414_);
	assign _0416_ = (\mchip.pong.game.vga.pix_ind [0] ? _0415_ : _0407_);
	assign _0417_ = ~(_4389_ | _4374_);
	assign _0418_ = (_4423_ ? _0417_ : _4434_);
	assign _0419_ = (_0127_ ? _0399_ : _0418_);
	assign _0420_ = ~_0134_;
	assign _0421_ = ~_0292_;
	assign _0422_ = (_4387_ ? _0421_ : _4381_);
	assign _0423_ = (_0056_ ? _0420_ : _0422_);
	assign _0424_ = (_0146_ ? _0419_ : _0423_);
	assign _0425_ = ~_4424_;
	assign _0426_ = (_4389_ ? _0425_ : _0065_);
	assign _0427_ = _4423_ & ~_0426_;
	assign _0428_ = (_0127_ ? _0154_ : _0427_);
	assign _0429_ = ~_0098_;
	assign _0430_ = (_4387_ ? _0114_ : _0093_);
	assign _0431_ = (_0056_ ? _0429_ : _0430_);
	assign _0432_ = (_0146_ ? _0428_ : _0431_);
	assign _0433_ = (\mchip.pong.game.vga.pix_ind [0] ? _0432_ : _0424_);
	assign _0434_ = (_1103_ ? _0416_ : _0433_);
	assign _0435_ = _4443_ | _4428_;
	assign _0436_ = (_4423_ ? _0435_ : _4425_);
	assign _0437_ = (_4387_ ? _0372_ : _0410_);
	assign _0438_ = (_0127_ ? _0436_ : _0437_);
	assign _0439_ = (_4387_ ? _4380_ : _4443_);
	assign _0440_ = _0439_ | _0127_;
	assign _0441_ = (_0146_ ? _0438_ : _0440_);
	assign _0442_ = (_4389_ ? _4407_ : _4375_);
	assign _0443_ = (_4380_ ? _4371_ : _4419_);
	assign _0444_ = ~_0443_;
	assign _0445_ = (_4387_ ? _0444_ : _0442_);
	assign _0446_ = ~_0412_;
	assign _0447_ = _4387_ & ~_0446_;
	assign _0448_ = ~_0447_;
	assign _0449_ = (_0127_ ? _0445_ : _0448_);
	assign _0450_ = ~(_4408_ | _4380_);
	assign _0451_ = ~_0450_;
	assign _0452_ = _4423_ & ~_0451_;
	assign _0453_ = ~_0452_;
	assign _0454_ = ~_0101_;
	assign _0455_ = (_4423_ ? _0153_ : _0454_);
	assign _0456_ = (_0127_ ? _0453_ : _0455_);
	assign _0457_ = (_0146_ ? _0449_ : _0456_);
	assign _0458_ = (\mchip.pong.game.vga.pix_ind [0] ? _0457_ : _0441_);
	assign _0459_ = _0054_ & ~_4423_;
	assign _0460_ = (_4423_ ? _0421_ : _0417_);
	assign _0461_ = (_0127_ ? _0459_ : _0460_);
	assign _0462_ = (_4387_ ? _0366_ : _0153_);
	assign _0463_ = _0462_ | _0127_;
	assign _0464_ = (_0146_ ? _0461_ : _0463_);
	assign _0465_ = (_0056_ ? _0154_ : _0179_);
	assign _0466_ = (_4387_ ? _0417_ : _4409_);
	assign _0467_ = _0466_ | _0127_;
	assign _0468_ = (_0146_ ? _0465_ : _0467_);
	assign _0469_ = (\mchip.pong.game.vga.pix_ind [0] ? _0468_ : _0464_);
	assign _0470_ = (_1103_ ? _0458_ : _0469_);
	assign _0471_ = (_0044_ ? _0434_ : _0470_);
	assign _0472_ = (_4389_ ? _4372_ : _4427_);
	assign _0473_ = (_4423_ ? _4417_ : _0472_);
	assign _0474_ = _4389_ & ~_0065_;
	assign _0475_ = ~_0474_;
	assign _0476_ = (_4387_ ? _0107_ : _0475_);
	assign _0477_ = (_0127_ ? _0473_ : _0476_);
	assign _0478_ = _4380_ & ~_4424_;
	assign _0479_ = ~_0478_;
	assign _0480_ = _0479_ | _4423_;
	assign _0481_ = (_4387_ ? _4380_ : _4434_);
	assign _0482_ = (_0127_ ? _0480_ : _0481_);
	assign _0483_ = (_0146_ ? _0477_ : _0482_);
	assign _0484_ = _4387_ & ~_4389_;
	assign _0485_ = (_4389_ ? _4374_ : _0065_);
	assign _0486_ = _0485_ | _4387_;
	assign _0487_ = (_0127_ ? _0484_ : _0486_);
	assign _0488_ = _4423_ | ~_0035_;
	assign _0489_ = (_4380_ ? _4427_ : _4407_);
	assign _0490_ = ~_0489_;
	assign _0491_ = (_4387_ ? _4380_ : _0490_);
	assign _0492_ = (_0127_ ? _0488_ : _0491_);
	assign _0493_ = (_0146_ ? _0487_ : _0492_);
	assign _0494_ = (\mchip.pong.game.vga.pix_ind [0] ? _0493_ : _0483_);
	assign _0495_ = ~_0153_;
	assign _0496_ = (_4423_ ? _4428_ : _0495_);
	assign _0497_ = (_4389_ ? _4408_ : _4427_);
	assign _0498_ = (_4423_ ? _0412_ : _0497_);
	assign _0499_ = (_0127_ ? _0496_ : _0498_);
	assign _0500_ = _4387_ & ~_0114_;
	assign _0501_ = ~_0500_;
	assign _0502_ = (_4389_ ? _4412_ : _0276_);
	assign _0503_ = ~_0502_;
	assign _0504_ = (_0127_ ? _0501_ : _0503_);
	assign _0505_ = (_0146_ ? _0499_ : _0504_);
	assign _0506_ = (_4371_ ? _4380_ : _4374_);
	assign _0507_ = (_4423_ ? _0107_ : _0506_);
	assign _0508_ = (_4387_ ? _0114_ : _4425_);
	assign _0509_ = (_0127_ ? _0507_ : _0508_);
	assign _0510_ = ~(_0502_ & _0056_);
	assign _0511_ = (_0146_ ? _0509_ : _0510_);
	assign _0512_ = (\mchip.pong.game.vga.pix_ind [0] ? _0511_ : _0505_);
	assign _0513_ = (_1103_ ? _0494_ : _0512_);
	assign _0514_ = ~_0426_;
	assign _0515_ = (_0276_ ? _0066_ : _0514_);
	assign _0516_ = _0474_ | _0366_;
	assign _0517_ = (_4387_ ? _0207_ : _0516_);
	assign _0518_ = (_0127_ ? _0515_ : _0517_);
	assign _0519_ = _4387_ & ~_4427_;
	assign _0520_ = ~_0519_;
	assign _0521_ = (_4389_ ? _0065_ : _4372_);
	assign _0522_ = ~_0521_;
	assign _0523_ = (_4423_ ? _0206_ : _0522_);
	assign _0524_ = (_0127_ ? _0520_ : _0523_);
	assign _0525_ = (_0146_ ? _0518_ : _0524_);
	assign _0526_ = (_4387_ ? _0203_ : _0066_);
	assign _0527_ = (_4423_ ? _0314_ : _0475_);
	assign _0528_ = (_0127_ ? _0526_ : _0527_);
	assign _0529_ = _0259_ & ~_4389_;
	assign _0530_ = ~_0529_;
	assign _0531_ = _4387_ & ~_0530_;
	assign _0532_ = ~_0531_;
	assign _0533_ = (_0056_ ? _0523_ : _0532_);
	assign _0534_ = (_0146_ ? _0528_ : _0533_);
	assign _0535_ = (\mchip.pong.game.vga.pix_ind [0] ? _0534_ : _0525_);
	assign _0536_ = (_4423_ ? _4417_ : _0054_);
	assign _0537_ = (_4387_ ? _0207_ : _0475_);
	assign _0538_ = (_0127_ ? _0536_ : _0537_);
	assign _0539_ = (_4389_ ? _4375_ : _0259_);
	assign _0540_ = ~_0539_;
	assign _0541_ = _0540_ | ~_4387_;
	assign _0542_ = (_4374_ ? _4371_ : _4380_);
	assign _0543_ = (_4387_ ? _0542_ : _0514_);
	assign _0544_ = (_0127_ ? _0541_ : _0543_);
	assign _0545_ = (_0146_ ? _0538_ : _0544_);
	assign _0546_ = (_4380_ ? _0425_ : _0065_);
	assign _0547_ = (_4387_ ? _0207_ : _0546_);
	assign _0548_ = (_0127_ ? _0536_ : _0547_);
	assign _0549_ = ~(_4443_ | _4423_);
	assign _0550_ = ~_0549_;
	assign _0551_ = (_4389_ ? _4419_ : _0425_);
	assign _0552_ = (_4423_ ? _0206_ : _0551_);
	assign _0553_ = (_0127_ ? _0550_ : _0552_);
	assign _0554_ = (_0146_ ? _0548_ : _0553_);
	assign _0555_ = (\mchip.pong.game.vga.pix_ind [0] ? _0554_ : _0545_);
	assign _0556_ = (_1103_ ? _0535_ : _0555_);
	assign _0557_ = (_0044_ ? _0513_ : _0556_);
	assign _0558_ = (_0088_ ? _0471_ : _0557_);
	assign _0559_ = (_4368_ ? _0398_ : _0558_);
	assign _0560_ = (_4380_ ? _4372_ : _4427_);
	assign _0561_ = (_4387_ ? _4380_ : _0560_);
	assign _0562_ = (_4423_ ? _0372_ : _0093_);
	assign _0563_ = (_0127_ ? _0561_ : _0562_);
	assign _0564_ = (_4423_ ? _4409_ : _0067_);
	assign _0565_ = (_0127_ ? _0162_ : _0564_);
	assign _0566_ = (_0146_ ? _0563_ : _0565_);
	assign _0567_ = _0459_ | _0272_;
	assign _0568_ = ~_0417_;
	assign _0569_ = (_4389_ ? _4374_ : _4371_);
	assign _0570_ = (_4423_ ? _0568_ : _0569_);
	assign _0571_ = (_0127_ ? _0567_ : _0570_);
	assign _0572_ = _0435_ | ~_4387_;
	assign _0573_ = (_4423_ ? _4409_ : _0404_);
	assign _0574_ = (_0127_ ? _0572_ : _0573_);
	assign _0575_ = (_0146_ ? _0571_ : _0574_);
	assign _0576_ = (\mchip.pong.game.vga.pix_ind [0] ? _0575_ : _0566_);
	assign _0577_ = ~_4374_;
	assign _0578_ = (_4389_ ? _0577_ : _4408_);
	assign _0579_ = (_4374_ ? _4372_ : _4389_);
	assign _0580_ = (_4423_ ? _0579_ : _0578_);
	assign _0581_ = (_0127_ ? _0567_ : _0580_);
	assign _0582_ = ~_4433_;
	assign _0583_ = (_4380_ ? _4408_ : _0582_);
	assign _0584_ = (_4423_ ? _0206_ : _0583_);
	assign _0585_ = (_0127_ ? _0520_ : _0584_);
	assign _0586_ = (_0146_ ? _0581_ : _0585_);
	assign _0587_ = (_4387_ ? _0054_ : _0066_);
	assign _0588_ = (_4423_ ? _0583_ : _4410_);
	assign _0590_ = (_0127_ ? _0587_ : _0588_);
	assign _0591_ = _4387_ & ~_0093_;
	assign _0592_ = ~_0591_;
	assign _0593_ = (_4423_ ? _4424_ : _0583_);
	assign _0594_ = (_0127_ ? _0592_ : _0593_);
	assign _0595_ = (_0146_ ? _0590_ : _0594_);
	assign _0596_ = (\mchip.pong.game.vga.pix_ind [0] ? _0595_ : _0586_);
	assign _0597_ = (_1103_ ? _0576_ : _0596_);
	assign _0598_ = (_4380_ ? _4371_ : _0259_);
	assign _0599_ = ~_0598_;
	assign _0601_ = _0361_ | _4409_;
	assign _0602_ = (_4423_ ? _0601_ : _0599_);
	assign _0603_ = _0361_ | _0066_;
	assign _0604_ = (_4423_ ? _0603_ : _0446_);
	assign _0605_ = (_0127_ ? _0602_ : _0604_);
	assign _0606_ = (_4380_ ? _4374_ : _0425_);
	assign _0607_ = _0606_ | _4423_;
	assign _0608_ = (_4389_ ? _4408_ : _4375_);
	assign _0609_ = (_4423_ ? _0153_ : _0608_);
	assign _0610_ = (_0127_ ? _0607_ : _0609_);
	assign _0612_ = (_0146_ ? _0605_ : _0610_);
	assign _0613_ = (_4380_ ? _4424_ : _4408_);
	assign _0614_ = (_4387_ ? _4437_ : _0613_);
	assign _0615_ = (_4389_ ? _4371_ : _4419_);
	assign _0616_ = (_4423_ ? _0119_ : _0615_);
	assign _0617_ = (_0127_ ? _0614_ : _0616_);
	assign _0618_ = _4387_ & ~_0472_;
	assign _0619_ = ~_0618_;
	assign _0620_ = (_4380_ ? _4371_ : _4375_);
	assign _0621_ = (_4389_ ? _4433_ : _0065_);
	assign _0623_ = ~_0621_;
	assign _0624_ = (_4423_ ? _0623_ : _0620_);
	assign _0625_ = (_0127_ ? _0619_ : _0624_);
	assign _0626_ = (_0146_ ? _0617_ : _0625_);
	assign _0627_ = (\mchip.pong.game.vga.pix_ind [0] ? _0626_ : _0612_);
	assign _0628_ = _0361_ | _4443_;
	assign _0629_ = (_4423_ ? _0628_ : _0506_);
	assign _0630_ = _0361_ | _0100_;
	assign _0631_ = (_4389_ ? _4408_ : _0065_);
	assign _0632_ = (_4423_ ? _0631_ : _0630_);
	assign _0634_ = (_0127_ ? _0629_ : _0632_);
	assign _0635_ = (_4423_ ? _4443_ : _0090_);
	assign _0636_ = (_0127_ ? _0520_ : _0635_);
	assign _0637_ = (_0146_ ? _0634_ : _0636_);
	assign _0638_ = (_4423_ ? _4427_ : _0506_);
	assign _0639_ = (_4380_ ? _0065_ : _4408_);
	assign _0640_ = (_4423_ ? _0372_ : _0639_);
	assign _0641_ = (_0127_ ? _0638_ : _0640_);
	assign _0642_ = (_4423_ ? _0446_ : _0207_);
	assign _0643_ = (_0127_ ? _0193_ : _0642_);
	assign _0645_ = (_0146_ ? _0641_ : _0643_);
	assign _0646_ = (\mchip.pong.game.vga.pix_ind [0] ? _0645_ : _0637_);
	assign _0647_ = (_1103_ ? _0627_ : _0646_);
	assign _0648_ = (_0044_ ? _0597_ : _0647_);
	assign _0649_ = (_4387_ ? _4381_ : _0446_);
	assign _0650_ = (_4423_ ? _0421_ : _0403_);
	assign _0651_ = (_0127_ ? _0649_ : _0650_);
	assign _0652_ = (_0127_ ? _0048_ : _0160_);
	assign _0653_ = (_0146_ ? _0651_ : _0652_);
	assign _0654_ = _4433_ & ~_4389_;
	assign _0656_ = ~_0654_;
	assign _0657_ = (_4387_ ? _0153_ : _0656_);
	assign _0658_ = (_4387_ ? _0403_ : _0560_);
	assign _0659_ = (_0127_ ? _0657_ : _0658_);
	assign _0660_ = (_4389_ ? _4374_ : _4407_);
	assign _0661_ = (_4423_ ? _0454_ : _0660_);
	assign _0662_ = (_0056_ ? _0429_ : _0661_);
	assign _0663_ = (_0146_ ? _0659_ : _0662_);
	assign _0664_ = (\mchip.pong.game.vga.pix_ind [0] ? _0663_ : _0653_);
	assign _0665_ = ~_0093_;
	assign _0667_ = (_4387_ ? _0665_ : _0656_);
	assign _0668_ = (_4387_ ? _4443_ : _4391_);
	assign _0669_ = (_0127_ ? _0667_ : _0668_);
	assign _0670_ = ~_0181_;
	assign _0671_ = _4389_ & ~_0259_;
	assign _0672_ = _0671_ | _0417_;
	assign _0673_ = (_4423_ ? _0451_ : _0672_);
	assign _0674_ = (_0056_ ? _0670_ : _0673_);
	assign _0675_ = (_0146_ ? _0669_ : _0674_);
	assign _0676_ = (_4387_ ? _0054_ : _0601_);
	assign _0678_ = (_4380_ ? _4419_ : _4427_);
	assign _0679_ = (_4423_ ? _0678_ : _0446_);
	assign _0680_ = (_0127_ ? _0676_ : _0679_);
	assign _0681_ = _0572_ & _0127_;
	assign _0682_ = _0238_ | _0681_;
	assign _0683_ = (_0146_ ? _0680_ : _0682_);
	assign _0684_ = (\mchip.pong.game.vga.pix_ind [0] ? _0683_ : _0675_);
	assign _0685_ = (_1103_ ? _0664_ : _0684_);
	assign _0686_ = (_4387_ ? _4389_ : _0435_);
	assign _0687_ = (_4380_ ? _4375_ : _0582_);
	assign _0689_ = (_4423_ ? _0615_ : _0687_);
	assign _0690_ = (_0127_ ? _0686_ : _0689_);
	assign _0691_ = (_0146_ ? _0690_ : _0242_);
	assign _0692_ = (_4387_ ? _4434_ : _0579_);
	assign _0693_ = (_4387_ ? _0117_ : _0107_);
	assign _0694_ = (_0127_ ? _0692_ : _0693_);
	assign _0695_ = (_0146_ ? _0694_ : _0126_);
	assign _0696_ = (\mchip.pong.game.vga.pix_ind [0] ? _0695_ : _0691_);
	assign _0697_ = (_4423_ ? _4389_ : _0153_);
	assign _0698_ = (_4423_ ? _0101_ : _0579_);
	assign _0700_ = (_0127_ ? _0697_ : _0698_);
	assign _0701_ = (_0146_ ? _0700_ : _0156_);
	assign _0702_ = (_4423_ ? _4389_ : _4409_);
	assign _0703_ = ~_0401_;
	assign _0704_ = (_4387_ ? _0703_ : _0093_);
	assign _0705_ = (_0127_ ? _0702_ : _0704_);
	assign _0706_ = (_0056_ ? _0420_ : _0399_);
	assign _0707_ = (_0146_ ? _0705_ : _0706_);
	assign _0708_ = (\mchip.pong.game.vga.pix_ind [0] ? _0707_ : _0701_);
	assign _0709_ = (_1103_ ? _0696_ : _0708_);
	assign _0711_ = (_0044_ ? _0685_ : _0709_);
	assign _0712_ = (_0088_ ? _0648_ : _0711_);
	assign _0713_ = (_4387_ ? _0113_ : _0404_);
	assign _0714_ = _0127_ & ~_0713_;
	assign _0715_ = (_0146_ ? _0714_ : _0340_);
	assign _0716_ = (\mchip.pong.game.vga.pix_ind [0] ? _0715_ : _0339_);
	assign _0717_ = (_1103_ ? _0337_ : _0716_);
	assign _0718_ = (_0044_ ? _0717_ : _0329_);
	assign _0719_ = (_0088_ ? _0718_ : _0307_);
	assign _0720_ = (_4368_ ? _0712_ : _0719_);
	assign _0722_ = (_4367_ ? _0559_ : _0720_);
	assign _0723_ = \mchip.pong.sync.o_out [0] & ~\mchip.pong.sync.o_out [1];
	assign _0724_ = _0128_ & ~_0056_;
	assign _0725_ = ~_0724_;
	assign _0726_ = ~(_0119_ & _4387_);
	assign _0727_ = ~_0726_;
	assign _0728_ = (_4387_ ? _0454_ : _0035_);
	assign _0729_ = (_0127_ ? _0727_ : _0728_);
	assign _0730_ = (_0146_ ? _0725_ : _0729_);
	assign _0731_ = _0127_ & ~_0686_;
	assign _0733_ = ~_0731_;
	assign _0734_ = (_0127_ ? _4387_ : _0420_);
	assign _0735_ = (_0146_ ? _0733_ : _0734_);
	assign _0736_ = (\mchip.pong.game.vga.pix_ind [0] ? _0735_ : _0730_);
	assign _0737_ = _0143_ | _0056_;
	assign _0738_ = (_4387_ ? _0295_ : _0119_);
	assign _0739_ = (_0056_ ? _0120_ : _0738_);
	assign _0740_ = (_0146_ ? _0737_ : _0739_);
	assign _0741_ = \mchip.pong.game.vga.pix_ind [0] & ~_0740_;
	assign _0742_ = _4423_ | _4381_;
	assign _0743_ = (_4387_ ? _0118_ : _4437_);
	assign _0744_ = (_0056_ ? _0742_ : _0743_);
	assign _0745_ = (_4387_ ? _4407_ : _0054_);
	assign _0746_ = (_0056_ ? _0383_ : _0745_);
	assign _0747_ = (_0146_ ? _0744_ : _0746_);
	assign _0748_ = _0747_ & ~\mchip.pong.game.vga.pix_ind [0];
	assign _0749_ = _0748_ | _0741_;
	assign _0750_ = (_1103_ ? _0736_ : _0749_);
	assign _0751_ = (_0044_ ? _0124_ : _0750_);
	assign _0752_ = (_0088_ ? _0084_ : _0751_);
	assign _0754_ = _4437_ & _4387_;
	assign _0755_ = ~_0754_;
	assign _0756_ = ~_0259_;
	assign _0757_ = (_4380_ ? _4407_ : _0756_);
	assign _0758_ = (_4387_ ? _0153_ : _0757_);
	assign _0759_ = (_0056_ ? _0755_ : _0758_);
	assign _0760_ = (_4387_ ? _4380_ : _0603_);
	assign _0761_ = (_4387_ ? _0117_ : _0391_);
	assign _0762_ = ~_0761_;
	assign _0763_ = (_0127_ ? _0760_ : _0762_);
	assign _0765_ = (_0146_ ? _0759_ : _0763_);
	assign _0766_ = (_4423_ ? _0131_ : _0113_);
	assign _0767_ = (_0127_ ? _0162_ : _0766_);
	assign _0768_ = ~_0767_;
	assign _0769_ = (_4387_ ? _4389_ : _0401_);
	assign _0770_ = (_4387_ ? _0035_ : _0153_);
	assign _0771_ = (_0127_ ? _0769_ : _0770_);
	assign _0772_ = (_0146_ ? _0768_ : _0771_);
	assign _0773_ = (\mchip.pong.game.vga.pix_ind [0] ? _0772_ : _0765_);
	assign _0774_ = (_0127_ ? _0166_ : _0500_);
	assign _0776_ = ~_0774_;
	assign _0777_ = _4428_ | _4387_;
	assign _0778_ = (_4423_ ? _0054_ : _0035_);
	assign _0779_ = (_0127_ ? _0777_ : _0778_);
	assign _0780_ = (_0146_ ? _0776_ : _0779_);
	assign _0781_ = _0127_ & ~_0697_;
	assign _0782_ = ~_0781_;
	assign _0783_ = _4387_ & ~_4417_;
	assign _0784_ = (_4387_ ? _0054_ : _4381_);
	assign _0785_ = (_0127_ ? _0783_ : _0784_);
	assign _0787_ = (_0146_ ? _0782_ : _0785_);
	assign _0788_ = (\mchip.pong.game.vga.pix_ind [0] ? _0787_ : _0780_);
	assign _0789_ = (_1103_ ? _0773_ : _0788_);
	assign _0790_ = (_4389_ ? _4423_ : _4424_);
	assign _0791_ = (_0056_ ? _4387_ : _0790_);
	assign _0792_ = ~_0114_;
	assign _0793_ = (_4423_ ? _4443_ : _0792_);
	assign _0794_ = (_0127_ ? _0488_ : _0793_);
	assign _0795_ = (_0146_ ? _0791_ : _0794_);
	assign _0796_ = (_4423_ ? _0066_ : _4381_);
	assign _0797_ = _0796_ | _0056_;
	assign _0798_ = (_4423_ ? _0153_ : _0792_);
	assign _0799_ = _0798_ | _0127_;
	assign _0800_ = (_0146_ ? _0797_ : _0799_);
	assign _0801_ = (\mchip.pong.game.vga.pix_ind [0] ? _0800_ : _0795_);
	assign _0802_ = (_0056_ ? _0193_ : _0784_);
	assign _0803_ = (_0146_ ? _0802_ : _0799_);
	assign _0804_ = _0179_ | ~_0046_;
	assign _0805_ = _0421_ & ~_4387_;
	assign _0806_ = (_0127_ ? _0804_ : _0805_);
	assign _0808_ = (_4389_ ? _4372_ : _0756_);
	assign _0809_ = _0808_ | _4387_;
	assign _0810_ = (_4387_ ? _0035_ : _4409_);
	assign _0811_ = (_0127_ ? _0809_ : _0810_);
	assign _0812_ = (_0146_ ? _0806_ : _0811_);
	assign _0813_ = (\mchip.pong.game.vga.pix_ind [0] ? _0812_ : _0803_);
	assign _0814_ = (_1103_ ? _0801_ : _0813_);
	assign _0815_ = (_0044_ ? _0789_ : _0814_);
	assign _0816_ = (_4387_ ? _0054_ : _0479_);
	assign _0817_ = (_4423_ ? _0035_ : _0372_);
	assign _0819_ = (_0127_ ? _0816_ : _0817_);
	assign _0820_ = (_4380_ ? _4419_ : _4407_);
	assign _0821_ = _0403_ | _0366_;
	assign _0822_ = (_4423_ ? _0821_ : _0820_);
	assign _0823_ = (_4387_ ? _0792_ : _4434_);
	assign _0824_ = (_0127_ ? _0822_ : _0823_);
	assign _0825_ = (_0146_ ? _0819_ : _0824_);
	assign _0826_ = (_4389_ ? _4372_ : _4424_);
	assign _0827_ = (_4387_ ? _4380_ : _0826_);
	assign _0828_ = ~(_0639_ | _4423_);
	assign _0830_ = ~_0828_;
	assign _0831_ = (_0127_ ? _0827_ : _0830_);
	assign _0832_ = (_4423_ ? _0474_ : _0401_);
	assign _0833_ = ~_0832_;
	assign _0834_ = (_4387_ ? _0792_ : _4409_);
	assign _0835_ = (_0127_ ? _0833_ : _0834_);
	assign _0836_ = (_0146_ ? _0831_ : _0835_);
	assign _0837_ = (\mchip.pong.game.vga.pix_ind [0] ? _0836_ : _0825_);
	assign _0838_ = (_4387_ ? _0035_ : _0444_);
	assign _0839_ = (_4380_ ? _4424_ : _4407_);
	assign _0841_ = ~_0839_;
	assign _0842_ = (_4423_ ? _0421_ : _0841_);
	assign _0843_ = (_0127_ ? _0838_ : _0842_);
	assign _0844_ = (_4423_ ? _0093_ : _0560_);
	assign _0845_ = ~_4380_;
	assign _0846_ = (_4423_ ? _0845_ : _0203_);
	assign _0847_ = (_0127_ ? _0844_ : _0846_);
	assign _0848_ = (_0146_ ? _0843_ : _0847_);
	assign _0849_ = _0035_ ^ _4423_;
	assign _0850_ = _4380_ & _4427_;
	assign _0852_ = ~_0850_;
	assign _0853_ = (_4423_ ? _0852_ : _0435_);
	assign _0854_ = (_0127_ ? _0849_ : _0853_);
	assign _0855_ = (_4423_ ? _0421_ : _4428_);
	assign _0856_ = (_4423_ ? _0845_ : _4428_);
	assign _0857_ = (_0127_ ? _0855_ : _0856_);
	assign _0858_ = (_0146_ ? _0854_ : _0857_);
	assign _0859_ = (\mchip.pong.game.vga.pix_ind [0] ? _0858_ : _0848_);
	assign _0860_ = (_1103_ ? _0837_ : _0859_);
	assign _0861_ = (_4387_ ? _0203_ : _0454_);
	assign _0863_ = (_4423_ ? _0542_ : _0472_);
	assign _0864_ = (_0127_ ? _0861_ : _0863_);
	assign _0865_ = (_4389_ ? _0065_ : _0577_);
	assign _0866_ = _0865_ | _4423_;
	assign _0867_ = (_4423_ ? _0206_ : _0792_);
	assign _0868_ = (_0127_ ? _0866_ : _0867_);
	assign _0869_ = (_0146_ ? _0864_ : _0868_);
	assign _0870_ = (_4387_ ? _0203_ : _4407_);
	assign _0871_ = ~(_4389_ & _4371_);
	assign _0872_ = _0871_ | _4387_;
	assign _0874_ = (_0127_ ? _0870_ : _0872_);
	assign _0875_ = _4387_ & ~_0421_;
	assign _0876_ = ~_0875_;
	assign _0877_ = (_0127_ ? _0876_ : _0867_);
	assign _0878_ = (_0146_ ? _0874_ : _0877_);
	assign _0879_ = (\mchip.pong.game.vga.pix_ind [0] ? _0878_ : _0869_);
	assign _0880_ = (_4374_ ? _4389_ : _4372_);
	assign _0881_ = (_4387_ ? _0054_ : _0880_);
	assign _0882_ = _0259_ & ~_4380_;
	assign _0883_ = ~_0882_;
	assign _0885_ = _0883_ | _4387_;
	assign _0886_ = (_0127_ ? _0881_ : _0885_);
	assign _0887_ = (_0127_ ? _0501_ : _0867_);
	assign _0888_ = (_0146_ ? _0886_ : _0887_);
	assign _0889_ = (_4387_ ? _0054_ : _0671_);
	assign _0890_ = (_4380_ ? _0425_ : _0756_);
	assign _0891_ = _0890_ | _4387_;
	assign _0892_ = (_0127_ ? _0889_ : _0891_);
	assign _0893_ = (_4423_ ? _0107_ : _0114_);
	assign _0894_ = (_0056_ ? _0867_ : _0893_);
	assign _0896_ = (_0146_ ? _0892_ : _0894_);
	assign _0897_ = (\mchip.pong.game.vga.pix_ind [0] ? _0896_ : _0888_);
	assign _0898_ = (_1103_ ? _0879_ : _0897_);
	assign _0899_ = (_0044_ ? _0860_ : _0898_);
	assign _0900_ = (_0088_ ? _0815_ : _0899_);
	assign _0901_ = (_4368_ ? _0752_ : _0900_);
	assign _0902_ = _0203_ | _4423_;
	assign _0903_ = ~_0254_;
	assign _0904_ = (_4387_ ? _4380_ : _0903_);
	assign _0905_ = (_0056_ ? _0902_ : _0904_);
	assign _0907_ = (_0127_ ? _0726_ : _0834_);
	assign _0908_ = (_0146_ ? _0905_ : _0907_);
	assign _0909_ = (_0127_ ? _0459_ : _0902_);
	assign _0910_ = (_0127_ ? _0572_ : _0834_);
	assign _0911_ = (_0146_ ? _0909_ : _0910_);
	assign _0912_ = (\mchip.pong.game.vga.pix_ind [0] ? _0911_ : _0908_);
	assign _0913_ = (_4387_ ? _0054_ : _4437_);
	assign _0914_ = _0361_ | _4423_;
	assign _0915_ = (_0127_ ? _0913_ : _0914_);
	assign _0916_ = (_4387_ ? _0451_ : _0114_);
	assign _0917_ = (_0056_ ? _0867_ : _0916_);
	assign _0918_ = (_0146_ ? _0915_ : _0917_);
	assign _0919_ = (_4423_ ? _0421_ : _0299_);
	assign _0920_ = (_0056_ ? _0867_ : _0919_);
	assign _0921_ = (_0146_ ? _0915_ : _0920_);
	assign _0922_ = (\mchip.pong.game.vga.pix_ind [0] ? _0921_ : _0918_);
	assign _0923_ = (_1103_ ? _0912_ : _0922_);
	assign _0924_ = (_4387_ ? _4381_ : _0479_);
	assign _0925_ = (_4423_ ? _4391_ : _0035_);
	assign _0926_ = (_0127_ ? _0924_ : _0925_);
	assign _0928_ = _0678_ | _4423_;
	assign _0929_ = (_4387_ ? _4390_ : _0153_);
	assign _0930_ = (_0127_ ? _0928_ : _0929_);
	assign _0931_ = (_0146_ ? _0926_ : _0930_);
	assign _0932_ = (_4387_ ? _4437_ : _0114_);
	assign _0933_ = (_4423_ ? _4391_ : _0792_);
	assign _0934_ = (_0127_ ? _0932_ : _0933_);
	assign _0935_ = (_0127_ ? _0550_ : _0823_);
	assign _0936_ = (_0146_ ? _0934_ : _0935_);
	assign _0937_ = (\mchip.pong.game.vga.pix_ind [0] ? _0936_ : _0931_);
	assign _0939_ = (_4423_ ? _0066_ : _0035_);
	assign _0940_ = (_4423_ ? _0421_ : _0792_);
	assign _0941_ = (_0127_ ? _0939_ : _0940_);
	assign _0942_ = (_4387_ ? _4428_ : _4443_);
	assign _0943_ = _0056_ & ~_0942_;
	assign _0944_ = ~_0943_;
	assign _0945_ = (_0146_ ? _0941_ : _0944_);
	assign _0946_ = (_4423_ ? _0671_ : _0035_);
	assign _0947_ = (_0056_ ? _0940_ : _0946_);
	assign _0948_ = (_4423_ ? _4389_ : _0792_);
	assign _0950_ = _0056_ & ~_0948_;
	assign _0951_ = ~_0950_;
	assign _0952_ = (_0146_ ? _0947_ : _0951_);
	assign _0953_ = (\mchip.pong.game.vga.pix_ind [0] ? _0952_ : _0945_);
	assign _0954_ = (_1103_ ? _0937_ : _0953_);
	assign _0955_ = (_0044_ ? _0923_ : _0954_);
	assign _0956_ = (_4387_ ? _4381_ : _0114_);
	assign _0957_ = (_4371_ ? _4374_ : _4380_);
	assign _0958_ = (_4387_ ? _4407_ : _0957_);
	assign _0959_ = (_0127_ ? _0956_ : _0958_);
	assign _0961_ = ~_4437_;
	assign _0962_ = (_4423_ ? _0070_ : _0961_);
	assign _0963_ = (_4423_ ? _0153_ : _0090_);
	assign _0964_ = (_0127_ ? _0962_ : _0963_);
	assign _0965_ = (_0146_ ? _0959_ : _0964_);
	assign _0966_ = (_4423_ ? _0100_ : _0153_);
	assign _0967_ = _4423_ | ~_0101_;
	assign _0968_ = (_0127_ ? _0966_ : _0967_);
	assign _0969_ = (_4423_ ? _0119_ : _0107_);
	assign _0970_ = ~_4389_;
	assign _0972_ = (_4387_ ? _0970_ : _4381_);
	assign _0973_ = (_0127_ ? _0969_ : _0972_);
	assign _0974_ = (_0146_ ? _0968_ : _0973_);
	assign _0975_ = (\mchip.pong.game.vga.pix_ind [0] ? _0974_ : _0965_);
	assign _0976_ = (_4387_ ? _0665_ : _0114_);
	assign _0977_ = (_4423_ ? _0421_ : _4390_);
	assign _0978_ = (_0127_ ? _0976_ : _0977_);
	assign _0979_ = (_4389_ ? _4372_ : _0065_);
	assign _0980_ = _0979_ | _4423_;
	assign _0981_ = (_4423_ ? _4409_ : _0035_);
	assign _0983_ = (_0127_ ? _0980_ : _0981_);
	assign _0984_ = (_0146_ ? _0978_ : _0983_);
	assign _0985_ = (_4387_ ? _0054_ : _0560_);
	assign _0986_ = _4391_ ^ _4387_;
	assign _0987_ = (_0127_ ? _0985_ : _0986_);
	assign _0988_ = (_4387_ ? _0090_ : _0582_);
	assign _0989_ = _4409_ | ~_0093_;
	assign _0990_ = (_4387_ ? _0361_ : _0989_);
	assign _0991_ = (_0127_ ? _0988_ : _0990_);
	assign _0992_ = (_0146_ ? _0987_ : _0991_);
	assign _0994_ = (\mchip.pong.game.vga.pix_ind [0] ? _0992_ : _0984_);
	assign _0995_ = (_1103_ ? _0975_ : _0994_);
	assign _0996_ = (_4387_ ? _0845_ : _4390_);
	assign _0997_ = (_0056_ ? _0193_ : _0996_);
	assign _0998_ = ~_0108_;
	assign _0999_ = (_4423_ ? _0035_ : _0578_);
	assign _1000_ = (_0056_ ? _0998_ : _0999_);
	assign _1001_ = (_0146_ ? _0997_ : _1000_);
	assign _1002_ = ~_4434_;
	assign _1003_ = (_4387_ ? _1002_ : _0506_);
	assign _1005_ = ~_1003_;
	assign _1006_ = (_4423_ ? _0451_ : _0852_);
	assign _1007_ = (_0127_ ? _1005_ : _1006_);
	assign _1008_ = _0065_ ^ _4380_;
	assign _1009_ = (_4389_ ? _4427_ : _4407_);
	assign _1010_ = ~_1009_;
	assign _1011_ = (_4423_ ? _1010_ : _1008_);
	assign _1012_ = (_4387_ ? _0903_ : _0035_);
	assign _1013_ = (_0127_ ? _1011_ : _1012_);
	assign _1014_ = (_0146_ ? _1007_ : _1013_);
	assign _1015_ = (\mchip.pong.game.vga.pix_ind [0] ? _1014_ : _1001_);
	assign _1016_ = (_4387_ ? _4389_ : _0067_);
	assign _1017_ = (_0127_ ? _0154_ : _1016_);
	assign _1018_ = (_4389_ ? _0425_ : _4408_);
	assign _1019_ = (_4423_ ? _4371_ : _1018_);
	assign _1020_ = (_4380_ ? _4407_ : _4375_);
	assign _1021_ = (_4423_ ? _4381_ : _1020_);
	assign _1022_ = (_0127_ ? _1019_ : _1021_);
	assign _1023_ = (_0146_ ? _1017_ : _1022_);
	assign _1024_ = ~(_0101_ & _0871_);
	assign _1025_ = (_4387_ ? _4409_ : _1024_);
	assign _1026_ = (_4387_ ? _1024_ : _0451_);
	assign _1027_ = (_0127_ ? _1025_ : _1026_);
	assign _1028_ = (_4374_ ? _4389_ : _4371_);
	assign _1029_ = (_4423_ ? _0391_ : _1028_);
	assign _1030_ = (_4389_ ? _4375_ : _0577_);
	assign _1031_ = (_4423_ ? _0054_ : _1030_);
	assign _1032_ = (_0127_ ? _1029_ : _1031_);
	assign _1033_ = (_0146_ ? _1027_ : _1032_);
	assign _1034_ = (\mchip.pong.game.vga.pix_ind [0] ? _1033_ : _1023_);
	assign _1035_ = (_1103_ ? _1015_ : _1034_);
	assign _1036_ = (_0044_ ? _0995_ : _1035_);
	assign _1037_ = (_0088_ ? _0955_ : _1036_);
	assign _1038_ = (_4387_ ? _4417_ : _0540_);
	assign _1039_ = (_4423_ ? _0093_ : _0404_);
	assign _1040_ = (_0127_ ? _1038_ : _1039_);
	assign _1041_ = ~(_4423_ | _4427_);
	assign _1042_ = (_0056_ ? _0386_ : _1041_);
	assign _1043_ = (_0146_ ? _1040_ : _1042_);
	assign _1044_ = (_4387_ ? _4443_ : _1024_);
	assign _1046_ = (_4423_ ? _0451_ : _0880_);
	assign _1047_ = (_0127_ ? _1044_ : _1046_);
	assign _1048_ = (_4423_ ? _0314_ : _0871_);
	assign _1049_ = (_0056_ ? _0383_ : _1048_);
	assign _1050_ = (_0146_ ? _1047_ : _1049_);
	assign _1051_ = (\mchip.pong.game.vga.pix_ind [0] ? _1050_ : _1043_);
	assign _1052_ = (_1103_ ? _0337_ : _1051_);
	assign _1053_ = (_0044_ ? _1052_ : _0329_);
	assign _1054_ = (_0088_ ? _1053_ : _0307_);
	assign _1055_ = (_4368_ ? _1037_ : _1054_);
	assign _1057_ = (_4367_ ? _0901_ : _1055_);
	assign _1058_ = \mchip.pong.sync.o_out [1] & ~\mchip.pong.sync.o_out [0];
	assign _1059_ = (_1058_ ? _1057_ : _0347_);
	assign _1060_ = (_0723_ ? _0722_ : _1059_);
	assign _1061_ = ~(\mchip.pong.sync.o_out [1] | \mchip.pong.sync.o_out [0]);
	assign _1062_ = (_1061_ ? _0347_ : _1060_);
	assign _1063_ = ~(\mchip.pong.game.ball.dpath.ballX [7] & \mchip.pong.game.ball.dpath.ballX [6]);
	assign _1064_ = _1063_ | _1241_;
	assign _1065_ = _1241_ & ~_1063_;
	assign _1066_ = _1065_ & ~_1294_;
	assign _1068_ = _1064_ & ~_1066_;
	assign _1069_ = _1338_ & ~_1068_;
	assign _1070_ = ~_4239_;
	assign _1071_ = \mchip.pong.game.ball.dpath.ballX [8] & ~_1068_;
	assign _1072_ = _1071_ ^ \mchip.pong.game.ball.dpath.ballX [9];
	assign _1073_ = _1072_ ^ _1070_;
	assign _1074_ = ~\mchip.pong.game.ball.dpath.ballX [8];
	assign _1075_ = _1068_ ^ _1074_;
	assign _1076_ = _1075_ ^ _4237_;
	assign _1077_ = _1076_ | ~_1073_;
	assign _1079_ = ~(_1077_ | _1069_);
	assign _1080_ = ~_4243_;
	assign _1081_ = _1294_ & _1241_;
	assign _1082_ = \mchip.pong.game.ball.dpath.ballX [6] & ~_1081_;
	assign _1083_ = _1082_ ^ \mchip.pong.game.ball.dpath.ballX [7];
	assign _1084_ = _1083_ ^ _1080_;
	assign _1085_ = ~\mchip.pong.game.ball.dpath.ballX [6];
	assign _1086_ = _1081_ ^ _1085_;
	assign _1087_ = _1086_ ^ _4244_;
	assign _1088_ = _1084_ & ~_1087_;
	assign _1090_ = _1294_ ^ \mchip.pong.game.ball.dpath.ballX [4];
	assign _1091_ = _1090_ ^ _4333_;
	assign _1092_ = _1294_ & ~\mchip.pong.game.ball.dpath.ballX [4];
	assign _1093_ = _1092_ ^ \mchip.pong.game.ball.dpath.ballX [5];
	assign _1094_ = ~(_1093_ ^ _4365_);
	assign _1095_ = _1094_ | _1091_;
	assign _1096_ = _1088_ & ~_1095_;
	assign _1097_ = _3381_ ^ \mchip.pong.game.ball.dpath.ballX [3];
	assign _1098_ = _1097_ ^ _4330_;
	assign _1099_ = ~(\mchip.pong.game.ball.dpath.ballX [1] ^ \mchip.pong.game.ball.dpath.ballX [2]);
	assign _1101_ = _1099_ ^ \mchip.pong.game.vga.pix_ind [2];
	assign _1102_ = _1098_ & ~_1101_;
	assign _1104_ = \mchip.pong.game.vga.pix_ind [0] & ~_1103_;
	assign _1105_ = _1104_ & _1102_;
	assign _1106_ = ~(_1105_ & _1096_);
	assign _1107_ = _1079_ & ~_1106_;
	assign _1108_ = _1072_ | _1070_;
	assign _1109_ = _1075_ | ~_4237_;
	assign _1110_ = _1073_ & ~_1109_;
	assign _1112_ = _1108_ & ~_1110_;
	assign _1113_ = _1083_ | _1080_;
	assign _1114_ = _1086_ | ~_4244_;
	assign _1115_ = _1084_ & ~_1114_;
	assign _1116_ = _1113_ & ~_1115_;
	assign _1117_ = _1093_ | _4365_;
	assign _1118_ = _4333_ & ~_1090_;
	assign _1119_ = _1118_ & ~_1094_;
	assign _1120_ = _1117_ & ~_1119_;
	assign _1121_ = _1088_ & ~_1120_;
	assign _1123_ = _1116_ & ~_1121_;
	assign _1124_ = _1097_ | _4330_;
	assign _1125_ = _1099_ | _4328_;
	assign _1126_ = _1098_ & ~_1125_;
	assign _1127_ = _1124_ & ~_1126_;
	assign _1128_ = ~(\mchip.pong.game.vga.pix_ind [1] & \mchip.pong.game.ball.dpath.ballX [1]);
	assign _1129_ = _1128_ & ~_1104_;
	assign _1130_ = _1102_ & ~_1129_;
	assign _1131_ = _1127_ & ~_1130_;
	assign _1132_ = _1096_ & ~_1131_;
	assign _1134_ = _1123_ & ~_1132_;
	assign _1135_ = ~(_1134_ | _1077_);
	assign _1136_ = _1112_ & ~_1135_;
	assign _1137_ = _1136_ | _1069_;
	assign _1138_ = ~(_1137_ | _1107_);
	assign _1139_ = _4239_ ^ _3370_;
	assign _1140_ = _4237_ ^ \mchip.pong.game.ball.dpath.ballX [8];
	assign _1141_ = _1139_ & ~_1140_;
	assign _1142_ = _4243_ ^ _3271_;
	assign _1143_ = _4244_ ^ \mchip.pong.game.ball.dpath.ballX [6];
	assign _1145_ = _1142_ & ~_1143_;
	assign _1146_ = ~(_4366_ & _4362_);
	assign _1147_ = _1145_ & ~_1146_;
	assign _1148_ = _1103_ & ~\mchip.pong.game.vga.pix_ind [0];
	assign _1149_ = _1148_ & _4358_;
	assign _1150_ = _1149_ & _1147_;
	assign _1151_ = ~(_1150_ & _1141_);
	assign _1152_ = _4239_ | _3370_;
	assign _1153_ = _4237_ | _1074_;
	assign _1154_ = _1139_ & ~_1153_;
	assign _1156_ = _1152_ & ~_1154_;
	assign _1157_ = _4243_ | _3271_;
	assign _1158_ = _4244_ | _1085_;
	assign _1159_ = _1142_ & ~_1158_;
	assign _1160_ = _1157_ & ~_1159_;
	assign _1161_ = ~(_4365_ & \mchip.pong.game.ball.dpath.ballX [5]);
	assign _1162_ = _4366_ & _4361_;
	assign _1163_ = _1161_ & ~_1162_;
	assign _1164_ = _1145_ & ~_1163_;
	assign _1165_ = _1160_ & ~_1164_;
	assign _1167_ = _4352_ & _4356_;
	assign _1168_ = _4351_ & ~_1167_;
	assign _1169_ = _0043_ & ~_1148_;
	assign _1170_ = _4358_ & ~_1169_;
	assign _1171_ = _1168_ & ~_1170_;
	assign _1172_ = _1147_ & ~_1171_;
	assign _1173_ = _1165_ & ~_1172_;
	assign _1174_ = _1141_ & ~_1173_;
	assign _1175_ = _1156_ & ~_1174_;
	assign _1176_ = _1151_ & ~_1175_;
	assign _1178_ = _4230_ ^ _1622_;
	assign _1179_ = _1600_ & ~_1178_;
	assign _1180_ = _1805_ | ~_4216_;
	assign _1181_ = ~(_4216_ ^ _1805_);
	assign _1182_ = _1761_ | ~_4217_;
	assign _1183_ = _1181_ & ~_1182_;
	assign _1184_ = _1180_ & ~_1183_;
	assign _1185_ = _4217_ ^ _1761_;
	assign _1186_ = _1181_ & ~_1185_;
	assign _1187_ = _1675_ | ~_4220_;
	assign _1188_ = _4220_ ^ _1675_;
	assign _1189_ = _4221_ & ~_1697_;
	assign _1190_ = _1189_ & ~_1188_;
	assign _1191_ = _1187_ & ~_1190_;
	assign _1192_ = _1186_ & ~_1191_;
	assign _1193_ = _1184_ & ~_1192_;
	assign _1194_ = _4221_ ^ _1697_;
	assign _1195_ = _1194_ | _1188_;
	assign _1196_ = _1186_ & ~_1195_;
	assign _1197_ = _4205_ | _1871_;
	assign _1198_ = _4205_ ^ _1871_;
	assign _1199_ = _4206_ | _1893_;
	assign _1200_ = _1198_ & ~_1199_;
	assign _1201_ = _1197_ & ~_1200_;
	assign _1202_ = _4318_ ^ _1893_;
	assign _1203_ = _1198_ & ~_1202_;
	assign _1204_ = _1937_ | ~_4317_;
	assign _1205_ = \mchip.pong.game.ball.dpath.ballY [0] | ~\mchip.pong.game.vga.line_ind [0];
	assign _1206_ = _4317_ ^ _1937_;
	assign _1207_ = _1205_ & ~_1206_;
	assign _1209_ = _1204_ & ~_1207_;
	assign _1210_ = _1203_ & ~_1209_;
	assign _1211_ = _1201_ & ~_1210_;
	assign _1212_ = _1196_ & ~_1211_;
	assign _1213_ = _1193_ & ~_1212_;
	assign _1214_ = _1179_ & ~_1213_;
	assign _1215_ = _1622_ | ~_4230_;
	assign _1216_ = _1600_ & ~_1215_;
	assign _1217_ = _1216_ | _1214_;
	assign _1218_ = \mchip.pong.game.ball.dpath.ballY [0] ^ \mchip.pong.game.vga.line_ind [0];
	assign _1220_ = ~(_1218_ | _1206_);
	assign _1221_ = _1220_ & _1203_;
	assign _1222_ = ~(_1221_ & _1196_);
	assign _1223_ = _1179_ & ~_1222_;
	assign _1224_ = _1217_ & ~_1223_;
	assign _1225_ = _4230_ ^ _1611_;
	assign _1226_ = _4406_ & _4402_;
	assign _1227_ = _4216_ ^ _2877_;
	assign _1228_ = _4217_ ^ \mchip.pong.game.ball.dpath.ballY [6];
	assign _1229_ = _1228_ | ~_1227_;
	assign _1231_ = _1226_ & ~_1229_;
	assign _1232_ = _4370_ | _4374_;
	assign _1233_ = ~(_1232_ | _4397_);
	assign _1234_ = _1233_ & _1231_;
	assign _1235_ = ~(_1234_ & _1225_);
	assign _1236_ = _4230_ | _1611_;
	assign _1237_ = _4216_ | _2877_;
	assign _1238_ = _4217_ | _1739_;
	assign _1239_ = _1227_ & ~_1238_;
	assign _1240_ = _1237_ & ~_1239_;
	assign _1242_ = _4220_ | _2658_;
	assign _1243_ = _4406_ & _4401_;
	assign _1244_ = _1242_ & ~_1243_;
	assign _1245_ = ~(_1244_ | _1229_);
	assign _1246_ = _1240_ & ~_1245_;
	assign _1247_ = _4319_ | _4393_;
	assign _1248_ = \mchip.pong.game.ball.dpath.ballY [2] & ~_4318_;
	assign _1249_ = _1248_ & ~_4385_;
	assign _1250_ = _1247_ & ~_1249_;
	assign _1251_ = _4317_ | _3073_;
	assign _1253_ = _4373_ & ~_4370_;
	assign _1254_ = _1253_ | ~_1251_;
	assign _1255_ = _1254_ & ~_4397_;
	assign _1256_ = _1250_ & ~_1255_;
	assign _1257_ = _1231_ & ~_1256_;
	assign _1258_ = _1246_ & ~_1257_;
	assign _1259_ = _1225_ & ~_1258_;
	assign _1260_ = _1236_ & ~_1259_;
	assign _1261_ = _1235_ & ~_1260_;
	assign _1262_ = _1261_ | _1224_;
	assign _1263_ = _1262_ | _1176_;
	assign _1264_ = ~(_1263_ | _1138_);
	assign _1265_ = _4230_ | _3899_;
	assign _1266_ = _4220_ ^ _3742_;
	assign _1267_ = _4221_ ^ \mchip.pong.game.left_paddle.coord [4];
	assign _1268_ = _1266_ & ~_1267_;
	assign _1269_ = _4217_ ^ \mchip.pong.game.left_paddle.coord [6];
	assign _1270_ = _4216_ ^ \mchip.pong.game.left_paddle.coord [7];
	assign _1271_ = _1270_ | _1269_;
	assign _1272_ = _1268_ & ~_1271_;
	assign _1273_ = _4319_ | _3786_;
	assign _1274_ = \mchip.pong.game.left_paddle.coord [2] & ~_4318_;
	assign _1275_ = _4319_ ^ \mchip.pong.game.left_paddle.coord [3];
	assign _1276_ = _1274_ & ~_1275_;
	assign _1277_ = _1273_ & ~_1276_;
	assign _1278_ = _4318_ ^ \mchip.pong.game.left_paddle.coord [2];
	assign _1279_ = ~(_1278_ | _1275_);
	assign _1280_ = _4317_ | _3830_;
	assign _1281_ = \mchip.pong.game.vga.line_ind [0] | \mchip.pong.game.left_paddle.coord [0];
	assign _1282_ = _4317_ ^ \mchip.pong.game.left_paddle.coord [1];
	assign _1284_ = _1281_ & ~_1282_;
	assign _1285_ = _1280_ & ~_1284_;
	assign _1286_ = _1279_ & ~_1285_;
	assign _1287_ = _1277_ & ~_1286_;
	assign _1288_ = _1272_ & ~_1287_;
	assign _1289_ = \mchip.pong.game.left_paddle.coord [7] & ~_4216_;
	assign _1290_ = \mchip.pong.game.left_paddle.coord [6] & ~_4217_;
	assign _1291_ = _1290_ & ~_1270_;
	assign _1292_ = _1291_ | _1289_;
	assign _1293_ = _4220_ | _3742_;
	assign _1295_ = _4221_ | _3720_;
	assign _1296_ = _1266_ & ~_1295_;
	assign _1297_ = _1293_ & ~_1296_;
	assign _1298_ = ~(_1297_ | _1271_);
	assign _1299_ = _1298_ | _1292_;
	assign _1300_ = ~(_1299_ | _1288_);
	assign _1301_ = _4230_ ^ _3899_;
	assign _1302_ = _1301_ & ~_1300_;
	assign _1303_ = _1265_ & ~_1302_;
	assign _1304_ = ~(\mchip.pong.game.vga.line_ind [0] ^ \mchip.pong.game.left_paddle.coord [0]);
	assign _1306_ = ~(_1304_ | _1282_);
	assign _1307_ = _1306_ & _1279_;
	assign _1308_ = ~(_1307_ & _1272_);
	assign _1309_ = _1301_ & ~_1308_;
	assign _1310_ = _1309_ | _1303_;
	assign _1311_ = _4230_ ^ _4003_;
	assign _1312_ = _4002_ & ~_1311_;
	assign _1313_ = ~_4216_;
	assign _1314_ = _1313_ | _4035_;
	assign _1315_ = _4216_ ^ _4009_;
	assign _1317_ = ~_4217_;
	assign _1318_ = _1317_ | _4011_;
	assign _1319_ = _1315_ & ~_1318_;
	assign _1320_ = _1314_ & ~_1319_;
	assign _1321_ = _4217_ ^ _4011_;
	assign _1322_ = _1321_ | ~_1315_;
	assign _1323_ = ~_4220_;
	assign _1324_ = _1323_ | _4017_;
	assign _1325_ = _4221_ & ~_4014_;
	assign _1326_ = _4220_ ^ _4017_;
	assign _1328_ = _1325_ & ~_1326_;
	assign _1329_ = _1328_ | ~_1324_;
	assign _1330_ = _1329_ & ~_1322_;
	assign _1331_ = _1320_ & ~_1330_;
	assign _1332_ = _4319_ ^ _4022_;
	assign _1333_ = _4318_ ^ _4024_;
	assign _1334_ = _1332_ & ~_1333_;
	assign _1335_ = _4027_ | ~_4317_;
	assign _1336_ = \mchip.pong.game.left_paddle.coord [0] | ~\mchip.pong.game.vga.line_ind [0];
	assign _1337_ = _4317_ ^ _4027_;
	assign _1339_ = _1336_ & ~_1337_;
	assign _1340_ = _1335_ & ~_1339_;
	assign _1341_ = _1334_ & ~_1340_;
	assign _1342_ = _4022_ & ~_4205_;
	assign _1343_ = _4206_ | _4024_;
	assign _1344_ = _1332_ & ~_1343_;
	assign _1345_ = _1344_ | _1342_;
	assign _1346_ = _1345_ | _1341_;
	assign _1347_ = _4221_ ^ _4014_;
	assign _1348_ = _1347_ | _1326_;
	assign _1350_ = _1348_ | _1322_;
	assign _1351_ = _1346_ & ~_1350_;
	assign _1352_ = _1331_ & ~_1351_;
	assign _1353_ = _1312_ & ~_1352_;
	assign _1354_ = _4003_ | ~_4230_;
	assign _1355_ = _4002_ & ~_1354_;
	assign _1356_ = _1355_ | _1353_;
	assign _1357_ = _1304_ & ~_1337_;
	assign _1358_ = ~(_1357_ & _1334_);
	assign _1359_ = _1358_ | _1350_;
	assign _1361_ = _1312_ & ~_1359_;
	assign _1362_ = _1356_ & ~_1361_;
	assign _1363_ = _1310_ & ~_1362_;
	assign _1364_ = _4239_ | _4237_;
	assign _1365_ = _4157_ & _4101_;
	assign _1366_ = _4244_ | _4243_;
	assign _1367_ = _4234_ & ~_1366_;
	assign _1368_ = ~(_1367_ & _1365_);
	assign _1369_ = _1368_ | _1364_;
	assign _1370_ = _1366_ | _4234_;
	assign _1372_ = _4101_ & ~_4157_;
	assign _1373_ = _1367_ & ~_1372_;
	assign _1374_ = _1370_ & ~_1373_;
	assign _1375_ = _1374_ | _1364_;
	assign _1376_ = _1369_ & ~_1375_;
	assign _1377_ = _1363_ & ~_1376_;
	assign _1378_ = _4102_ & ~_4158_;
	assign _1379_ = _4245_ & _4099_;
	assign _1380_ = ~(_1379_ & _1378_);
	assign _1381_ = _1380_ | _1364_;
	assign _1383_ = _4245_ & ~_1364_;
	assign _1384_ = _4158_ | ~_4099_;
	assign _1385_ = _1383_ & ~_1384_;
	assign _1386_ = ~(_1366_ | _1364_);
	assign _1387_ = _1386_ | _1385_;
	assign _1388_ = _1381_ & ~_1387_;
	assign _1389_ = _1377_ & ~_1388_;
	assign _1390_ = _4230_ ^ _2013_;
	assign _1391_ = ~(_4216_ & _1783_);
	assign _1392_ = _4216_ ^ _1783_;
	assign _1394_ = ~(_4217_ & _1728_);
	assign _1395_ = _1392_ & ~_1394_;
	assign _1396_ = _1391_ & ~_1395_;
	assign _1397_ = _4217_ ^ \mchip.pong.game.right_paddle.coord [6];
	assign _1398_ = _1392_ & ~_1397_;
	assign _1399_ = ~(_4220_ & _1654_);
	assign _1400_ = _4220_ ^ _1654_;
	assign _1401_ = ~(_4221_ & _2111_);
	assign _1402_ = _1400_ & ~_1401_;
	assign _1403_ = _1399_ & ~_1402_;
	assign _1405_ = _1398_ & ~_1403_;
	assign _1406_ = _1396_ & ~_1405_;
	assign _1407_ = _4221_ ^ _2111_;
	assign _1408_ = ~(_1407_ & _1400_);
	assign _1409_ = _1398_ & ~_1408_;
	assign _1410_ = _4205_ | \mchip.pong.game.right_paddle.coord [3];
	assign _1411_ = _4319_ ^ _1849_;
	assign _1412_ = _4206_ | \mchip.pong.game.right_paddle.coord [2];
	assign _1413_ = _1411_ & ~_1412_;
	assign _1414_ = _1410_ & ~_1413_;
	assign _1416_ = _4318_ ^ \mchip.pong.game.right_paddle.coord [2];
	assign _1417_ = _1411_ & ~_1416_;
	assign _1418_ = ~(_4317_ & _1926_);
	assign _1419_ = ~(\mchip.pong.game.vga.line_ind [0] & \mchip.pong.game.right_paddle.coord [0]);
	assign _1420_ = _4317_ ^ \mchip.pong.game.right_paddle.coord [1];
	assign _1421_ = _1419_ & ~_1420_;
	assign _1422_ = _1418_ & ~_1421_;
	assign _1423_ = _1417_ & ~_1422_;
	assign _1424_ = _1414_ & ~_1423_;
	assign _1425_ = _1409_ & ~_1424_;
	assign _1427_ = _1406_ & ~_1425_;
	assign _1428_ = _1390_ & ~_1427_;
	assign _1429_ = _4230_ & ~\mchip.pong.game.right_paddle.coord [8];
	assign _1430_ = _1429_ | _1428_;
	assign _1431_ = ~(\mchip.pong.game.vga.line_ind [0] ^ \mchip.pong.game.right_paddle.coord [0]);
	assign _1432_ = ~(_1431_ | _1420_);
	assign _1433_ = _1432_ & _1417_;
	assign _1434_ = ~(_1433_ & _1409_);
	assign _1435_ = _1390_ & ~_1434_;
	assign _1436_ = _1435_ | _1430_;
	assign _1438_ = _4230_ ^ _2504_;
	assign _1439_ = _2493_ & ~_1438_;
	assign _1440_ = _1313_ | _2888_;
	assign _1441_ = _4216_ ^ _2570_;
	assign _1442_ = _1317_ | _2592_;
	assign _1443_ = _1441_ & ~_1442_;
	assign _1444_ = _1440_ & ~_1443_;
	assign _1445_ = _4217_ ^ _2592_;
	assign _1446_ = _1445_ | ~_1441_;
	assign _1447_ = _1323_ | _2680_;
	assign _1449_ = _4221_ & ~_2636_;
	assign _1450_ = _4220_ ^ _2680_;
	assign _1451_ = _1449_ & ~_1450_;
	assign _1452_ = _1451_ | ~_1447_;
	assign _1453_ = _1452_ & ~_1446_;
	assign _1454_ = _1444_ & ~_1453_;
	assign _1455_ = _4319_ ^ _2734_;
	assign _1456_ = _4318_ ^ _2756_;
	assign _1457_ = _1455_ & ~_1456_;
	assign _1458_ = _2789_ | ~_4317_;
	assign _1460_ = \mchip.pong.game.right_paddle.coord [0] | ~\mchip.pong.game.vga.line_ind [0];
	assign _1461_ = _4317_ ^ _2789_;
	assign _1462_ = _1460_ & ~_1461_;
	assign _1463_ = _1458_ & ~_1462_;
	assign _1464_ = _1457_ & ~_1463_;
	assign _1465_ = _2734_ & ~_4205_;
	assign _1466_ = _4206_ | _2756_;
	assign _1467_ = _1455_ & ~_1466_;
	assign _1468_ = _1467_ | _1465_;
	assign _1469_ = _1468_ | _1464_;
	assign _1471_ = _4221_ ^ _2636_;
	assign _1472_ = _1471_ | _1450_;
	assign _1473_ = _1472_ | _1446_;
	assign _1474_ = _1469_ & ~_1473_;
	assign _1475_ = _1454_ & ~_1474_;
	assign _1476_ = _1439_ & ~_1475_;
	assign _1477_ = _2504_ | ~_4230_;
	assign _1478_ = _2493_ & ~_1477_;
	assign _1479_ = _1478_ | _1476_;
	assign _1480_ = \mchip.pong.game.vga.line_ind [0] ^ \mchip.pong.game.right_paddle.coord [0];
	assign _1482_ = ~(_1480_ | _1461_);
	assign _1483_ = ~(_1482_ & _1457_);
	assign _1484_ = _1483_ | _1473_;
	assign _1485_ = _1439_ & ~_1484_;
	assign _1486_ = _1479_ & ~_1485_;
	assign _1487_ = _1436_ & ~_1486_;
	assign _1488_ = \mchip.pong.game.vga.pix_ind [1] | ~\mchip.pong.game.vga.pix_ind [0];
	assign _1489_ = ~(_1488_ | _4158_);
	assign _1490_ = _1489_ & _1379_;
	assign _1491_ = ~(_1490_ & _4240_);
	assign _1493_ = _4245_ & ~_4099_;
	assign _1494_ = _1080_ & ~_1493_;
	assign _1495_ = _4157_ & ~_4158_;
	assign _1496_ = _1379_ & ~_1495_;
	assign _1497_ = _1494_ & ~_1496_;
	assign _1498_ = _4240_ & ~_1497_;
	assign _1499_ = _4239_ & _4237_;
	assign _1500_ = _1499_ | _1498_;
	assign _1501_ = _1491_ & ~_1500_;
	assign _1502_ = _1487_ & ~_1501_;
	assign _1504_ = \mchip.pong.game.vga.pix_ind [3] & ~\mchip.pong.game.vga.pix_ind [2];
	assign _1505_ = _1504_ & _4157_;
	assign _1506_ = _1505_ & _1379_;
	assign _1507_ = ~(_1506_ & _4240_);
	assign _1508_ = _1080_ & ~_4237_;
	assign _1509_ = _4244_ & ~_4365_;
	assign _1510_ = _4365_ & _4244_;
	assign _1511_ = \mchip.pong.game.vga.pix_ind [4] & ~\mchip.pong.game.vga.pix_ind [3];
	assign _1512_ = _1510_ & ~_1511_;
	assign _1513_ = _1512_ | _1509_;
	assign _1515_ = _1508_ & ~_1513_;
	assign _1516_ = _1515_ | _1070_;
	assign _1517_ = _1507_ & ~_1516_;
	assign _1518_ = _1502_ & ~_1517_;
	assign _1519_ = _1518_ | _1389_;
	assign \mchip.pong.VGA_G2  = (_1264_ ? _1062_ : _1519_);
	assign _1520_ = _0056_ & ~_0726_;
	assign _1521_ = (_0159_ ? _0351_ : _1520_);
	assign _1522_ = _0114_ & _4423_;
	assign _1524_ = ~(_0114_ | _4423_);
	assign _1525_ = _1524_ | _1522_;
	assign _1526_ = _0056_ & ~_1525_;
	assign _1527_ = (_4387_ ? _0107_ : _0118_);
	assign _1528_ = _0127_ & ~_1527_;
	assign _1529_ = (_0146_ ? _1526_ : _1528_);
	assign _1530_ = (\mchip.pong.game.vga.pix_ind [0] ? _1529_ : _1521_);
	assign _1531_ = _0193_ & ~_0127_;
	assign _1532_ = _4389_ & ~_4387_;
	assign _1533_ = _0127_ & ~_1532_;
	assign _1535_ = (_0146_ ? _1531_ : _1533_);
	assign _1536_ = _0056_ & ~_0783_;
	assign _1537_ = _0127_ & ~_1522_;
	assign _1538_ = (_0146_ ? _1536_ : _1537_);
	assign _1539_ = (\mchip.pong.game.vga.pix_ind [0] ? _1538_ : _1535_);
	assign _1540_ = (_1103_ ? _1530_ : _1539_);
	assign _1541_ = _0237_ | _0056_;
	assign _1542_ = _0410_ | _4423_;
	assign _1543_ = _1542_ | _0127_;
	assign _1544_ = (_0146_ ? _1541_ : _1543_);
	assign _1546_ = _1544_ & ~\mchip.pong.game.vga.pix_ind [0];
	assign _1547_ = _0127_ & ~_0197_;
	assign _1548_ = ~(_4387_ & _0090_);
	assign _1549_ = _0056_ & ~_1548_;
	assign _1550_ = (_0146_ ? _1547_ : _1549_);
	assign _1551_ = \mchip.pong.game.vga.pix_ind [0] & ~_1550_;
	assign _1552_ = ~(_1551_ | _1546_);
	assign _1553_ = _4443_ & _4423_;
	assign _1554_ = (_0127_ ? _1553_ : _0500_);
	assign _1555_ = _0035_ & ~_4423_;
	assign _1557_ = _4423_ & ~_0119_;
	assign _1558_ = (_0056_ ? _1555_ : _1557_);
	assign _1559_ = (_0146_ ? _1554_ : _1558_);
	assign _1560_ = ~(_4423_ | _4389_);
	assign _1561_ = (_0056_ ? _1560_ : _1557_);
	assign _1562_ = _4423_ & _4389_;
	assign _1563_ = (_0127_ ? _1562_ : _0500_);
	assign _1564_ = (_0146_ ? _1561_ : _1563_);
	assign _1565_ = (\mchip.pong.game.vga.pix_ind [0] ? _1564_ : _1559_);
	assign _1566_ = (_1103_ ? _1552_ : _1565_);
	assign _1568_ = (_0044_ ? _1540_ : _1566_);
	assign _1569_ = (_4387_ ? _0107_ : _0114_);
	assign _1570_ = _0127_ & ~_1569_;
	assign _1571_ = (_4387_ ? _0119_ : _0131_);
	assign _1572_ = _0056_ & ~_1571_;
	assign _1573_ = (_0146_ ? _1570_ : _1572_);
	assign _1574_ = _4387_ | ~_0035_;
	assign _1575_ = _0127_ & ~_1574_;
	assign _1576_ = _0056_ & ~_0766_;
	assign _1577_ = (_0146_ ? _1575_ : _1576_);
	assign _1579_ = (\mchip.pong.game.vga.pix_ind [0] ? _1577_ : _1573_);
	assign _1580_ = _0127_ & ~_0134_;
	assign _1581_ = (_0159_ ? _0111_ : _1580_);
	assign _1582_ = _0410_ | _4387_;
	assign _1583_ = _0127_ & ~_1582_;
	assign _1584_ = (_0146_ ? _1583_ : _0096_);
	assign _1585_ = (\mchip.pong.game.vga.pix_ind [0] ? _1584_ : _1581_);
	assign _1586_ = (_1103_ ? _1579_ : _1585_);
	assign _1587_ = (\mchip.pong.game.vga.pix_ind [0] ? _0130_ : _0168_);
	assign _1588_ = _0056_ & ~_0330_;
	assign _1590_ = _0127_ & ~_0766_;
	assign _1591_ = (_0159_ ? _1588_ : _1590_);
	assign _1592_ = _0056_ & ~_1569_;
	assign _1593_ = (_0146_ ? _0335_ : _1592_);
	assign _1594_ = (\mchip.pong.game.vga.pix_ind [0] ? _1593_ : _1591_);
	assign _1595_ = (_1103_ ? _1587_ : _1594_);
	assign _1596_ = (_0044_ ? _1586_ : _1595_);
	assign _1597_ = (_0088_ ? _1568_ : _1596_);
	assign _1598_ = (_1103_ ? _0233_ : _0248_);
	assign _1599_ = ~(_0160_ & _0056_);
	assign _1601_ = _0162_ | _0056_;
	assign _1602_ = (_0159_ ? _1599_ : _1601_);
	assign _1603_ = (_0146_ ? _1601_ : _0192_);
	assign _1604_ = (\mchip.pong.game.vga.pix_ind [0] ? _1602_ : _1603_);
	assign _1605_ = _1604_ | _1103_;
	assign _1606_ = _0218_ | _0063_;
	assign _1607_ = ~(_1606_ & _1605_);
	assign _1608_ = (_0044_ ? _1598_ : _1607_);
	assign _1609_ = _0173_ | _0127_;
	assign _1610_ = (_0146_ ? _0200_ : _1609_);
	assign _1612_ = ~(_0361_ & _4387_);
	assign _1613_ = _1612_ | _0056_;
	assign _1614_ = (_0146_ ? _1613_ : _1609_);
	assign _1615_ = (\mchip.pong.game.vga.pix_ind [0] ? _1614_ : _1610_);
	assign _1616_ = (_1103_ ? _1615_ : _0191_);
	assign _1617_ = _0044_ & ~_1616_;
	assign _1618_ = _0228_ & ~_0044_;
	assign _1619_ = _1618_ | _1617_;
	assign _1620_ = (_0088_ ? _1608_ : _1619_);
	assign _1621_ = (_4368_ ? _1597_ : _1620_);
	assign _1623_ = (\mchip.pong.game.vga.pix_ind [0] ? _0191_ : _0218_);
	assign _1624_ = (_1103_ ? _0218_ : _1623_);
	assign _1625_ = _0308_ & ~_1624_;
	assign _1626_ = (\mchip.pong.game.vga.pix_ind [0] ? _1610_ : _1614_);
	assign _1627_ = (_1103_ ? _1626_ : _1610_);
	assign _1628_ = _0044_ & ~_1627_;
	assign _1629_ = _1628_ | _1625_;
	assign _1630_ = ~(_0872_ | _0127_);
	assign _1631_ = (_0146_ ? _0163_ : _1630_);
	assign _1632_ = (\mchip.pong.game.vga.pix_ind [0] ? _1631_ : _0164_);
	assign _1634_ = (_1103_ ? _0165_ : _1632_);
	assign _1635_ = _0056_ & ~_1574_;
	assign _1636_ = (_0146_ ? _0129_ : _1635_);
	assign _1637_ = _0127_ & ~_0110_;
	assign _1638_ = (_0146_ ? _1637_ : _0135_);
	assign _1639_ = (\mchip.pong.game.vga.pix_ind [0] ? _1638_ : _1636_);
	assign _1640_ = (_1103_ ? _1639_ : _0169_);
	assign _1641_ = (_0044_ ? _1634_ : _1640_);
	assign _1642_ = (_0088_ ? _1629_ : _1641_);
	assign _1644_ = (_4423_ ? _0117_ : _0792_);
	assign _1645_ = _0056_ & ~_1644_;
	assign _1646_ = (_4387_ ? _0113_ : _0118_);
	assign _1647_ = _0127_ & ~_1646_;
	assign _1648_ = (_0146_ ? _1645_ : _1647_);
	assign _1649_ = ~(_0451_ & _4387_);
	assign _1650_ = _0056_ & ~_1649_;
	assign _1651_ = ~(_0421_ & _4423_);
	assign _1652_ = _0127_ & ~_1651_;
	assign _1653_ = (_0146_ ? _1650_ : _1652_);
	assign _1655_ = (\mchip.pong.game.vga.pix_ind [0] ? _1653_ : _1648_);
	assign _1656_ = (_0127_ ? _4418_ : _0484_);
	assign _1657_ = (_0127_ ? _1532_ : _1524_);
	assign _1658_ = (_0146_ ? _1656_ : _1657_);
	assign _1659_ = _4443_ & ~_4387_;
	assign _1660_ = (_0127_ ? _1659_ : _1524_);
	assign _1661_ = (_0056_ ? _1555_ : _0270_);
	assign _1662_ = (_0146_ ? _1660_ : _1661_);
	assign _1663_ = (\mchip.pong.game.vga.pix_ind [0] ? _1662_ : _1658_);
	assign _1664_ = (_1103_ ? _1655_ : _1663_);
	assign _1666_ = (_0159_ ? _0194_ : _0198_);
	assign _1667_ = \mchip.pong.game.vga.pix_ind [0] & ~_1666_;
	assign _1668_ = _4423_ & ~_4428_;
	assign _1669_ = _0127_ & ~_1668_;
	assign _1670_ = (_0146_ ? _1536_ : _1669_);
	assign _1671_ = (\mchip.pong.game.vga.pix_ind [0] ? _1535_ : _1670_);
	assign _1672_ = (_1103_ ? _1667_ : _1671_);
	assign _1673_ = (_0044_ ? _1664_ : _1672_);
	assign _1674_ = (_0056_ ? _4429_ : _1532_);
	assign _1676_ = _0056_ & ~_0193_;
	assign _1677_ = (_0146_ ? _1674_ : _1676_);
	assign _1678_ = _0127_ & ~_0237_;
	assign _1679_ = _0255_ | _4423_;
	assign _1680_ = _0056_ & ~_1679_;
	assign _1681_ = (_0146_ ? _1678_ : _1680_);
	assign _1682_ = (\mchip.pong.game.vga.pix_ind [0] ? _1681_ : _1677_);
	assign _1683_ = _0102_ | _4387_;
	assign _1684_ = _0127_ & ~_1683_;
	assign _1685_ = _0056_ & ~_0402_;
	assign _1687_ = (_0146_ ? _1684_ : _1685_);
	assign _1688_ = _0056_ & ~_0288_;
	assign _1689_ = (_0146_ ? _0321_ : _1688_);
	assign _1690_ = (\mchip.pong.game.vga.pix_ind [0] ? _1689_ : _1687_);
	assign _1691_ = (_1103_ ? _1682_ : _1690_);
	assign _1692_ = _0056_ & ~_0128_;
	assign _1693_ = (_0146_ ? _0324_ : _1692_);
	assign _1694_ = (_0146_ ? _0331_ : _1572_);
	assign _1695_ = (\mchip.pong.game.vga.pix_ind [0] ? _1694_ : _1693_);
	assign _1696_ = _0056_ & ~_0334_;
	assign _1698_ = (_0146_ ? _0335_ : _1696_);
	assign _1699_ = _0127_ & ~_1571_;
	assign _1700_ = (_0146_ ? _1699_ : _1588_);
	assign _1701_ = (\mchip.pong.game.vga.pix_ind [0] ? _1700_ : _1698_);
	assign _1702_ = (_1103_ ? _1695_ : _1701_);
	assign _1703_ = (_0044_ ? _1702_ : _1691_);
	assign _1704_ = (_0088_ ? _1703_ : _1673_);
	assign _1705_ = (_4368_ ? _1642_ : _1704_);
	assign _1706_ = (_4367_ ? _1621_ : _1705_);
	assign _1708_ = _1592_ | _0167_;
	assign _1709_ = (_4423_ ? _0054_ : _4428_);
	assign _1710_ = (_0127_ ? _0793_ : _1709_);
	assign _1711_ = (_0146_ ? _1708_ : _1710_);
	assign _1712_ = _4423_ & ~_0880_;
	assign _1713_ = (_0127_ ? _0356_ : _1712_);
	assign _1714_ = (_4387_ ? _0792_ : _0035_);
	assign _1715_ = (_0127_ ? _0793_ : _1714_);
	assign _1716_ = (_0146_ ? _1713_ : _1715_);
	assign _1717_ = (\mchip.pong.game.vga.pix_ind [0] ? _1716_ : _1711_);
	assign _1719_ = ~_0320_;
	assign _1720_ = ~_0766_;
	assign _1721_ = (_0056_ ? _1719_ : _1720_);
	assign _1722_ = (_4423_ ? _0421_ : _0522_);
	assign _1723_ = (_4423_ ? _0035_ : _0401_);
	assign _1724_ = (_0127_ ? _1722_ : _1723_);
	assign _1725_ = (_0146_ ? _1721_ : _1724_);
	assign _1726_ = (_0056_ ? _0051_ : _0334_);
	assign _1727_ = ~_1726_;
	assign _1729_ = ~_1569_;
	assign _1730_ = (_4387_ ? _4428_ : _0451_);
	assign _1731_ = (_0056_ ? _1729_ : _1730_);
	assign _1732_ = (_0146_ ? _1727_ : _1731_);
	assign _1733_ = (\mchip.pong.game.vga.pix_ind [0] ? _1732_ : _1725_);
	assign _1734_ = (_1103_ ? _1717_ : _1733_);
	assign _1735_ = (_0044_ ? _1586_ : _1734_);
	assign _1736_ = (_0088_ ? _1568_ : _1735_);
	assign _1737_ = ~_0783_;
	assign _1738_ = ~_0162_;
	assign _1740_ = (_0056_ ? _1737_ : _1738_);
	assign _1741_ = (_4389_ ? _4371_ : _4375_);
	assign _1742_ = (_4423_ ? _0153_ : _1741_);
	assign _1743_ = _1742_ | _0127_;
	assign _1744_ = (_0146_ ? _1740_ : _1743_);
	assign _1745_ = _4423_ | ~_0207_;
	assign _1746_ = (_0127_ ? _0154_ : _1745_);
	assign _1747_ = _4387_ & ~_0410_;
	assign _1748_ = ~_1747_;
	assign _1749_ = (_4387_ ? _4371_ : _4381_);
	assign _1751_ = (_0127_ ? _1748_ : _1749_);
	assign _1752_ = (_0146_ ? _1746_ : _1751_);
	assign _1753_ = (\mchip.pong.game.vga.pix_ind [0] ? _1752_ : _1744_);
	assign _1754_ = (_4387_ ? _0118_ : _0852_);
	assign _1755_ = (_0127_ ? _0154_ : _1754_);
	assign _1756_ = _1548_ & _0098_;
	assign _1757_ = ~_1756_;
	assign _1758_ = (_0127_ ? _4423_ : _1757_);
	assign _1759_ = (_0146_ ? _1755_ : _1758_);
	assign _1760_ = (_4387_ ? _0118_ : _0442_);
	assign _1762_ = (_0127_ ? _0399_ : _1760_);
	assign _1763_ = (_4423_ ? _0665_ : _0792_);
	assign _1764_ = (_4387_ ? _0970_ : _0054_);
	assign _1765_ = (_0127_ ? _1763_ : _1764_);
	assign _1766_ = (_0146_ ? _1762_ : _1765_);
	assign _1767_ = (\mchip.pong.game.vga.pix_ind [0] ? _1766_ : _1759_);
	assign _1768_ = (_1103_ ? _1753_ : _1767_);
	assign _1769_ = (_4423_ ? _0114_ : _0472_);
	assign _1770_ = _0127_ & ~_1769_;
	assign _1771_ = ~_1770_;
	assign _1773_ = (_4423_ ? _4409_ : _0101_);
	assign _1774_ = _1773_ | _0127_;
	assign _1775_ = (_0146_ ? _1771_ : _1774_);
	assign _1776_ = _0472_ & ~_4423_;
	assign _1777_ = _0127_ & ~_1776_;
	assign _1778_ = ~_1777_;
	assign _1779_ = (_0146_ ? _1778_ : _1774_);
	assign _1780_ = (\mchip.pong.game.vga.pix_ind [0] ? _1779_ : _1775_);
	assign _1781_ = (_4389_ ? _4374_ : _4372_);
	assign _1782_ = ~_1781_;
	assign _1784_ = ~(_1782_ | _4423_);
	assign _1785_ = (_0056_ ? _0480_ : _1784_);
	assign _1786_ = (_4423_ ? _4409_ : _0656_);
	assign _1787_ = _1786_ | _0127_;
	assign _1788_ = (_0146_ ? _1785_ : _1787_);
	assign _1789_ = (_0127_ ? _0048_ : _0726_);
	assign _1790_ = (_4389_ ? _4408_ : _4374_);
	assign _1791_ = (_4423_ ? _0153_ : _1790_);
	assign _1792_ = _1791_ | _0127_;
	assign _1793_ = (_0146_ ? _1789_ : _1792_);
	assign _1795_ = (\mchip.pong.game.vga.pix_ind [0] ? _1793_ : _1788_);
	assign _1796_ = (_1103_ ? _1780_ : _1795_);
	assign _1797_ = (_0044_ ? _1768_ : _1796_);
	assign _1798_ = ~_0154_;
	assign _1799_ = _1024_ | _4387_;
	assign _1800_ = (_0127_ ? _1798_ : _1799_);
	assign _1801_ = (_4423_ ? _0435_ : _0101_);
	assign _1802_ = (_0127_ ? _0755_ : _1801_);
	assign _1803_ = (_0146_ ? _1800_ : _1802_);
	assign _1804_ = (_4389_ ? _4372_ : _0582_);
	assign _1806_ = _4387_ & ~_1804_;
	assign _1807_ = ~_1806_;
	assign _1808_ = (_4389_ ? _4424_ : _4375_);
	assign _1809_ = ~_1808_;
	assign _1810_ = (_4387_ ? _0451_ : _1809_);
	assign _1811_ = (_0127_ ? _1807_ : _1810_);
	assign _1812_ = (_4423_ ? _4443_ : _0101_);
	assign _1813_ = _1812_ | _0127_;
	assign _1814_ = (_0146_ ? _1811_ : _1813_);
	assign _1815_ = (\mchip.pong.game.vga.pix_ind [0] ? _1814_ : _1803_);
	assign _1817_ = _4423_ & ~_0421_;
	assign _1818_ = ~_1817_;
	assign _1819_ = (_0127_ ? _0619_ : _1818_);
	assign _1820_ = (_4423_ ? _4434_ : _0101_);
	assign _1821_ = _1820_ | _0127_;
	assign _1822_ = (_0146_ ? _1819_ : _1821_);
	assign _1823_ = _0618_ & ~_0056_;
	assign _1824_ = ~_1823_;
	assign _1825_ = (_0146_ ? _1824_ : _1821_);
	assign _1826_ = (\mchip.pong.game.vga.pix_ind [0] ? _1825_ : _1822_);
	assign _1828_ = (_1103_ ? _1815_ : _1826_);
	assign _1829_ = (_4387_ ? _0495_ : _0254_);
	assign _1830_ = (_4423_ ? _0093_ : _0475_);
	assign _1831_ = (_0127_ ? _1829_ : _1830_);
	assign _1832_ = (_4389_ ? _4375_ : _4372_);
	assign _1833_ = (_4423_ ? _1832_ : _0474_);
	assign _1834_ = _0056_ & ~_1833_;
	assign _1835_ = _1834_ | _0681_;
	assign _1836_ = (_0146_ ? _1831_ : _1835_);
	assign _1837_ = (_4423_ ? _0454_ : _0206_);
	assign _1839_ = ~_1837_;
	assign _1840_ = (_0127_ ? _1829_ : _1839_);
	assign _1841_ = _4387_ & ~_0628_;
	assign _1842_ = _0127_ & ~_1841_;
	assign _1843_ = _1842_ | _1834_;
	assign _1844_ = (_0146_ ? _1840_ : _1843_);
	assign _1845_ = (\mchip.pong.game.vga.pix_ind [0] ? _1844_ : _1836_);
	assign _1846_ = _0366_ | _0100_;
	assign _1847_ = (_4387_ ? _0451_ : _1846_);
	assign _1848_ = (_0127_ ? _1798_ : _1847_);
	assign _1850_ = _4387_ & ~_0656_;
	assign _1851_ = ~_1850_;
	assign _1852_ = (_4389_ ? _4375_ : _4407_);
	assign _1853_ = ~_1852_;
	assign _1854_ = (_4423_ ? _0435_ : _1853_);
	assign _1855_ = (_0127_ ? _1851_ : _1854_);
	assign _1856_ = (_0146_ ? _1848_ : _1855_);
	assign _1857_ = (_4423_ ? _1024_ : _0451_);
	assign _1858_ = (_0127_ ? _1798_ : _1857_);
	assign _1859_ = (_4389_ ? _0065_ : _4408_);
	assign _1861_ = (_4423_ ? _0435_ : _1859_);
	assign _1862_ = (_0127_ ? _0592_ : _1861_);
	assign _1863_ = (_0146_ ? _1858_ : _1862_);
	assign _1864_ = (\mchip.pong.game.vga.pix_ind [0] ? _1863_ : _1856_);
	assign _1865_ = (_1103_ ? _1845_ : _1864_);
	assign _1866_ = (_0044_ ? _1828_ : _1865_);
	assign _1867_ = (_0088_ ? _1797_ : _1866_);
	assign _1868_ = (_4368_ ? _1736_ : _1867_);
	assign _1869_ = (_4423_ ? _0101_ : _1804_);
	assign _1870_ = (_4389_ ? _4371_ : _0425_);
	assign _1872_ = (_4423_ ? _0117_ : _1870_);
	assign _1873_ = (_0127_ ? _1869_ : _1872_);
	assign _1874_ = (_4387_ ? _0475_ : _1853_);
	assign _1875_ = _1874_ | _0127_;
	assign _1876_ = (_0146_ ? _1873_ : _1875_);
	assign _1877_ = (_4423_ ? _0665_ : _0153_);
	assign _1878_ = ~_1877_;
	assign _1879_ = (_4423_ ? _0117_ : _0207_);
	assign _1880_ = (_0127_ ? _1878_ : _1879_);
	assign _1881_ = (_4387_ ? _0207_ : _1853_);
	assign _1883_ = _1881_ | _0127_;
	assign _1884_ = (_0146_ ? _1880_ : _1883_);
	assign _1885_ = (\mchip.pong.game.vga.pix_ind [0] ? _1884_ : _1876_);
	assign _1886_ = (_4387_ ? _0475_ : _0530_);
	assign _1887_ = (_0127_ ? _1878_ : _1886_);
	assign _1888_ = _0852_ | _4423_;
	assign _1889_ = (_4380_ ? _4408_ : _4427_);
	assign _1890_ = (_4387_ ? _0883_ : _1889_);
	assign _1891_ = (_0127_ ? _1888_ : _1890_);
	assign _1892_ = (_0146_ ? _1887_ : _1891_);
	assign _1894_ = (_0127_ ? _1829_ : _1886_);
	assign _1895_ = (_4423_ ? _0391_ : _0883_);
	assign _1896_ = (_0127_ ? _0550_ : _1895_);
	assign _1897_ = (_0146_ ? _1894_ : _1896_);
	assign _1898_ = (\mchip.pong.game.vga.pix_ind [0] ? _1897_ : _1892_);
	assign _1899_ = (_1103_ ? _1885_ : _1898_);
	assign _1900_ = (_4387_ ? _0054_ : _0530_);
	assign _1901_ = (_4387_ ? _0631_ : _0530_);
	assign _1902_ = (_0127_ ? _1900_ : _1901_);
	assign _1903_ = (_4389_ ? _4371_ : _4424_);
	assign _1905_ = ~(_1903_ & _4387_);
	assign _1906_ = (_0056_ ? _0834_ : _1905_);
	assign _1907_ = (_0146_ ? _1902_ : _1906_);
	assign _1908_ = ~_0608_;
	assign _1909_ = (_4423_ ? _0961_ : _1908_);
	assign _1910_ = (_4423_ ? _0117_ : _0639_);
	assign _1911_ = (_0127_ ? _1909_ : _1910_);
	assign _1912_ = (_4423_ ? _4409_ : _1853_);
	assign _1913_ = (_0127_ ? _0572_ : _1912_);
	assign _1914_ = (_0146_ ? _1911_ : _1913_);
	assign _1916_ = (\mchip.pong.game.vga.pix_ind [0] ? _1914_ : _1907_);
	assign _1917_ = (_4423_ ? _0530_ : _1908_);
	assign _1918_ = (_4423_ ? _0117_ : _0264_);
	assign _1919_ = (_0127_ ? _1917_ : _1918_);
	assign _1920_ = (_4423_ ? _4408_ : _0254_);
	assign _1921_ = (_0127_ ? _1888_ : _1920_);
	assign _1922_ = (_0146_ ? _1919_ : _1921_);
	assign _1923_ = (_4423_ ? _0852_ : _0472_);
	assign _1924_ = (_4387_ ? _4371_ : _0117_);
	assign _1925_ = (_0127_ ? _1923_ : _1924_);
	assign _1927_ = (_4380_ ? _4374_ : _0582_);
	assign _1928_ = (_4387_ ? _0070_ : _1927_);
	assign _1929_ = _1928_ | _0127_;
	assign _1930_ = (_0146_ ? _1925_ : _1929_);
	assign _1931_ = (\mchip.pong.game.vga.pix_ind [0] ? _1930_ : _1922_);
	assign _1932_ = (_1103_ ? _1916_ : _1931_);
	assign _1933_ = (_0044_ ? _1899_ : _1932_);
	assign _1934_ = (_4387_ ? _0495_ : _0792_);
	assign _1935_ = ~_1934_;
	assign _1936_ = (_4387_ ? _0451_ : _0852_);
	assign _1938_ = (_0127_ ? _1935_ : _1936_);
	assign _1939_ = (_0056_ ? _0098_ : _1649_);
	assign _1940_ = ~_1939_;
	assign _1941_ = (_0146_ ? _1938_ : _1940_);
	assign _1942_ = (_4423_ ? _0117_ : _4381_);
	assign _1943_ = (_4387_ ? _0451_ : _0101_);
	assign _1944_ = (_0127_ ? _1942_ : _1943_);
	assign _1945_ = (_4423_ ? _0792_ : _0207_);
	assign _1946_ = (_0056_ ? _0160_ : _1945_);
	assign _1947_ = (_0146_ ? _1944_ : _1946_);
	assign _1949_ = (\mchip.pong.game.vga.pix_ind [0] ? _1947_ : _1941_);
	assign _1950_ = (_4387_ ? _0451_ : _1853_);
	assign _1951_ = (_0127_ ? _1942_ : _1950_);
	assign _1952_ = (_4423_ ? _0119_ : _0426_);
	assign _1953_ = (_0056_ ? _0160_ : _1952_);
	assign _1954_ = (_0146_ ? _1951_ : _1953_);
	assign _1955_ = (_4387_ ? _4381_ : _0530_);
	assign _1956_ = _0631_ | _4423_;
	assign _1957_ = (_0127_ ? _1955_ : _1956_);
	assign _1959_ = ~_0872_;
	assign _1960_ = _0883_ | _4423_;
	assign _1961_ = (_0056_ ? _1959_ : _1960_);
	assign _1962_ = (_0146_ ? _1957_ : _1961_);
	assign _1963_ = (\mchip.pong.game.vga.pix_ind [0] ? _1962_ : _1954_);
	assign _1964_ = (_1103_ ? _1949_ : _1963_);
	assign _1965_ = (_4387_ ? _4443_ : _0117_);
	assign _1966_ = (_4387_ ? _4389_ : _0639_);
	assign _1967_ = (_0127_ ? _1965_ : _1966_);
	assign _1968_ = (_0146_ ? _1967_ : _1635_);
	assign _1970_ = (_4387_ ? _4389_ : _0117_);
	assign _1971_ = _4387_ & ~_0372_;
	assign _1972_ = ~_1971_;
	assign _1973_ = (_0127_ ? _1970_ : _1972_);
	assign _1974_ = (_0146_ ? _1973_ : _0135_);
	assign _1975_ = (\mchip.pong.game.vga.pix_ind [0] ? _1974_ : _1968_);
	assign _1976_ = (_4387_ ? _4409_ : _0114_);
	assign _1977_ = (_0127_ ? _1976_ : _0140_);
	assign _1978_ = (_0146_ ? _1977_ : _0135_);
	assign _1979_ = (_0056_ ? _1574_ : _1935_);
	assign _1981_ = _1846_ & ~_4423_;
	assign _1982_ = ~_1981_;
	assign _1983_ = (_0056_ ? _0098_ : _1982_);
	assign _1984_ = ~_1983_;
	assign _1985_ = (_0146_ ? _1979_ : _1984_);
	assign _1986_ = (\mchip.pong.game.vga.pix_ind [0] ? _1985_ : _1978_);
	assign _1987_ = (_1103_ ? _1975_ : _1986_);
	assign _1988_ = (_0044_ ? _1964_ : _1987_);
	assign _1989_ = (_0088_ ? _1933_ : _1988_);
	assign _1990_ = (_4387_ ? _0119_ : _0489_);
	assign _1992_ = _0127_ & ~_1990_;
	assign _1993_ = (_0146_ ? _1992_ : _1588_);
	assign _1994_ = (\mchip.pong.game.vga.pix_ind [0] ? _1993_ : _1698_);
	assign _1995_ = (_1103_ ? _1695_ : _1994_);
	assign _1996_ = (_0044_ ? _1995_ : _1691_);
	assign _1997_ = (_0088_ ? _1996_ : _1673_);
	assign _1998_ = (_4368_ ? _1989_ : _1997_);
	assign _1999_ = (_4367_ ? _1868_ : _1998_);
	assign _2000_ = _0127_ & ~_1965_;
	assign _2001_ = (_4387_ ? _4380_ : _0035_);
	assign _2003_ = _0056_ & ~_2001_;
	assign _2004_ = (_0146_ ? _2000_ : _2003_);
	assign _2005_ = \mchip.pong.game.vga.pix_ind [0] & ~_2004_;
	assign _2006_ = _0127_ & ~_1976_;
	assign _2007_ = (_4423_ ? _0054_ : _0280_);
	assign _2008_ = _0056_ & ~_2007_;
	assign _2009_ = (_0146_ ? _2006_ : _2008_);
	assign _2010_ = _4442_ & ~_2009_;
	assign _2011_ = _2010_ | _2005_;
	assign _2012_ = (_0056_ ? _0549_ : _0766_);
	assign _2014_ = _4387_ & ~_0035_;
	assign _2015_ = (_4407_ ? _4423_ : _4389_);
	assign _2016_ = (_0127_ ? _2014_ : _2015_);
	assign _2017_ = (_0146_ ? _2012_ : _2016_);
	assign _2018_ = _4442_ & ~_2017_;
	assign _2019_ = (_4423_ ? _0114_ : _4409_);
	assign _2020_ = _0056_ & ~_2019_;
	assign _2021_ = (_0146_ ? _0335_ : _2020_);
	assign _2022_ = _2021_ & ~_4442_;
	assign _2023_ = _2022_ | _2018_;
	assign _2025_ = (_1103_ ? _2011_ : _2023_);
	assign _2026_ = (_0044_ ? _1586_ : _2025_);
	assign _2027_ = (_0088_ ? _1568_ : _2026_);
	assign _2028_ = (_4380_ ? _4424_ : _0582_);
	assign _2029_ = (_4387_ ? _4381_ : _2028_);
	assign _2030_ = (_0056_ ? _0501_ : _2029_);
	assign _2031_ = ~_0367_;
	assign _2032_ = _2031_ | _4387_;
	assign _2033_ = (_0056_ ? _0770_ : _2032_);
	assign _2034_ = (_0146_ ? _2030_ : _2033_);
	assign _2036_ = (_4423_ ? _0292_ : _0089_);
	assign _2037_ = (_0127_ ? _1934_ : _2036_);
	assign _2038_ = ~_2037_;
	assign _2039_ = (_0127_ ? _0453_ : _0762_);
	assign _2040_ = (_0146_ ? _2038_ : _2039_);
	assign _2041_ = (\mchip.pong.game.vga.pix_ind [0] ? _2040_ : _2034_);
	assign _2042_ = _1934_ & ~_0056_;
	assign _2043_ = ~_2042_;
	assign _2044_ = _0784_ | _0127_;
	assign _2045_ = (_0146_ ? _2043_ : _2044_);
	assign _2047_ = ~_2006_;
	assign _2048_ = (_4423_ ? _0054_ : _0412_);
	assign _2049_ = _2048_ | _0127_;
	assign _2050_ = (_0146_ ? _2047_ : _2049_);
	assign _2051_ = (\mchip.pong.game.vga.pix_ind [0] ? _2050_ : _2045_);
	assign _2052_ = (_1103_ ? _2041_ : _2051_);
	assign _2053_ = ~_0054_;
	assign _2054_ = (_4387_ ? _2053_ : _0035_);
	assign _2055_ = ~(_2054_ & _0127_);
	assign _2056_ = (_4387_ ? _4428_ : _4409_);
	assign _2057_ = _2056_ | _0127_;
	assign _2058_ = (_0146_ ? _2055_ : _2057_);
	assign _2059_ = _0567_ | _0056_;
	assign _2060_ = _0834_ | _0127_;
	assign _2061_ = (_0146_ ? _2059_ : _2060_);
	assign _2062_ = (\mchip.pong.game.vga.pix_ind [0] ? _2061_ : _2058_);
	assign _2063_ = ~(_2062_ & _1103_);
	assign _2064_ = (_4423_ ? _4443_ : _4381_);
	assign _2065_ = _0127_ & ~_2064_;
	assign _2066_ = _0056_ & ~_0834_;
	assign _2068_ = (_0146_ ? _2065_ : _2066_);
	assign _2069_ = (_4423_ ? _0118_ : _4381_);
	assign _2070_ = _0127_ & ~_2069_;
	assign _2071_ = _0056_ & ~_0770_;
	assign _2072_ = (_0146_ ? _2070_ : _2071_);
	assign _2073_ = (\mchip.pong.game.vga.pix_ind [0] ? _2072_ : _2068_);
	assign _2074_ = ~(_2073_ | _1103_);
	assign _2075_ = _2074_ | ~_2063_;
	assign _2076_ = (_0044_ ? _2052_ : _2075_);
	assign _2077_ = (_4387_ ? _0421_ : _0107_);
	assign _2079_ = (_0127_ ? _1555_ : _2077_);
	assign _2080_ = (_4423_ ? _0113_ : _0114_);
	assign _2081_ = (_0127_ ? _0500_ : _2080_);
	assign _2082_ = ~_2081_;
	assign _2083_ = (_0146_ ? _2079_ : _2082_);
	assign _2084_ = (_4423_ ? _0454_ : _0361_);
	assign _2085_ = _0421_ | _4423_;
	assign _2086_ = (_0127_ ? _2084_ : _2085_);
	assign _2087_ = _0820_ | _4423_;
	assign _2088_ = (_0056_ ? _0793_ : _2087_);
	assign _2090_ = (_0146_ ? _2086_ : _2088_);
	assign _2091_ = (\mchip.pong.game.vga.pix_ind [0] ? _2090_ : _2083_);
	assign _2092_ = (_4387_ ? _0054_ : _1024_);
	assign _2093_ = (_0056_ ? _0501_ : _2092_);
	assign _2094_ = (_4387_ ? _4428_ : _4434_);
	assign _2095_ = (_0127_ ? _0448_ : _2094_);
	assign _2096_ = (_0146_ ? _2093_ : _2095_);
	assign _2097_ = ~_2036_;
	assign _2098_ = (_4387_ ? _0054_ : _0114_);
	assign _2099_ = (_0056_ ? _2097_ : _2098_);
	assign _2101_ = (_0127_ ? _2085_ : _2094_);
	assign _2102_ = (_0146_ ? _2099_ : _2101_);
	assign _2103_ = (\mchip.pong.game.vga.pix_ind [0] ? _2102_ : _2096_);
	assign _2104_ = (_1103_ ? _2091_ : _2103_);
	assign _2105_ = (_4423_ ? _4443_ : _0035_);
	assign _2106_ = (_0056_ ? _0453_ : _2105_);
	assign _2107_ = (_0146_ ? _2106_ : _2082_);
	assign _2108_ = (_4423_ ? _0206_ : _0035_);
	assign _2109_ = (_4387_ ? _0421_ : _0451_);
	assign _2110_ = (_0127_ ? _2108_ : _2109_);
	assign _2112_ = (_0127_ ? _0875_ : _2080_);
	assign _2113_ = ~_2112_;
	assign _2114_ = (_0146_ ? _2110_ : _2113_);
	assign _2115_ = (\mchip.pong.game.vga.pix_ind [0] ? _2114_ : _2107_);
	assign _2116_ = (_0127_ ? _1555_ : _2109_);
	assign _2117_ = (_0146_ ? _2116_ : _2113_);
	assign _2118_ = (_1103_ ? _2115_ : _2117_);
	assign _2119_ = (_0044_ ? _2104_ : _2118_);
	assign _2120_ = (_0088_ ? _2076_ : _2119_);
	assign _2121_ = (_4368_ ? _2027_ : _2120_);
	assign _2123_ = (_4423_ ? _0117_ : _0361_);
	assign _2124_ = (_0056_ ? _0140_ : _2123_);
	assign _2125_ = _0056_ & ~_0793_;
	assign _2126_ = ~_2125_;
	assign _2127_ = (_0146_ ? _2124_ : _2126_);
	assign _2128_ = (_4423_ ? _4389_ : _0035_);
	assign _2129_ = (_0056_ ? _1818_ : _2128_);
	assign _2130_ = (_0146_ ? _2129_ : _2113_);
	assign _2131_ = (\mchip.pong.game.vga.pix_ind [0] ? _2130_ : _2127_);
	assign _2132_ = _0127_ & ~_2128_;
	assign _2134_ = ~_2132_;
	assign _2135_ = (_0127_ ? _1737_ : _0793_);
	assign _2136_ = (_0146_ ? _2134_ : _2135_);
	assign _2137_ = _4387_ & ~_0871_;
	assign _2138_ = (_0056_ ? _2080_ : _2137_);
	assign _2139_ = ~_2138_;
	assign _2140_ = (_0146_ ? _2134_ : _2139_);
	assign _2141_ = (\mchip.pong.game.vga.pix_ind [0] ? _2140_ : _2136_);
	assign _2142_ = (_1103_ ? _2131_ : _2141_);
	assign _2143_ = (_4387_ ? _0054_ : _0903_);
	assign _2145_ = (_4387_ ? _0421_ : _0372_);
	assign _2146_ = (_0127_ ? _2143_ : _2145_);
	assign _2147_ = (_0056_ ? _0834_ : _1972_);
	assign _2148_ = (_0146_ ? _2146_ : _2147_);
	assign _2149_ = (_4387_ ? _0054_ : _0100_);
	assign _2150_ = (_0056_ ? _2145_ : _2149_);
	assign _2151_ = (_0146_ ? _2150_ : _2057_);
	assign _2152_ = (\mchip.pong.game.vga.pix_ind [0] ? _2151_ : _2148_);
	assign _2153_ = (_4387_ ? _0054_ : _0153_);
	assign _2154_ = (_0056_ ? _2145_ : _2153_);
	assign _2156_ = (_0146_ ? _2154_ : _2060_);
	assign _2157_ = (_4387_ ? _0054_ : _0989_);
	assign _2158_ = (_0056_ ? _2145_ : _2157_);
	assign _2159_ = _0056_ & ~_0823_;
	assign _2160_ = ~_2159_;
	assign _2161_ = (_0146_ ? _2158_ : _2160_);
	assign _2162_ = (\mchip.pong.game.vga.pix_ind [0] ? _2161_ : _2156_);
	assign _2163_ = (_1103_ ? _2152_ : _2162_);
	assign _2164_ = (_0044_ ? _2142_ : _2163_);
	assign _2165_ = (_4423_ ? _0421_ : _0451_);
	assign _2167_ = (_0127_ ? _0154_ : _2165_);
	assign _2168_ = ~(_0094_ & _4387_);
	assign _2169_ = (_0056_ ? _0972_ : _2168_);
	assign _2170_ = (_0146_ ? _2167_ : _2169_);
	assign _2171_ = (_0056_ ? _0140_ : _2069_);
	assign _2172_ = (_4423_ ? _0421_ : _0372_);
	assign _2173_ = (_4387_ ? _4380_ : _0153_);
	assign _2174_ = (_0127_ ? _2172_ : _2173_);
	assign _2175_ = (_0146_ ? _2171_ : _2174_);
	assign _2176_ = (\mchip.pong.game.vga.pix_ind [0] ? _2175_ : _2170_);
	assign _2178_ = (_4387_ ? _0114_ : _0372_);
	assign _2179_ = (_0127_ ? _0048_ : _2178_);
	assign _2180_ = (_0127_ ? _1924_ : _2153_);
	assign _2181_ = (_0146_ ? _2179_ : _2180_);
	assign _2182_ = (_0127_ ? _0048_ : _2145_);
	assign _2183_ = (_4423_ ? _0100_ : _0035_);
	assign _2184_ = (_0127_ ? _0572_ : _2183_);
	assign _2185_ = (_0146_ ? _2182_ : _2184_);
	assign _2186_ = (\mchip.pong.game.vga.pix_ind [0] ? _2185_ : _2181_);
	assign _2187_ = (_1103_ ? _2176_ : _2186_);
	assign _2189_ = _4387_ & ~_0254_;
	assign _2190_ = ~_2189_;
	assign _2191_ = (_4387_ ? _4443_ : _0114_);
	assign _2192_ = (_0056_ ? _2190_ : _2191_);
	assign _2193_ = (_4380_ ? _4408_ : _0065_);
	assign _2194_ = (_4423_ ? _0961_ : _2193_);
	assign _2195_ = (_0056_ ? _2001_ : _2194_);
	assign _2196_ = (_0146_ ? _2192_ : _2195_);
	assign _2197_ = (_4387_ ? _0845_ : _4437_);
	assign _2198_ = (_0056_ ? _2085_ : _2197_);
	assign _2200_ = (_4374_ ? _4372_ : _4380_);
	assign _2201_ = ~_2200_;
	assign _2202_ = (_4389_ ? _4375_ : _4419_);
	assign _2203_ = ~_2202_;
	assign _2204_ = (_4412_ ? _2201_ : _2203_);
	assign _2205_ = (_0056_ ? _1764_ : _2204_);
	assign _2206_ = (_0146_ ? _2198_ : _2205_);
	assign _2207_ = (\mchip.pong.game.vga.pix_ind [0] ? _2206_ : _2196_);
	assign _2208_ = (_4423_ ? _0444_ : _0490_);
	assign _2209_ = (_4423_ ? _0054_ : _1010_);
	assign _2211_ = (_0127_ ? _2208_ : _2209_);
	assign _2212_ = (_0146_ ? _2047_ : _2211_);
	assign _2213_ = (_4423_ ? _0118_ : _0153_);
	assign _2214_ = (_0056_ ? _0755_ : _2213_);
	assign _2215_ = (_4423_ ? _0119_ : _0530_);
	assign _2216_ = (_4423_ ? _4381_ : _0957_);
	assign _2217_ = (_0127_ ? _2215_ : _2216_);
	assign _2218_ = (_0146_ ? _2214_ : _2217_);
	assign _2219_ = (\mchip.pong.game.vga.pix_ind [0] ? _2218_ : _2212_);
	assign _2220_ = (_1103_ ? _2207_ : _2219_);
	assign _2222_ = (_0044_ ? _2187_ : _2220_);
	assign _2223_ = (_0088_ ? _2164_ : _2222_);
	assign _2224_ = _0254_ | _4387_;
	assign _2225_ = (_4371_ ? _4423_ : _4389_);
	assign _2226_ = (_0056_ ? _2224_ : _2225_);
	assign _2227_ = _4423_ | _4409_;
	assign _2228_ = (_0127_ ? _2227_ : _0334_);
	assign _2229_ = ~_2228_;
	assign _2230_ = (_0146_ ? _2226_ : _2229_);
	assign _2231_ = (_4387_ ? _0118_ : _0372_);
	assign _2233_ = _0127_ & ~_2231_;
	assign _2234_ = ~_2233_;
	assign _2235_ = ~_0330_;
	assign _2236_ = (_4423_ ? _4428_ : _0403_);
	assign _2237_ = (_0056_ ? _2235_ : _2236_);
	assign _2238_ = (_0146_ ? _2234_ : _2237_);
	assign _2239_ = (\mchip.pong.game.vga.pix_ind [0] ? _2238_ : _2230_);
	assign _2240_ = (_1103_ ? _1695_ : _2239_);
	assign _2241_ = (_0044_ ? _2240_ : _1691_);
	assign _2242_ = (_0088_ ? _2241_ : _1673_);
	assign _2244_ = (_4368_ ? _2223_ : _2242_);
	assign _2245_ = (_4367_ ? _2121_ : _2244_);
	assign _2246_ = (_1058_ ? _2245_ : _1706_);
	assign _2247_ = (_0723_ ? _1999_ : _2246_);
	assign _2248_ = (_1061_ ? _1706_ : _2247_);
	assign \mchip.pong.VGA_G3  = (_1264_ ? _2248_ : _1519_);
	assign _2249_ = ~_0115_;
	assign _2250_ = _0660_ & ~_4387_;
	assign _2251_ = (_0056_ ? _2249_ : _2250_);
	assign _2252_ = (_0146_ ? _0349_ : _2251_);
	assign _2254_ = (\mchip.pong.game.vga.pix_ind [0] ? _0112_ : _2252_);
	assign _2255_ = (_1103_ ? _2254_ : _0106_);
	assign _2256_ = ~(_0035_ | _4417_);
	assign _2257_ = ~_2256_;
	assign _2258_ = (_4387_ ? _0206_ : _2257_);
	assign _2259_ = (_0127_ ? _0356_ : _2258_);
	assign _2260_ = (_4423_ ? _0118_ : _0361_);
	assign _2261_ = (_0056_ ? _0035_ : _2260_);
	assign _2262_ = (_0146_ ? _2259_ : _2261_);
	assign _2263_ = (_4380_ ? _4427_ : _4408_);
	assign _2265_ = (_4387_ ? _4417_ : _2263_);
	assign _2266_ = (_0127_ ? _0365_ : _2265_);
	assign _2267_ = (_4423_ ? _4443_ : _0366_);
	assign _2268_ = (_4423_ ? _0054_ : _4390_);
	assign _2269_ = (_0127_ ? _2267_ : _2268_);
	assign _2270_ = (_0146_ ? _2266_ : _2269_);
	assign _2271_ = (\mchip.pong.game.vga.pix_ind [0] ? _2270_ : _2262_);
	assign _2272_ = ~(_4387_ | _4427_);
	assign _2273_ = (_0127_ ? _0378_ : _2272_);
	assign _2274_ = (_4423_ ? _0421_ : _0101_);
	assign _2276_ = (_0056_ ? _0792_ : _2274_);
	assign _2277_ = (_0146_ ? _2273_ : _2276_);
	assign _2278_ = (_4380_ ? _4424_ : _4375_);
	assign _2279_ = _2278_ & ~_4387_;
	assign _2280_ = (_0127_ ? _0386_ : _2279_);
	assign _2281_ = (_0056_ ? _0390_ : _0402_);
	assign _2282_ = (_0146_ ? _2280_ : _2281_);
	assign _2283_ = (\mchip.pong.game.vga.pix_ind [0] ? _2282_ : _2277_);
	assign _2284_ = (_1103_ ? _2271_ : _2283_);
	assign _2285_ = (_0044_ ? _2255_ : _2284_);
	assign _2287_ = (_0088_ ? _0084_ : _2285_);
	assign _2288_ = (_4387_ ? _0671_ : _0792_);
	assign _2289_ = (_0127_ ? _0154_ : _2288_);
	assign _2290_ = (_4380_ ? _0577_ : _0582_);
	assign _2291_ = (_4423_ ? _4381_ : _2290_);
	assign _2292_ = _2291_ & ~_0127_;
	assign _2293_ = (_0146_ ? _2289_ : _2292_);
	assign _2294_ = (_4423_ ? _4380_ : _4443_);
	assign _2295_ = (_0127_ ? _0048_ : _2294_);
	assign _2296_ = _4387_ & ~_0426_;
	assign _2298_ = (_4387_ ? _0100_ : _0153_);
	assign _2299_ = (_0127_ ? _2296_ : _2298_);
	assign _2300_ = (_0146_ ? _2295_ : _2299_);
	assign _2301_ = (\mchip.pong.game.vga.pix_ind [0] ? _2300_ : _2293_);
	assign _2302_ = (_4387_ ? _4413_ : _0961_);
	assign _2303_ = (_0127_ ? _0399_ : _2302_);
	assign _2304_ = (_4423_ ? _0054_ : _0542_);
	assign _2305_ = (_0127_ ? _0386_ : _2304_);
	assign _2306_ = (_0146_ ? _2303_ : _2305_);
	assign _2307_ = _0118_ | ~_0114_;
	assign _2309_ = (_4387_ ? _4417_ : _2307_);
	assign _2310_ = (_0127_ ? _0154_ : _2309_);
	assign _2311_ = (_4423_ ? _4381_ : _0035_);
	assign _2312_ = (_4387_ ? _0280_ : _4381_);
	assign _2313_ = (_0127_ ? _2311_ : _2312_);
	assign _2314_ = (_0146_ ? _2310_ : _2313_);
	assign _2315_ = (\mchip.pong.game.vga.pix_ind [0] ? _2314_ : _2306_);
	assign _2316_ = (_1103_ ? _2301_ : _2315_);
	assign _2317_ = (_4387_ ? _0425_ : _4391_);
	assign _2318_ = _0127_ & ~_2317_;
	assign _2320_ = (_4423_ ? _0113_ : _0478_);
	assign _2321_ = _0056_ & ~_2320_;
	assign _2322_ = (_0146_ ? _2318_ : _2321_);
	assign _2323_ = (_4387_ ? _0599_ : _0442_);
	assign _2324_ = _2323_ & ~_0056_;
	assign _2325_ = (_4423_ ? _0153_ : _0613_);
	assign _2326_ = (_0127_ ? _0208_ : _2325_);
	assign _2327_ = (_0146_ ? _2324_ : _2326_);
	assign _2328_ = (\mchip.pong.game.vga.pix_ind [0] ? _2327_ : _2322_);
	assign _2329_ = _1908_ & ~_4423_;
	assign _2331_ = ~_1679_;
	assign _2332_ = (_0127_ ? _2329_ : _2331_);
	assign _2333_ = (_4423_ ? _0153_ : _0568_);
	assign _2334_ = (_0127_ ? _0208_ : _2333_);
	assign _2335_ = (_0146_ ? _2332_ : _2334_);
	assign _2336_ = ~(_0207_ | _4423_);
	assign _2337_ = (_0127_ ? _0179_ : _2336_);
	assign _2338_ = (_4389_ ? _4408_ : _4433_);
	assign _2339_ = _4423_ & ~_2338_;
	assign _2340_ = (_4387_ ? _4408_ : _4409_);
	assign _2342_ = (_0127_ ? _2339_ : _2340_);
	assign _2343_ = (_0146_ ? _2337_ : _2342_);
	assign _2344_ = (\mchip.pong.game.vga.pix_ind [0] ? _2343_ : _2335_);
	assign _2345_ = (_1103_ ? _2328_ : _2344_);
	assign _2346_ = (_0044_ ? _2316_ : _2345_);
	assign _2347_ = _2263_ & ~_4387_;
	assign _2348_ = (_0127_ ? _2092_ : _2347_);
	assign _2349_ = _4408_ & ~_4423_;
	assign _2350_ = (_4387_ ? _0852_ : _0687_);
	assign _2351_ = (_0127_ ? _2349_ : _2350_);
	assign _2353_ = (_0146_ ? _2348_ : _2351_);
	assign _2354_ = (_4387_ ? _4417_ : _4427_);
	assign _2355_ = (_0127_ ? _0484_ : _2354_);
	assign _2356_ = _1870_ & ~_4423_;
	assign _2357_ = (_4387_ ? _0852_ : _0490_);
	assign _2358_ = (_0127_ ? _2356_ : _2357_);
	assign _2359_ = (_0146_ ? _2355_ : _2358_);
	assign _2360_ = (\mchip.pong.game.vga.pix_ind [0] ? _2359_ : _2353_);
	assign _2361_ = (_4380_ ? _4371_ : _4408_);
	assign _2362_ = _2361_ & ~_4387_;
	assign _2364_ = (_0127_ ? _1555_ : _2362_);
	assign _2365_ = _1020_ & ~_4423_;
	assign _2366_ = (_0056_ ? _4389_ : _2365_);
	assign _2367_ = (_0146_ ? _2364_ : _2366_);
	assign _2368_ = _1630_ | _0226_;
	assign _2369_ = (_4423_ ? _4380_ : _0478_);
	assign _2370_ = _0056_ & ~_2369_;
	assign _2371_ = (_0146_ ? _2368_ : _2370_);
	assign _2372_ = (\mchip.pong.game.vga.pix_ind [0] ? _2371_ : _2367_);
	assign _2373_ = (_1103_ ? _2360_ : _2372_);
	assign _2375_ = (_4387_ ? _0203_ : _0067_);
	assign _2376_ = (_4380_ ? _4372_ : _4424_);
	assign _2377_ = (_4387_ ? _4413_ : _2376_);
	assign _2378_ = (_0127_ ? _2375_ : _2377_);
	assign _2379_ = (_4412_ ? _4437_ : _0100_);
	assign _2380_ = (_4387_ ? _4389_ : _0045_);
	assign _2381_ = (_0127_ ? _2379_ : _2380_);
	assign _2382_ = (_0146_ ? _2378_ : _2381_);
	assign _2383_ = (_4387_ ? _0203_ : _0119_);
	assign _2385_ = (_4423_ ? _4372_ : _0206_);
	assign _2386_ = (_0127_ ? _2383_ : _2385_);
	assign _2387_ = _4387_ & ~_0100_;
	assign _2388_ = (_4387_ ? _0568_ : _0045_);
	assign _2389_ = (_0127_ ? _2387_ : _2388_);
	assign _2390_ = (_0146_ ? _2386_ : _2389_);
	assign _2391_ = (\mchip.pong.game.vga.pix_ind [0] ? _2390_ : _2382_);
	assign _2392_ = (_4423_ ? _0119_ : _0472_);
	assign _2393_ = (_4380_ ? _4424_ : _0756_);
	assign _2394_ = (_4387_ ? _0118_ : _2393_);
	assign _2396_ = (_0127_ ? _2392_ : _2394_);
	assign _2397_ = (_0127_ ? _4387_ : _2388_);
	assign _2398_ = (_0146_ ? _2396_ : _2397_);
	assign _2399_ = (_4387_ ? _0054_ : _0451_);
	assign _2400_ = _0366_ | _0066_;
	assign _2401_ = (_4387_ ? _4417_ : _2400_);
	assign _2402_ = (_0127_ ? _2399_ : _2401_);
	assign _2403_ = (_4389_ ? _4433_ : _4407_);
	assign _2404_ = _4387_ & ~_2403_;
	assign _2406_ = (_4387_ ? _0568_ : _1808_);
	assign _2407_ = (_0127_ ? _2404_ : _2406_);
	assign _2408_ = (_0146_ ? _2402_ : _2407_);
	assign _2409_ = (\mchip.pong.game.vga.pix_ind [0] ? _2408_ : _2398_);
	assign _2410_ = (_1103_ ? _2391_ : _2409_);
	assign _2411_ = (_0044_ ? _2373_ : _2410_);
	assign _2412_ = (_0088_ ? _2346_ : _2411_);
	assign _2413_ = (_4368_ ? _2287_ : _2412_);
	assign _2414_ = (_4423_ ? _4380_ : _0871_);
	assign _2415_ = (_4423_ ? _0066_ : _0314_);
	assign _2417_ = (_0127_ ? _2414_ : _2415_);
	assign _2418_ = (_4387_ ? _4428_ : _0114_);
	assign _2419_ = (_4423_ ? _4408_ : _1889_);
	assign _2420_ = (_0127_ ? _2418_ : _2419_);
	assign _2421_ = (_0146_ ? _2417_ : _2420_);
	assign _2422_ = (_4423_ ? _1010_ : _0472_);
	assign _2423_ = (_4389_ ? _4374_ : _4419_);
	assign _2424_ = (_4423_ ? _4425_ : _2423_);
	assign _2425_ = (_0127_ ? _2422_ : _2424_);
	assign _2426_ = (_4387_ ? _4428_ : _1809_);
	assign _2428_ = (_4387_ ? _0568_ : _1790_);
	assign _2429_ = (_0127_ ? _2426_ : _2428_);
	assign _2430_ = (_0146_ ? _2425_ : _2429_);
	assign _2431_ = (\mchip.pong.game.vga.pix_ind [0] ? _2430_ : _2421_);
	assign _2432_ = (_4389_ ? _4374_ : _4408_);
	assign _2433_ = (_4387_ ? _0472_ : _2432_);
	assign _2434_ = (_4389_ ? _0577_ : _4419_);
	assign _2435_ = (_4423_ ? _4390_ : _2434_);
	assign _2436_ = (_0127_ ? _2433_ : _2435_);
	assign _2437_ = (_4387_ ? _4380_ : _0454_);
	assign _2439_ = (_4387_ ? _0961_ : _0506_);
	assign _2440_ = (_0127_ ? _2437_ : _2439_);
	assign _2441_ = (_0146_ ? _2436_ : _2440_);
	assign _2442_ = (_4423_ ? _4380_ : _1908_);
	assign _2443_ = (_4387_ ? _4417_ : _0054_);
	assign _2444_ = (_0127_ ? _2442_ : _2443_);
	assign _2445_ = (_4387_ ? _4375_ : _1020_);
	assign _2446_ = (_4387_ ? _4391_ : _0506_);
	assign _2447_ = (_0127_ ? _2445_ : _2446_);
	assign _2448_ = (_0146_ ? _2444_ : _2447_);
	assign _2450_ = (\mchip.pong.game.vga.pix_ind [0] ? _2448_ : _2441_);
	assign _2451_ = (_1103_ ? _2431_ : _2450_);
	assign _2452_ = (_4423_ ? _0417_ : _0599_);
	assign _2453_ = (_4423_ ? _0280_ : _0101_);
	assign _2454_ = (_0127_ ? _2452_ : _2453_);
	assign _2455_ = (_4423_ ? _0852_ : _0599_);
	assign _2456_ = (_4389_ ? _4374_ : _4375_);
	assign _2457_ = (_4423_ ? _0153_ : _2456_);
	assign _2458_ = (_0127_ ? _2455_ : _2457_);
	assign _2459_ = (_0146_ ? _2454_ : _2458_);
	assign _2461_ = (_0276_ ? _0067_ : _4437_);
	assign _2462_ = (_4389_ ? _4371_ : _4387_);
	assign _2463_ = (_0127_ ? _2461_ : _2462_);
	assign _2464_ = (_4387_ ? _0678_ : _0444_);
	assign _2465_ = (_4380_ ? _4371_ : _0756_);
	assign _2466_ = (_4423_ ? _0623_ : _2465_);
	assign _2467_ = (_0127_ ? _2464_ : _2466_);
	assign _2468_ = (_0146_ ? _2463_ : _2467_);
	assign _2469_ = (\mchip.pong.game.vga.pix_ind [0] ? _2468_ : _2459_);
	assign _2470_ = (_4423_ ? _4380_ : _0506_);
	assign _2472_ = (_4371_ ? _4389_ : _4374_);
	assign _2473_ = (_4387_ ? _1870_ : _2472_);
	assign _2474_ = (_0127_ ? _2470_ : _2473_);
	assign _2475_ = (_4389_ ? _4408_ : _0577_);
	assign _2476_ = (_4423_ ? _2475_ : _2456_);
	assign _2477_ = _0359_ | _4387_;
	assign _2478_ = (_0127_ ? _2476_ : _2477_);
	assign _2479_ = (_0146_ ? _2474_ : _2478_);
	assign _2480_ = (_4423_ ? _0404_ : _2257_);
	assign _2481_ = (_4387_ ? _0989_ : _0479_);
	assign _2483_ = (_0127_ ? _2480_ : _2481_);
	assign _2484_ = (_4374_ ? _4372_ : _0970_);
	assign _2485_ = _2484_ | _4423_;
	assign _2486_ = (_4380_ ? _4427_ : _0582_);
	assign _2487_ = (_4423_ ? _0093_ : _2486_);
	assign _2488_ = (_0127_ ? _2485_ : _2487_);
	assign _2489_ = (_0146_ ? _2483_ : _2488_);
	assign _2490_ = (\mchip.pong.game.vga.pix_ind [0] ? _2489_ : _2479_);
	assign _2491_ = (_1103_ ? _2469_ : _2490_);
	assign _2492_ = (_0044_ ? _2451_ : _2491_);
	assign _2494_ = (_4387_ ? _4381_ : _0560_);
	assign _2495_ = (_4380_ ? _0577_ : _4427_);
	assign _2496_ = (_4387_ ? _0820_ : _2495_);
	assign _2497_ = (_0127_ ? _2494_ : _2496_);
	assign _2498_ = _0235_ | _0161_;
	assign _2499_ = (_0146_ ? _2497_ : _2498_);
	assign _2500_ = (_4423_ ? _0421_ : _0153_);
	assign _2501_ = (_4389_ ? _4374_ : _4424_);
	assign _2502_ = (_4387_ ? _2031_ : _2501_);
	assign _2503_ = (_0127_ ? _2500_ : _2502_);
	assign _2505_ = (_0056_ ? _0429_ : _0861_);
	assign _2506_ = (_0146_ ? _2503_ : _2505_);
	assign _2507_ = (\mchip.pong.game.vga.pix_ind [0] ? _2506_ : _2499_);
	assign _2508_ = (_4387_ ? _0665_ : _2475_);
	assign _2509_ = (_4423_ ? _0660_ : _1853_);
	assign _2510_ = (_0127_ ? _2508_ : _2509_);
	assign _2511_ = (_4387_ ? _4419_ : _1781_);
	assign _2512_ = (_0056_ ? _0670_ : _2511_);
	assign _2513_ = (_0146_ ? _2510_ : _2512_);
	assign _2514_ = (_4387_ ? _0054_ : _2290_);
	assign _2516_ = (_4387_ ? _0101_ : _2376_);
	assign _2517_ = (_0127_ ? _2514_ : _2516_);
	assign _2518_ = ~_0237_;
	assign _2519_ = (_4423_ ? _0372_ : _0613_);
	assign _2520_ = (_0056_ ? _2518_ : _2519_);
	assign _2521_ = (_0146_ ? _2517_ : _2520_);
	assign _2522_ = (\mchip.pong.game.vga.pix_ind [0] ? _2521_ : _2513_);
	assign _2523_ = (_1103_ ? _2507_ : _2522_);
	assign _2524_ = (_4387_ ? _4389_ : _0442_);
	assign _2525_ = (_4389_ ? _4419_ : _0582_);
	assign _2527_ = (_4387_ ? _0687_ : _2525_);
	assign _2528_ = (_0127_ ? _2524_ : _2527_);
	assign _2529_ = (_0146_ ? _2528_ : _0242_);
	assign _2530_ = (_4423_ ? _0454_ : _4434_);
	assign _2531_ = (_4423_ ? _4389_ : _0117_);
	assign _2532_ = (_0127_ ? _2530_ : _2531_);
	assign _2533_ = (_0146_ ? _2532_ : _0126_);
	assign _2534_ = (\mchip.pong.game.vga.pix_ind [0] ? _2533_ : _2529_);
	assign _2535_ = (_4380_ ? _4372_ : _0582_);
	assign _2536_ = (_4387_ ? _0153_ : _2535_);
	assign _2538_ = (_4387_ ? _0206_ : _0093_);
	assign _2539_ = (_0127_ ? _2536_ : _2538_);
	assign _2540_ = (_0146_ ? _2539_ : _0156_);
	assign _2541_ = (_4387_ ? _4409_ : _2535_);
	assign _2542_ = (_4387_ ? _0206_ : _0372_);
	assign _2543_ = (_0127_ ? _2541_ : _2542_);
	assign _2544_ = (_0146_ ? _2543_ : _0706_);
	assign _2545_ = (\mchip.pong.game.vga.pix_ind [0] ? _2544_ : _2540_);
	assign _2546_ = (_1103_ ? _2534_ : _2545_);
	assign _2547_ = (_0044_ ? _2523_ : _2546_);
	assign _2549_ = (_0088_ ? _2492_ : _2547_);
	assign _2550_ = (_4423_ ? _0107_ : _0113_);
	assign _2551_ = _0127_ & ~_2550_;
	assign _2552_ = (_0146_ ? _2551_ : _0340_);
	assign _2553_ = (\mchip.pong.game.vga.pix_ind [0] ? _2552_ : _0339_);
	assign _2554_ = (_1103_ ? _0337_ : _2553_);
	assign _2555_ = (_0044_ ? _2554_ : _0329_);
	assign _2556_ = (_0088_ ? _2555_ : _0307_);
	assign _2557_ = (_4368_ ? _2549_ : _2556_);
	assign _2558_ = (_4367_ ? _2413_ : _2557_);
	assign _2560_ = (_4423_ ? _4417_ : _0153_);
	assign _2561_ = (_0056_ ? _0755_ : _2560_);
	assign _2562_ = (_0146_ ? _2561_ : _0763_);
	assign _2563_ = (\mchip.pong.game.vga.pix_ind [0] ? _0772_ : _2562_);
	assign _2564_ = (_1103_ ? _2563_ : _0788_);
	assign _2565_ = (_4380_ ? _4424_ : _0065_);
	assign _2566_ = (_4387_ ? _4381_ : _2565_);
	assign _2567_ = _2566_ | _0056_;
	assign _2568_ = (_0146_ ? _2567_ : _0799_);
	assign _2569_ = (\mchip.pong.game.vga.pix_ind [0] ? _2568_ : _0795_);
	assign _2571_ = (_4387_ ? _0054_ : _0454_);
	assign _2572_ = (_0056_ ? _0193_ : _2571_);
	assign _2573_ = (_0146_ ? _2572_ : _0799_);
	assign _2574_ = (\mchip.pong.game.vga.pix_ind [0] ? _0812_ : _2573_);
	assign _2575_ = (_1103_ ? _2569_ : _2574_);
	assign _2576_ = (_0044_ ? _2564_ : _2575_);
	assign _2577_ = (_4423_ ? _4437_ : _0957_);
	assign _2578_ = (_0127_ ? _0816_ : _2577_);
	assign _2579_ = (_0146_ ? _2578_ : _0824_);
	assign _2580_ = (_4387_ ? _4380_ : _0579_);
	assign _2582_ = (_4423_ ? _0114_ : _0957_);
	assign _2583_ = (_0127_ ? _2580_ : _2582_);
	assign _2584_ = (_0146_ ? _2583_ : _0835_);
	assign _2585_ = (\mchip.pong.game.vga.pix_ind [0] ? _2584_ : _2579_);
	assign _2586_ = (_4423_ ? _0114_ : _0542_);
	assign _2587_ = (_0127_ ? _0838_ : _2586_);
	assign _2588_ = (_0146_ ? _2587_ : _0847_);
	assign _2589_ = (\mchip.pong.game.vga.pix_ind [0] ? _0858_ : _2588_);
	assign _2590_ = (_1103_ ? _2585_ : _2589_);
	assign _2591_ = (_4423_ ? _0890_ : _0603_);
	assign _2593_ = (_0127_ ? _0861_ : _2591_);
	assign _2594_ = (_0146_ ? _2593_ : _0868_);
	assign _2595_ = (_4387_ ? _0203_ : _0757_);
	assign _2596_ = (_0056_ ? _0872_ : _2595_);
	assign _2597_ = (_0146_ ? _2596_ : _0877_);
	assign _2598_ = (\mchip.pong.game.vga.pix_ind [0] ? _2597_ : _2594_);
	assign _2599_ = (_4387_ ? _0119_ : _0883_);
	assign _2600_ = (_0127_ ? _0881_ : _2599_);
	assign _2601_ = (_0146_ ? _2600_ : _0887_);
	assign _2602_ = (_4387_ ? _0054_ : _0403_);
	assign _2604_ = (_4387_ ? _0090_ : _0672_);
	assign _2605_ = (_0127_ ? _2602_ : _2604_);
	assign _2606_ = (_0146_ ? _2605_ : _0894_);
	assign _2607_ = (\mchip.pong.game.vga.pix_ind [0] ? _2606_ : _2601_);
	assign _2608_ = (_1103_ ? _2598_ : _2607_);
	assign _2609_ = (_0044_ ? _2590_ : _2608_);
	assign _2610_ = (_0088_ ? _2576_ : _2609_);
	assign _2611_ = (_4368_ ? _0752_ : _2610_);
	assign _2612_ = (_0127_ ? _0484_ : _0902_);
	assign _2613_ = (_0127_ ? _0550_ : _0834_);
	assign _2615_ = (_0146_ ? _2612_ : _2613_);
	assign _2616_ = (\mchip.pong.game.vga.pix_ind [0] ? _0911_ : _2615_);
	assign _2617_ = (_0056_ ? _0902_ : _0913_);
	assign _2618_ = (_0146_ ? _2617_ : _0917_);
	assign _2619_ = (_0056_ ? _0914_ : _2143_);
	assign _2620_ = (_4387_ ? _4371_ : _0421_);
	assign _2621_ = (_0056_ ? _0867_ : _2620_);
	assign _2622_ = (_0146_ ? _2619_ : _2621_);
	assign _2623_ = (\mchip.pong.game.vga.pix_ind [0] ? _2622_ : _2618_);
	assign _2624_ = (_1103_ ? _2616_ : _2623_);
	assign _2626_ = (_4423_ ? _4389_ : _4381_);
	assign _2627_ = (_0056_ ? _0933_ : _2626_);
	assign _2628_ = (_0146_ ? _2627_ : _0930_);
	assign _2629_ = (_4387_ ? _4437_ : _0880_);
	assign _2630_ = (_0056_ ? _0933_ : _2629_);
	assign _2631_ = (_0146_ ? _2630_ : _0935_);
	assign _2632_ = (\mchip.pong.game.vga.pix_ind [0] ? _2631_ : _2628_);
	assign _2633_ = (_4387_ ? _0035_ : _2565_);
	assign _2634_ = (_0056_ ? _0940_ : _2633_);
	assign _2635_ = (_0146_ ? _2634_ : _0944_);
	assign _2637_ = (\mchip.pong.game.vga.pix_ind [0] ? _0952_ : _2635_);
	assign _2638_ = (_1103_ ? _2632_ : _2637_);
	assign _2639_ = (_0044_ ? _2624_ : _2638_);
	assign _2640_ = (_4423_ ? _0957_ : _0757_);
	assign _2641_ = (_0127_ ? _0956_ : _2640_);
	assign _2642_ = (_4380_ ? _0577_ : _0425_);
	assign _2643_ = (_4423_ ? _0070_ : _2642_);
	assign _2644_ = (_4387_ ? _0255_ : _0495_);
	assign _2645_ = ~_2644_;
	assign _2646_ = (_0127_ ? _2643_ : _2645_);
	assign _2648_ = (_0146_ ? _2641_ : _2646_);
	assign _2649_ = (_4423_ ? _0903_ : _0153_);
	assign _2650_ = (_0056_ ? _0967_ : _2649_);
	assign _2651_ = (_0146_ ? _2650_ : _0973_);
	assign _2652_ = (\mchip.pong.game.vga.pix_ind [0] ? _2651_ : _2648_);
	assign _2653_ = (_0127_ ? _0567_ : _0986_);
	assign _2654_ = (_0146_ ? _2653_ : _0991_);
	assign _2655_ = (\mchip.pong.game.vga.pix_ind [0] ? _2654_ : _0984_);
	assign _2656_ = (_1103_ ? _2652_ : _2655_);
	assign _2657_ = (_0056_ ? _4389_ : _0996_);
	assign _2659_ = (_0146_ ? _2657_ : _1000_);
	assign _2660_ = (_4387_ ? _0852_ : _0530_);
	assign _2661_ = (_0127_ ? _1005_ : _2660_);
	assign _2662_ = (_0146_ ? _2661_ : _1013_);
	assign _2663_ = (\mchip.pong.game.vga.pix_ind [0] ? _2662_ : _2659_);
	assign _2664_ = (_4387_ ? _0117_ : _0119_);
	assign _2665_ = (_0127_ ? _0154_ : _2664_);
	assign _2666_ = (_4423_ ? _4371_ : _0606_);
	assign _2667_ = (_0056_ ? _1021_ : _2666_);
	assign _2668_ = (_0146_ ? _2665_ : _2667_);
	assign _2670_ = (_4423_ ? _0391_ : _0615_);
	assign _2671_ = (_0056_ ? _1031_ : _2670_);
	assign _2672_ = (_0146_ ? _1027_ : _2671_);
	assign _2673_ = (\mchip.pong.game.vga.pix_ind [0] ? _2672_ : _2668_);
	assign _2674_ = (_1103_ ? _2663_ : _2673_);
	assign _2675_ = (_0044_ ? _2656_ : _2674_);
	assign _2676_ = (_0088_ ? _2639_ : _2675_);
	assign _2677_ = (_4423_ ? _4389_ : _0070_);
	assign _2678_ = (_0127_ ? _1038_ : _2677_);
	assign _2679_ = (_0146_ ? _2678_ : _1042_);
	assign _2681_ = (_4387_ ? _0880_ : _0474_);
	assign _2682_ = (_0127_ ? _1044_ : _2681_);
	assign _2683_ = (_0146_ ? _2682_ : _1049_);
	assign _2684_ = (\mchip.pong.game.vga.pix_ind [0] ? _2683_ : _2679_);
	assign _2685_ = (_1103_ ? _0337_ : _2684_);
	assign _2686_ = (_0044_ ? _2685_ : _0329_);
	assign _2687_ = (_0088_ ? _2686_ : _0307_);
	assign _2688_ = (_4368_ ? _2676_ : _2687_);
	assign _2689_ = (_4367_ ? _2611_ : _2688_);
	assign _2690_ = (_1058_ ? _2689_ : _0347_);
	assign _2692_ = (_0723_ ? _2558_ : _2690_);
	assign _2693_ = (_1061_ ? _0347_ : _2692_);
	assign \mchip.pong.VGA_B2  = (_1264_ ? _2693_ : _1519_);
	assign _2694_ = _4417_ & _4387_;
	assign _2695_ = (_0056_ ? _2694_ : _0399_);
	assign _2696_ = (_0127_ ? _4429_ : _0420_);
	assign _2697_ = (_0146_ ? _2695_ : _2696_);
	assign _2698_ = _4428_ & ~_4387_;
	assign _2699_ = (_0127_ ? _0356_ : _2698_);
	assign _2700_ = (_4387_ ? _0203_ : _0035_);
	assign _2702_ = (_0127_ ? _1524_ : _2700_);
	assign _2703_ = (_0146_ ? _2699_ : _2702_);
	assign _2704_ = (\mchip.pong.game.vga.pix_ind [0] ? _2703_ : _2697_);
	assign _2705_ = _1590_ | _0135_;
	assign _2706_ = (_0056_ ? _2235_ : _1524_);
	assign _2707_ = (_0146_ ? _2705_ : _2706_);
	assign _2708_ = (_0127_ ? _4429_ : _1729_);
	assign _2709_ = (_0146_ ? _1727_ : _2708_);
	assign _2710_ = (\mchip.pong.game.vga.pix_ind [0] ? _2709_ : _2707_);
	assign _2711_ = (_1103_ ? _2704_ : _2710_);
	assign _2713_ = (_0044_ ? _1586_ : _2711_);
	assign _2714_ = (_0088_ ? _1568_ : _2713_);
	assign _2715_ = (_0127_ ? _0048_ : _1522_);
	assign _2716_ = (_4387_ ? _4428_ : _0153_);
	assign _2717_ = _2716_ | _0127_;
	assign _2718_ = (_0146_ ? _2715_ : _2717_);
	assign _2719_ = (_0127_ ? _0154_ : _1532_);
	assign _2720_ = _0442_ | _4423_;
	assign _2721_ = (_4387_ ? _0792_ : _4381_);
	assign _2722_ = (_0127_ ? _2720_ : _2721_);
	assign _2724_ = (_0146_ ? _2719_ : _2722_);
	assign _2725_ = (\mchip.pong.game.vga.pix_ind [0] ? _2724_ : _2718_);
	assign _2726_ = (_0127_ ? _0154_ : _2336_);
	assign _2727_ = _1652_ | _0156_;
	assign _2728_ = (_0146_ ? _2726_ : _2727_);
	assign _2729_ = (_0127_ ? _0399_ : _2336_);
	assign _2730_ = (_4423_ ? _2053_ : _0961_);
	assign _2731_ = _0056_ & ~_2730_;
	assign _2732_ = (_0146_ ? _2729_ : _2731_);
	assign _2733_ = (\mchip.pong.game.vga.pix_ind [0] ? _2732_ : _2728_);
	assign _2735_ = (_1103_ ? _2725_ : _2733_);
	assign _2736_ = (_4423_ ? _0117_ : _1908_);
	assign _2737_ = _2736_ | _0056_;
	assign _2738_ = (_0146_ ? _2737_ : _2060_);
	assign _2739_ = (_4423_ ? _4409_ : _0401_);
	assign _2740_ = _2739_ | _0127_;
	assign _2741_ = (_0146_ ? _1778_ : _2740_);
	assign _2742_ = (\mchip.pong.game.vga.pix_ind [0] ? _2741_ : _2738_);
	assign _2743_ = (_0056_ ? _0550_ : _1784_);
	assign _2744_ = (_4387_ ? _0203_ : _4409_);
	assign _2746_ = _2744_ | _0127_;
	assign _2747_ = (_0146_ ? _2743_ : _2746_);
	assign _2748_ = _0160_ | _0127_;
	assign _2749_ = (_0146_ ? _1740_ : _2748_);
	assign _2750_ = (\mchip.pong.game.vga.pix_ind [0] ? _2749_ : _2747_);
	assign _2751_ = (_1103_ ? _2742_ : _2750_);
	assign _2752_ = (_0044_ ? _2735_ : _2751_);
	assign _2753_ = _4387_ | _4381_;
	assign _2754_ = (_4387_ ? _0495_ : _2307_);
	assign _2755_ = (_0056_ ? _2753_ : _2754_);
	assign _2757_ = (_0146_ ? _2755_ : _0794_);
	assign _2758_ = (_4423_ ? _4381_ : _0451_);
	assign _2759_ = (_0127_ ? _1807_ : _2758_);
	assign _2760_ = (_0146_ ? _2759_ : _2082_);
	assign _2761_ = (\mchip.pong.game.vga.pix_ind [0] ? _2760_ : _2757_);
	assign _2762_ = (_4380_ ? _4372_ : _4407_);
	assign _2763_ = _2762_ | _4387_;
	assign _2764_ = (_0127_ ? _0619_ : _2763_);
	assign _2765_ = (_0146_ ? _2764_ : _2160_);
	assign _2766_ = (_0127_ ? _0619_ : _0872_);
	assign _2768_ = (_0146_ ? _2766_ : _2160_);
	assign _2769_ = (\mchip.pong.game.vga.pix_ind [0] ? _2768_ : _2765_);
	assign _2770_ = (_1103_ ? _2761_ : _2769_);
	assign _2771_ = (_4423_ ? _0118_ : _0495_);
	assign _2772_ = (_4380_ ? _4371_ : _0425_);
	assign _2773_ = (_4387_ ? _0475_ : _2772_);
	assign _2774_ = (_0127_ ? _2771_ : _2773_);
	assign _2775_ = (_0127_ ? _0572_ : _2105_);
	assign _2776_ = (_0146_ ? _2774_ : _2775_);
	assign _2777_ = (_4423_ ? _4371_ : _0207_);
	assign _2779_ = (_0127_ ? _2771_ : _2777_);
	assign _2780_ = (_0127_ ? _0550_ : _0793_);
	assign _2781_ = (_0146_ ? _2779_ : _2780_);
	assign _2782_ = (\mchip.pong.game.vga.pix_ind [0] ? _2781_ : _2776_);
	assign _2783_ = (_4423_ ? _0118_ : _0035_);
	assign _2784_ = (_4387_ ? _0119_ : _1846_);
	assign _2785_ = (_0127_ ? _2783_ : _2784_);
	assign _2786_ = (_0146_ ? _2785_ : _2780_);
	assign _2787_ = (_4423_ ? _4417_ : _0495_);
	assign _2788_ = (_0056_ ? _1857_ : _2787_);
	assign _2790_ = (_0127_ ? _0193_ : _0793_);
	assign _2791_ = (_0146_ ? _2788_ : _2790_);
	assign _2792_ = (\mchip.pong.game.vga.pix_ind [0] ? _2791_ : _2786_);
	assign _2793_ = (_1103_ ? _2782_ : _2792_);
	assign _2794_ = (_0044_ ? _2770_ : _2793_);
	assign _2795_ = (_0088_ ? _2752_ : _2794_);
	assign _2796_ = (_4368_ ? _2714_ : _2795_);
	assign _2797_ = (_4423_ ? _4389_ : _0361_);
	assign _2798_ = (_0056_ ? _1924_ : _2797_);
	assign _2799_ = _0635_ | _0127_;
	assign _2801_ = (_0146_ ? _2798_ : _2799_);
	assign _2802_ = (_0056_ ? _1879_ : _2105_);
	assign _2803_ = (_4387_ ? _4380_ : _0678_);
	assign _2804_ = _2803_ | _0127_;
	assign _2805_ = (_0146_ ? _2802_ : _2804_);
	assign _2806_ = (\mchip.pong.game.vga.pix_ind [0] ? _2805_ : _2801_);
	assign _2807_ = (_4423_ ? _0117_ : _0475_);
	assign _2808_ = (_0127_ ? _2105_ : _2807_);
	assign _2809_ = (_0127_ ? _0193_ : _2105_);
	assign _2810_ = (_0146_ ? _2808_ : _2809_);
	assign _2812_ = (_4423_ ? _4443_ : _0506_);
	assign _2813_ = (_4423_ ? _0852_ : _0475_);
	assign _2814_ = (_0127_ ? _2812_ : _2813_);
	assign _2815_ = (_0127_ ? _0550_ : _2105_);
	assign _2816_ = (_0146_ ? _2814_ : _2815_);
	assign _2817_ = (\mchip.pong.game.vga.pix_ind [0] ? _2816_ : _2810_);
	assign _2818_ = (_1103_ ? _2806_ : _2817_);
	assign _2819_ = (_4387_ ? _0054_ : _0852_);
	assign _2820_ = (_4389_ ? _4408_ : _4372_);
	assign _2821_ = (_4423_ ? _4389_ : _2820_);
	assign _2823_ = (_0127_ ? _2819_ : _2821_);
	assign _2824_ = _4387_ & ~_2307_;
	assign _2825_ = ~_2824_;
	assign _2826_ = (_0056_ ? _0834_ : _2825_);
	assign _2827_ = (_0146_ ? _2823_ : _2826_);
	assign _2828_ = (_4423_ ? _4389_ : _1908_);
	assign _2829_ = (_0056_ ? _2015_ : _2828_);
	assign _2830_ = (_4423_ ? _4409_ : _0583_);
	assign _2831_ = (_0127_ ? _1748_ : _2830_);
	assign _2832_ = (_0146_ ? _2829_ : _2831_);
	assign _2834_ = (\mchip.pong.game.vga.pix_ind [0] ? _2832_ : _2827_);
	assign _2835_ = (_4387_ ? _4380_ : _1028_);
	assign _2836_ = (_0127_ ? _0550_ : _2835_);
	assign _2837_ = (_0146_ ? _2829_ : _2836_);
	assign _2838_ = (_4423_ ? _4389_ : _2484_);
	assign _2839_ = (_0056_ ? _1924_ : _2838_);
	assign _2840_ = (_4387_ ? _0090_ : _4434_);
	assign _2841_ = (_0127_ ? _1888_ : _2840_);
	assign _2842_ = (_0146_ ? _2839_ : _2841_);
	assign _2843_ = (\mchip.pong.game.vga.pix_ind [0] ? _2842_ : _2837_);
	assign _2845_ = (_1103_ ? _2834_ : _2843_);
	assign _2846_ = (_0044_ ? _2818_ : _2845_);
	assign _2847_ = (_4423_ ? _0852_ : _0639_);
	assign _2848_ = (_0127_ ? _0697_ : _2847_);
	assign _2849_ = (_0146_ ? _2848_ : _1940_);
	assign _2850_ = (_4387_ ? _4409_ : _0391_);
	assign _2851_ = (_0127_ ? _2626_ : _2850_);
	assign _2852_ = (_4423_ ? _0792_ : _0426_);
	assign _2853_ = (_0056_ ? _0160_ : _2852_);
	assign _2854_ = (_0146_ ? _2851_ : _2853_);
	assign _2856_ = (\mchip.pong.game.vga.pix_ind [0] ? _2854_ : _2849_);
	assign _2857_ = _4387_ | ~_1853_;
	assign _2858_ = ~(_2857_ & _0095_);
	assign _2859_ = (_0127_ ? _2626_ : _2858_);
	assign _2860_ = (_4380_ ? _0065_ : _0756_);
	assign _2861_ = (_4423_ ? _0119_ : _2860_);
	assign _2862_ = (_0056_ ? _0160_ : _2861_);
	assign _2863_ = (_0146_ ? _2859_ : _2862_);
	assign _2864_ = (_4387_ ? _4381_ : _0852_);
	assign _2865_ = (_4423_ ? _0101_ : _2820_);
	assign _2867_ = (_0127_ ? _2864_ : _2865_);
	assign _2868_ = (_4371_ ? _4380_ : _0577_);
	assign _2869_ = _2868_ | _4423_;
	assign _2870_ = (_0056_ ? _1959_ : _2869_);
	assign _2871_ = (_0146_ ? _2867_ : _2870_);
	assign _2872_ = (\mchip.pong.game.vga.pix_ind [0] ? _2871_ : _2863_);
	assign _2873_ = (_1103_ ? _2856_ : _2872_);
	assign _2874_ = (_4387_ ? _4389_ : _0264_);
	assign _2875_ = (_0127_ ? _1965_ : _2874_);
	assign _2876_ = (_0146_ ? _2875_ : _1635_);
	assign _2878_ = (_4423_ ? _0107_ : _0372_);
	assign _2879_ = (_0127_ ? _4389_ : _2878_);
	assign _2880_ = (_0146_ ? _2879_ : _0135_);
	assign _2881_ = (\mchip.pong.game.vga.pix_ind [0] ? _2880_ : _2876_);
	assign _2882_ = (_0127_ ? _0702_ : _1574_);
	assign _2883_ = (_0146_ ? _2882_ : _0135_);
	assign _2884_ = (_0127_ ? _0697_ : _0323_);
	assign _2885_ = (_0146_ ? _2884_ : _1984_);
	assign _2886_ = (\mchip.pong.game.vga.pix_ind [0] ? _2885_ : _2883_);
	assign _2887_ = (_1103_ ? _2881_ : _2886_);
	assign _2889_ = (_0044_ ? _2873_ : _2887_);
	assign _2890_ = (_0088_ ? _2846_ : _2889_);
	assign _2891_ = (_4368_ ? _2890_ : _1997_);
	assign _2892_ = (_4367_ ? _2796_ : _2891_);
	assign _2893_ = (_4387_ ? _4381_ : _0703_);
	assign _2894_ = (_0056_ ? _0501_ : _2893_);
	assign _2895_ = (_0146_ ? _2894_ : _2033_);
	assign _2896_ = (\mchip.pong.game.vga.pix_ind [0] ? _2040_ : _2895_);
	assign _2897_ = (_1103_ ? _2896_ : _2051_);
	assign _2898_ = ~_2070_;
	assign _2900_ = ~_2071_;
	assign _2901_ = (_0146_ ? _2898_ : _2900_);
	assign _2902_ = _2626_ | _0056_;
	assign _2903_ = (_0146_ ? _2902_ : _2060_);
	assign _2904_ = (\mchip.pong.game.vga.pix_ind [0] ? _2901_ : _2903_);
	assign _2905_ = (_1103_ ? _2062_ : _2904_);
	assign _2906_ = (_0044_ ? _2897_ : _2905_);
	assign _2907_ = (_4423_ ? _0451_ : _0254_);
	assign _2908_ = (_0127_ ? _2105_ : _2907_);
	assign _2909_ = (_0146_ ? _2908_ : _2082_);
	assign _2910_ = (\mchip.pong.game.vga.pix_ind [0] ? _2114_ : _2909_);
	assign _2911_ = (_1103_ ? _2910_ : _2117_);
	assign _2912_ = (_0044_ ? _2104_ : _2911_);
	assign _2913_ = (_0088_ ? _2906_ : _2912_);
	assign _2914_ = (_4368_ ? _2027_ : _2913_);
	assign _2915_ = (_4387_ ? _0035_ : _0579_);
	assign _2916_ = _2915_ | _0056_;
	assign _2917_ = (_0146_ ? _2916_ : _2139_);
	assign _2918_ = (\mchip.pong.game.vga.pix_ind [0] ? _2917_ : _2136_);
	assign _2919_ = (_1103_ ? _2131_ : _2918_);
	assign _2921_ = (_4387_ ? _0054_ : _2278_);
	assign _2922_ = (_0056_ ? _2145_ : _2921_);
	assign _2923_ = (_0146_ ? _2922_ : _2147_);
	assign _2924_ = (_4387_ ? _0054_ : _1903_);
	assign _2925_ = (_0056_ ? _2145_ : _2924_);
	assign _2926_ = (_0146_ ? _2925_ : _2057_);
	assign _2927_ = (\mchip.pong.game.vga.pix_ind [0] ? _2926_ : _2923_);
	assign _2928_ = (_1103_ ? _2927_ : _2162_);
	assign _2929_ = (_0044_ ? _2919_ : _2928_);
	assign _2930_ = _4380_ | ~_4433_;
	assign _2932_ = (_4423_ ? _0421_ : _2930_);
	assign _2933_ = (_0127_ ? _0154_ : _2932_);
	assign _2934_ = _0264_ | ~_4387_;
	assign _2935_ = (_0056_ ? _0972_ : _2934_);
	assign _2936_ = (_0146_ ? _2933_ : _2935_);
	assign _2937_ = (_0056_ ? _0140_ : _2064_);
	assign _2938_ = (_0146_ ? _2937_ : _2174_);
	assign _2939_ = (\mchip.pong.game.vga.pix_ind [0] ? _2938_ : _2936_);
	assign _2940_ = (_4387_ ? _4381_ : _4437_);
	assign _2941_ = (_0056_ ? _2145_ : _2940_);
	assign _2943_ = (_0146_ ? _2941_ : _2184_);
	assign _2944_ = (\mchip.pong.game.vga.pix_ind [0] ? _2943_ : _2181_);
	assign _2945_ = (_1103_ ? _2939_ : _2944_);
	assign _2946_ = (_0056_ ? _0592_ : _1976_);
	assign _2947_ = (_4423_ ? _0444_ : _2361_);
	assign _2948_ = (_0056_ ? _2209_ : _2947_);
	assign _2949_ = (_0146_ ? _2946_ : _2948_);
	assign _2950_ = (\mchip.pong.game.vga.pix_ind [0] ? _2218_ : _2949_);
	assign _2951_ = (_1103_ ? _2207_ : _2950_);
	assign _2952_ = (_0044_ ? _2945_ : _2951_);
	assign _2954_ = (_0088_ ? _2929_ : _2952_);
	assign _2955_ = (_4368_ ? _2954_ : _2242_);
	assign _2956_ = (_4367_ ? _2914_ : _2955_);
	assign _2957_ = (_1058_ ? _2956_ : _1706_);
	assign _2958_ = (_0723_ ? _2892_ : _2957_);
	assign _2959_ = (_1061_ ? _1706_ : _2958_);
	assign \mchip.pong.VGA_B3  = (_1264_ ? _2959_ : _1519_);
	assign _2960_ = (_1103_ ? _0061_ : _0081_);
	assign _2961_ = _1103_ & ~_4432_;
	assign _2962_ = (\mchip.pong.game.vga.pix_ind [0] ? _4440_ : _0039_);
	assign _2964_ = _2962_ & ~_1103_;
	assign _2965_ = _2964_ | _2961_;
	assign _2966_ = (_0044_ ? _2965_ : _2960_);
	assign _2967_ = _0044_ & ~_0124_;
	assign _2968_ = _0308_ & ~_0149_;
	assign _2969_ = _2968_ | _2967_;
	assign _2970_ = (_0088_ ? _2966_ : _2969_);
	assign _2971_ = _0088_ & ~_0186_;
	assign _2972_ = _0214_ & ~_0088_;
	assign _2973_ = _2972_ | _2971_;
	assign _2975_ = (_4368_ ? _2970_ : _2973_);
	assign _2976_ = _0088_ | ~_0307_;
	assign _2977_ = _0344_ & ~_0152_;
	assign _2978_ = _2976_ & ~_2977_;
	assign _2979_ = ~(_0241_ & _0044_);
	assign _2980_ = _0249_ & ~_0044_;
	assign _2981_ = _2979_ & ~_2980_;
	assign _2982_ = _0220_ & _0044_;
	assign _2983_ = _0308_ & ~_0230_;
	assign _2984_ = _2983_ | _2982_;
	assign _2986_ = (_0088_ ? _2984_ : _2981_);
	assign _2987_ = (_4368_ ? _2986_ : _2978_);
	assign _2988_ = (_4367_ ? _2975_ : _2987_);
	assign _2989_ = _1103_ | ~_0106_;
	assign _2990_ = ~(_2820_ & _4423_);
	assign _2991_ = (_0056_ ? _0115_ : _2990_);
	assign _2992_ = (_0146_ ? _0348_ : _2991_);
	assign _2993_ = ~_0109_;
	assign _2994_ = ~_0111_;
	assign _2995_ = (_0146_ ? _2993_ : _2994_);
	assign _2997_ = (\mchip.pong.game.vga.pix_ind [0] ? _2995_ : _2992_);
	assign _2998_ = _1103_ & ~_2997_;
	assign _2999_ = _2989_ & ~_2998_;
	assign _3000_ = (_4423_ ? _0295_ : _0119_);
	assign _3001_ = (_0127_ ? _0128_ : _3000_);
	assign _3002_ = ~(_0530_ & _4387_);
	assign _3003_ = (_4387_ ? _4391_ : _0117_);
	assign _3004_ = (_0127_ ? _3002_ : _3003_);
	assign _3005_ = (_0146_ ? _3001_ : _3004_);
	assign _3006_ = (_4387_ ? _0107_ : _1832_);
	assign _3008_ = (_0127_ ? _0132_ : _3006_);
	assign _3009_ = ~_0606_;
	assign _3010_ = (_4423_ ? _0703_ : _3009_);
	assign _3011_ = (_4387_ ? _0295_ : _2053_);
	assign _3012_ = (_0127_ ? _3010_ : _3011_);
	assign _3013_ = (_0146_ ? _3008_ : _3012_);
	assign _3014_ = (\mchip.pong.game.vga.pix_ind [0] ? _3013_ : _3005_);
	assign _3015_ = (_0056_ ? _0091_ : _0138_);
	assign _3016_ = (_4387_ ? _0281_ : _0792_);
	assign _3017_ = (_0056_ ? _0140_ : _3016_);
	assign _3019_ = (_0146_ ? _3015_ : _3017_);
	assign _3020_ = (_0056_ ? _0350_ : _0143_);
	assign _3021_ = (_4423_ ? _0495_ : _0521_);
	assign _3022_ = (_0056_ ? _0120_ : _3021_);
	assign _3023_ = (_0146_ ? _3020_ : _3022_);
	assign _3024_ = (\mchip.pong.game.vga.pix_ind [0] ? _3023_ : _3019_);
	assign _3025_ = (_1103_ ? _3014_ : _3024_);
	assign _3026_ = (_0044_ ? _2999_ : _3025_);
	assign _3027_ = (_0088_ ? _2966_ : _3026_);
	assign _3028_ = (_0127_ ? _1798_ : _1560_);
	assign _3030_ = (_4423_ ? _4381_ : _1927_);
	assign _3031_ = _0056_ & ~_3030_;
	assign _3032_ = (_0146_ ? _3028_ : _3031_);
	assign _3033_ = (_0056_ ? _0549_ : _0162_);
	assign _3034_ = _4387_ & ~_2860_;
	assign _3035_ = (_4423_ ? _0495_ : _1009_);
	assign _3036_ = (_0127_ ? _3034_ : _3035_);
	assign _3037_ = (_0146_ ? _3033_ : _3036_);
	assign _3038_ = (\mchip.pong.game.vga.pix_ind [0] ? _3037_ : _3032_);
	assign _3039_ = (_4387_ ? _0113_ : _0850_);
	assign _3041_ = (_0127_ ? _0166_ : _3039_);
	assign _3042_ = (_4387_ ? _4389_ : _1808_);
	assign _3043_ = (_4423_ ? _2053_ : _0281_);
	assign _3044_ = (_0127_ ? _3042_ : _3043_);
	assign _3045_ = (_0146_ ? _3041_ : _3044_);
	assign _3046_ = (_4389_ ? _4374_ : _4427_);
	assign _3047_ = (_4387_ ? _0119_ : _3046_);
	assign _3048_ = (_0127_ ? _1798_ : _3047_);
	assign _3049_ = (_4387_ ? _0035_ : _0521_);
	assign _3050_ = _1612_ & _0098_;
	assign _3052_ = (_0127_ ? _3049_ : _3050_);
	assign _3053_ = (_0146_ ? _3048_ : _3052_);
	assign _3054_ = (\mchip.pong.game.vga.pix_ind [0] ? _3053_ : _3045_);
	assign _3055_ = (_1103_ ? _3038_ : _3054_);
	assign _3056_ = (_4387_ ? _0826_ : _0530_);
	assign _3057_ = _0127_ & ~_3056_;
	assign _3058_ = (_4423_ ? _4443_ : _2307_);
	assign _3059_ = _0056_ & ~_3058_;
	assign _3060_ = (_0146_ ? _3057_ : _3059_);
	assign _3061_ = ~_0410_;
	assign _3063_ = (_0276_ ? _3061_ : _0443_);
	assign _3064_ = (_0056_ ? _0875_ : _3063_);
	assign _3065_ = (_4423_ ? _0153_ : _0391_);
	assign _3066_ = _0056_ & ~_3065_;
	assign _3067_ = (_0146_ ? _3064_ : _3066_);
	assign _3068_ = (\mchip.pong.game.vga.pix_ind [0] ? _3067_ : _3060_);
	assign _3069_ = (_0127_ ? _0055_ : _0447_);
	assign _3070_ = (_4423_ ? _0153_ : _1028_);
	assign _3071_ = _0056_ & ~_3070_;
	assign _3072_ = (_0146_ ? _3069_ : _3071_);
	assign _3074_ = ~_0179_;
	assign _3075_ = _4387_ & ~_0880_;
	assign _3076_ = (_0127_ ? _3074_ : _3075_);
	assign _3077_ = (_4423_ ? _4409_ : _0623_);
	assign _3078_ = ~(_3077_ | _0127_);
	assign _3079_ = (_0146_ ? _3076_ : _3078_);
	assign _3080_ = (\mchip.pong.game.vga.pix_ind [0] ? _3079_ : _3072_);
	assign _3081_ = (_1103_ ? _3068_ : _3080_);
	assign _3082_ = (_0044_ ? _3055_ : _3081_);
	assign _3083_ = ~(_1809_ | _4387_);
	assign _3085_ = (_0127_ ? _0618_ : _3083_);
	assign _3086_ = (_4423_ ? _1002_ : _1903_);
	assign _3087_ = (_0127_ ? _0754_ : _3086_);
	assign _3088_ = (_0146_ ? _3085_ : _3087_);
	assign _3089_ = (_4387_ ? _0450_ : _0410_);
	assign _3090_ = (_0127_ ? _2137_ : _3089_);
	assign _3091_ = (_4423_ ? _0490_ : _2307_);
	assign _3092_ = _0056_ & ~_3091_;
	assign _3093_ = (_0146_ ? _3090_ : _3092_);
	assign _3094_ = (\mchip.pong.game.vga.pix_ind [0] ? _3093_ : _3088_);
	assign _3096_ = (_4423_ ? _4389_ : _2307_);
	assign _3097_ = _0056_ & ~_3096_;
	assign _3098_ = (_0146_ ? _0155_ : _3097_);
	assign _3099_ = (_1103_ ? _3094_ : _3098_);
	assign _3100_ = (_4389_ ? _4372_ : _4419_);
	assign _3101_ = _4387_ & ~_3100_;
	assign _3102_ = (_4423_ ? _0454_ : _0882_);
	assign _3103_ = (_0127_ ? _3101_ : _3102_);
	assign _3104_ = _4387_ & ~_0579_;
	assign _3105_ = (_4412_ ? _0367_ : _0207_);
	assign _3107_ = (_0127_ ? _3104_ : _3105_);
	assign _3108_ = (_0146_ ? _3103_ : _3107_);
	assign _3109_ = (_0056_ ? _0452_ : _3101_);
	assign _3110_ = (_4387_ ? _2256_ : _1809_);
	assign _3111_ = (_0127_ ? _0591_ : _3110_);
	assign _3112_ = (_0146_ ? _3109_ : _3111_);
	assign _3113_ = (\mchip.pong.game.vga.pix_ind [0] ? _3112_ : _3108_);
	assign _3114_ = (_4387_ ? _0450_ : _0263_);
	assign _3115_ = (_0127_ ? _0618_ : _3114_);
	assign _3116_ = ~_0045_;
	assign _3118_ = (_4387_ ? _0153_ : _3116_);
	assign _3119_ = (_0127_ ? _1841_ : _3118_);
	assign _3120_ = (_0146_ ? _3115_ : _3119_);
	assign _3121_ = (_0276_ ? _0371_ : _0450_);
	assign _3122_ = (_0127_ ? _0618_ : _3121_);
	assign _3123_ = (_4387_ ? _1903_ : _1809_);
	assign _3124_ = _3123_ & ~_0127_;
	assign _3125_ = (_0146_ ? _3122_ : _3124_);
	assign _3126_ = (\mchip.pong.game.vga.pix_ind [0] ? _3125_ : _3120_);
	assign _3127_ = (_1103_ ? _3113_ : _3126_);
	assign _3129_ = (_0044_ ? _3099_ : _3127_);
	assign _3130_ = (_0088_ ? _3082_ : _3129_);
	assign _3131_ = (_4368_ ? _3027_ : _3130_);
	assign _3132_ = (_4423_ ? _0292_ : _4424_);
	assign _3133_ = (_0127_ ? _0399_ : _3132_);
	assign _3134_ = (_4387_ ? _0090_ : _0613_);
	assign _3135_ = _0056_ & ~_3134_;
	assign _3136_ = (_0146_ ? _3133_ : _3135_);
	assign _3137_ = ~_2807_;
	assign _3138_ = _4387_ & ~_1908_;
	assign _3140_ = (_0056_ ? _3137_ : _3138_);
	assign _3141_ = _0056_ & ~_2835_;
	assign _3142_ = (_0146_ ? _3140_ : _3141_);
	assign _3143_ = (\mchip.pong.game.vga.pix_ind [0] ? _3142_ : _3136_);
	assign _3144_ = (_4387_ ? _0100_ : _0529_);
	assign _3145_ = (_0127_ ? _0618_ : _3144_);
	assign _3146_ = _4387_ & ~_0101_;
	assign _3147_ = (_4387_ ? _4389_ : _0207_);
	assign _3148_ = (_0127_ ? _3146_ : _3147_);
	assign _3149_ = (_0146_ ? _3145_ : _3148_);
	assign _3151_ = _4423_ & ~_0530_;
	assign _3152_ = (_0127_ ? _0618_ : _3151_);
	assign _3153_ = (_4389_ ? _0425_ : _4433_);
	assign _3154_ = (_4387_ ? _4389_ : _3153_);
	assign _3155_ = (_0127_ ? _1555_ : _3154_);
	assign _3156_ = (_0146_ ? _3152_ : _3155_);
	assign _3157_ = (\mchip.pong.game.vga.pix_ind [0] ? _3156_ : _3149_);
	assign _3158_ = (_1103_ ? _3143_ : _3157_);
	assign _3159_ = (_4387_ ? _0598_ : _4437_);
	assign _3160_ = _4437_ | _4387_;
	assign _3162_ = _0631_ & ~_4423_;
	assign _3163_ = _3160_ & ~_3162_;
	assign _3164_ = (_0127_ ? _3159_ : _3163_);
	assign _3165_ = ~_0609_;
	assign _3166_ = _4387_ & ~_0756_;
	assign _3167_ = (_0056_ ? _3165_ : _3166_);
	assign _3168_ = (_0146_ ? _3164_ : _3167_);
	assign _3169_ = (_4437_ ? _4423_ : _4387_);
	assign _3170_ = _4423_ | ~_0639_;
	assign _3171_ = _0530_ & ~_4387_;
	assign _3173_ = _3170_ & ~_3171_;
	assign _3174_ = (_0127_ ? _3169_ : _3173_);
	assign _3175_ = (_4387_ ? _4372_ : _0621_);
	assign _3176_ = (_0127_ ? _1747_ : _3175_);
	assign _3177_ = (_0146_ ? _3174_ : _3176_);
	assign _3178_ = (\mchip.pong.game.vga.pix_ind [0] ? _3177_ : _3168_);
	assign _3179_ = (_0056_ ? _0828_ : _1877_);
	assign _3180_ = ~_0572_;
	assign _3181_ = (_4423_ ? _0113_ : _0882_);
	assign _3182_ = (_0127_ ? _3180_ : _3181_);
	assign _3184_ = (_0146_ ? _3179_ : _3182_);
	assign _3185_ = _4387_ & ~_0314_;
	assign _3186_ = (_0127_ ? _0154_ : _3185_);
	assign _3187_ = (_4387_ ? _0089_ : _0654_);
	assign _3188_ = (_0127_ ? _0531_ : _3187_);
	assign _3189_ = (_0146_ ? _3186_ : _3188_);
	assign _3190_ = (\mchip.pong.game.vga.pix_ind [0] ? _3189_ : _3184_);
	assign _3191_ = (_1103_ ? _3178_ : _3190_);
	assign _3192_ = (_0044_ ? _3158_ : _3191_);
	assign _3193_ = (_4423_ ? _0292_ : _0391_);
	assign _3195_ = (_0056_ ? _3151_ : _3193_);
	assign _3196_ = ~_0160_;
	assign _3197_ = (_0127_ ? _0103_ : _3196_);
	assign _3198_ = (_0146_ ? _3195_ : _3197_);
	assign _3199_ = (_0056_ ? _1837_ : _1934_);
	assign _3200_ = (_4423_ ? _0101_ : _0371_);
	assign _3201_ = (_0056_ ? _0098_ : _3200_);
	assign _3202_ = (_0146_ ? _3199_ : _3201_);
	assign _3203_ = (\mchip.pong.game.vga.pix_ind [0] ? _3202_ : _3198_);
	assign _3204_ = ~_0976_;
	assign _3206_ = (_4387_ ? _0839_ : _1852_);
	assign _3207_ = (_0127_ ? _3204_ : _3206_);
	assign _3208_ = (_4423_ ? _0450_ : _0206_);
	assign _3209_ = (_0056_ ? _0181_ : _3208_);
	assign _3210_ = (_0146_ ? _3207_ : _3209_);
	assign _3211_ = ~(_0093_ & _4423_);
	assign _3212_ = _3211_ & ~_3162_;
	assign _3213_ = (_0127_ ? _2054_ : _3212_);
	assign _3214_ = _4387_ & ~_0065_;
	assign _3215_ = (_0056_ ? _0237_ : _3214_);
	assign _3217_ = (_0146_ ? _3213_ : _3215_);
	assign _3218_ = (\mchip.pong.game.vga.pix_ind [0] ? _3217_ : _3210_);
	assign _3219_ = (_1103_ ? _3203_ : _3218_);
	assign _3220_ = ~_0242_;
	assign _3221_ = ~(_0689_ & _0056_);
	assign _3222_ = (_4387_ ? _0970_ : _0529_);
	assign _3223_ = _0127_ & ~_3222_;
	assign _3224_ = _3221_ & ~_3223_;
	assign _3225_ = (_0146_ ? _3224_ : _3220_);
	assign _3226_ = ~_0126_;
	assign _3228_ = (_4423_ ? _0035_ : _1002_);
	assign _3229_ = (_4387_ ? _0529_ : _4417_);
	assign _3230_ = (_0127_ ? _3228_ : _3229_);
	assign _3231_ = (_0146_ ? _3230_ : _3226_);
	assign _3232_ = (\mchip.pong.game.vga.pix_ind [0] ? _3231_ : _3225_);
	assign _3233_ = (_0056_ ? _1817_ : _1934_);
	assign _3234_ = (_0127_ ? _0052_ : _0098_);
	assign _3235_ = (_0146_ ? _3233_ : _3234_);
	assign _3236_ = ~_0706_;
	assign _3237_ = ~_0140_;
	assign _3239_ = (_4423_ ? _0292_ : _4410_);
	assign _3240_ = (_0056_ ? _3237_ : _3239_);
	assign _3241_ = (_0159_ ? _3236_ : _3240_);
	assign _3242_ = (\mchip.pong.game.vga.pix_ind [0] ? _3241_ : _3235_);
	assign _3243_ = (_1103_ ? _3232_ : _3242_);
	assign _3244_ = (_0044_ ? _3219_ : _3243_);
	assign _3245_ = (_0088_ ? _3192_ : _3244_);
	assign _3246_ = _3245_ & _4368_;
	assign _3247_ = ~(_0719_ | _4368_);
	assign _3248_ = _3247_ | _3246_;
	assign _3250_ = (_4367_ ? _3131_ : _3248_);
	assign _3251_ = (_0146_ ? _0724_ : _2003_);
	assign _3252_ = _0056_ & ~_0778_;
	assign _3253_ = (_0146_ ? _0731_ : _3252_);
	assign _3254_ = (\mchip.pong.game.vga.pix_ind [0] ? _3253_ : _3251_);
	assign _3255_ = ~_0744_;
	assign _3256_ = (_4387_ ? _4408_ : _0292_);
	assign _3257_ = (_4387_ ? _0117_ : _0114_);
	assign _3258_ = (_0127_ ? _3256_ : _3257_);
	assign _3259_ = (_0146_ ? _3255_ : _3258_);
	assign _3261_ = (\mchip.pong.game.vga.pix_ind [0] ? _0740_ : _3259_);
	assign _3262_ = (_1103_ ? _3254_ : _3261_);
	assign _3263_ = _3262_ & ~_0044_;
	assign _3264_ = _3263_ | _2967_;
	assign _3265_ = (_0088_ ? _2966_ : _3264_);
	assign _3266_ = _0044_ | ~_0814_;
	assign _3267_ = (_4387_ ? _0495_ : _0506_);
	assign _3268_ = (_0056_ ? _0754_ : _3267_);
	assign _3269_ = (_4387_ ? _4389_ : _2338_);
	assign _3270_ = (_0056_ ? _0761_ : _3269_);
	assign _3272_ = (_0146_ ? _3268_ : _3270_);
	assign _3273_ = (_4387_ ? _4380_ : _0450_);
	assign _3274_ = (_4387_ ? _0117_ : _0495_);
	assign _3275_ = (_0127_ ? _3273_ : _3274_);
	assign _3276_ = (_0146_ ? _0767_ : _3275_);
	assign _3277_ = (\mchip.pong.game.vga.pix_ind [0] ? _3276_ : _3272_);
	assign _3278_ = _0056_ & ~_0374_;
	assign _3279_ = (_0146_ ? _0774_ : _3278_);
	assign _3280_ = (_4387_ ? _0412_ : _4381_);
	assign _3281_ = _0056_ & ~_3280_;
	assign _3283_ = (_0146_ ? _0781_ : _3281_);
	assign _3284_ = (\mchip.pong.game.vga.pix_ind [0] ? _3283_ : _3279_);
	assign _3285_ = (_1103_ ? _3277_ : _3284_);
	assign _3286_ = _0044_ & ~_3285_;
	assign _3287_ = _3266_ & ~_3286_;
	assign _3288_ = _0146_ | ~_0824_;
	assign _3289_ = _4408_ | _4387_;
	assign _3290_ = (_4387_ ? _0054_ : _0826_);
	assign _3291_ = (_0056_ ? _3289_ : _3290_);
	assign _3292_ = _3291_ & ~_0159_;
	assign _3294_ = _3288_ & ~_3292_;
	assign _3295_ = ~_0834_;
	assign _3296_ = (_0127_ ? _0832_ : _3295_);
	assign _3297_ = _0127_ & ~_0827_;
	assign _3298_ = (_0146_ ? _3297_ : _3296_);
	assign _3299_ = (\mchip.pong.game.vga.pix_ind [0] ? _3298_ : _3294_);
	assign _3300_ = _0127_ & ~_0838_;
	assign _3301_ = ~_0846_;
	assign _3302_ = (_4423_ ? _0665_ : _1903_);
	assign _3303_ = (_0056_ ? _3301_ : _3302_);
	assign _3305_ = (_0146_ ? _3300_ : _3303_);
	assign _3306_ = _0127_ & ~_0849_;
	assign _3307_ = (_4387_ ? _0131_ : _0529_);
	assign _3308_ = _3307_ & ~_0127_;
	assign _3309_ = _3308_ | _3306_;
	assign _3310_ = ~_0856_;
	assign _3311_ = (_4389_ ? _0065_ : _4427_);
	assign _3312_ = (_4423_ ? _0292_ : _3311_);
	assign _3313_ = (_0056_ ? _3310_ : _3312_);
	assign _3314_ = (_0146_ ? _3309_ : _3313_);
	assign _3316_ = (\mchip.pong.game.vga.pix_ind [0] ? _3314_ : _3305_);
	assign _3317_ = (_1103_ ? _3299_ : _3316_);
	assign _3318_ = (_4387_ ? _0295_ : _0113_);
	assign _3319_ = ~(_2387_ | _2362_);
	assign _3320_ = (_0127_ ? _3318_ : _3319_);
	assign _3321_ = ~_0867_;
	assign _3322_ = (_0056_ ? _3321_ : _3075_);
	assign _3323_ = (_0146_ ? _3320_ : _3322_);
	assign _3324_ = (_0127_ ? _0875_ : _3321_);
	assign _3325_ = _4423_ & ~_2361_;
	assign _3327_ = (_0127_ ? _0738_ : _3325_);
	assign _3328_ = (_0146_ ? _3327_ : _3324_);
	assign _3329_ = (\mchip.pong.game.vga.pix_ind [0] ? _3328_ : _3323_);
	assign _3330_ = (_0127_ ? _0500_ : _3321_);
	assign _3331_ = (_4387_ ? _2053_ : _0119_);
	assign _3332_ = (_0056_ ? _3325_ : _3331_);
	assign _3333_ = (_0146_ ? _3332_ : _3330_);
	assign _3334_ = ~_0894_;
	assign _3335_ = ~_0536_;
	assign _3336_ = (_0056_ ? _0452_ : _3335_);
	assign _3338_ = (_0159_ ? _3334_ : _3336_);
	assign _3339_ = (\mchip.pong.game.vga.pix_ind [0] ? _3338_ : _3333_);
	assign _3340_ = (_1103_ ? _3329_ : _3339_);
	assign _3341_ = (_0044_ ? _3317_ : _3340_);
	assign _3342_ = (_0088_ ? _3287_ : _3341_);
	assign _3343_ = (_4368_ ? _3265_ : _3342_);
	assign _3344_ = _4423_ & ~_0372_;
	assign _3345_ = (_0127_ ? _0502_ : _3344_);
	assign _3346_ = (_0127_ ? _0727_ : _3295_);
	assign _3347_ = (_0146_ ? _3345_ : _3346_);
	assign _3349_ = (_0127_ ? _0549_ : _3295_);
	assign _3350_ = (_4423_ ? _4380_ : _2053_);
	assign _3351_ = (_0056_ ? _1817_ : _3350_);
	assign _3352_ = (_0159_ ? _3349_ : _3351_);
	assign _3353_ = (\mchip.pong.game.vga.pix_ind [0] ? _3352_ : _3347_);
	assign _3354_ = _0127_ & ~_0816_;
	assign _3355_ = _4387_ & ~_0401_;
	assign _3356_ = _0350_ & ~_3355_;
	assign _3357_ = (_0056_ ? _3321_ : _3356_);
	assign _3358_ = (_0146_ ? _3354_ : _3357_);
	assign _3360_ = (_4387_ ? _0054_ : _0579_);
	assign _3361_ = _0127_ & ~_3360_;
	assign _3362_ = (_4423_ ? _0292_ : _0118_);
	assign _3363_ = (_0056_ ? _3321_ : _3362_);
	assign _3364_ = (_0146_ ? _3361_ : _3363_);
	assign _3365_ = (\mchip.pong.game.vga.pix_ind [0] ? _3364_ : _3358_);
	assign _3366_ = (_1103_ ? _3353_ : _3365_);
	assign _3367_ = ~_0924_;
	assign _3368_ = _4437_ & _4423_;
	assign _3369_ = (_0127_ ? _3367_ : _3368_);
	assign _3371_ = ~_0929_;
	assign _3372_ = (_0056_ ? _3371_ : _2824_);
	assign _3373_ = (_0146_ ? _3369_ : _3372_);
	assign _3374_ = ~_0823_;
	assign _3375_ = (_0127_ ? _0549_ : _3374_);
	assign _3376_ = _0127_ & ~_0932_;
	assign _3377_ = (_0159_ ? _3375_ : _3376_);
	assign _3378_ = (\mchip.pong.game.vga.pix_ind [0] ? _3377_ : _3373_);
	assign _3379_ = (_0146_ ? _2132_ : _0943_);
	assign _3380_ = (_0159_ ? _0950_ : _3306_);
	assign _3382_ = (\mchip.pong.game.vga.pix_ind [0] ? _3380_ : _3379_);
	assign _3383_ = (_1103_ ? _3378_ : _3382_);
	assign _3384_ = (_0044_ ? _3366_ : _3383_);
	assign _3385_ = ~_0956_;
	assign _3386_ = (_4387_ ? _0539_ : _0474_);
	assign _3387_ = (_0127_ ? _3385_ : _3386_);
	assign _3388_ = (_4423_ ? _4413_ : _0094_);
	assign _3389_ = (_0056_ ? _2644_ : _3388_);
	assign _3390_ = (_0146_ ? _3387_ : _3389_);
	assign _3391_ = (_4387_ ? _0792_ : _0371_);
	assign _3393_ = (_4423_ ? _0871_ : _0495_);
	assign _3394_ = (_0127_ ? _3393_ : _3391_);
	assign _3395_ = ~_0972_;
	assign _3396_ = (_0056_ ? _3395_ : _1557_);
	assign _3397_ = (_0146_ ? _3394_ : _3396_);
	assign _3398_ = (\mchip.pong.game.vga.pix_ind [0] ? _3397_ : _3390_);
	assign _3399_ = (_4423_ ? _4389_ : _0665_);
	assign _3400_ = _0127_ & ~_3399_;
	assign _3401_ = ~_0981_;
	assign _3402_ = (_4423_ ? _0292_ : _0281_);
	assign _3404_ = (_0056_ ? _3401_ : _3402_);
	assign _3405_ = (_0146_ ? _3400_ : _3404_);
	assign _3406_ = _0146_ | ~_0991_;
	assign _3407_ = _0146_ & ~_3361_;
	assign _3408_ = _3406_ & ~_3407_;
	assign _3409_ = (\mchip.pong.game.vga.pix_ind [0] ? _3408_ : _3405_);
	assign _3410_ = (_1103_ ? _3398_ : _3409_);
	assign _3411_ = ~_0996_;
	assign _3412_ = (_0056_ ? _0549_ : _3411_);
	assign _3413_ = (_4387_ ? _0206_ : _0417_);
	assign _3415_ = (_4423_ ? _4389_ : _2256_);
	assign _3416_ = (_0127_ ? _3413_ : _3415_);
	assign _3417_ = (_0146_ ? _3412_ : _3416_);
	assign _3418_ = (_0276_ ? _0474_ : _0850_);
	assign _3419_ = (_0127_ ? _1003_ : _3418_);
	assign _3420_ = ~_2001_;
	assign _3421_ = _0852_ & _4387_;
	assign _3422_ = _3211_ & ~_3421_;
	assign _3423_ = (_0056_ ? _3420_ : _3422_);
	assign _3424_ = (_0146_ ? _3419_ : _3423_);
	assign _3426_ = (\mchip.pong.game.vga.pix_ind [0] ? _3424_ : _3417_);
	assign _3427_ = (_4387_ ? _4380_ : _0474_);
	assign _3428_ = (_0127_ ? _1798_ : _3427_);
	assign _3429_ = (_4423_ ? _0454_ : _0412_);
	assign _3430_ = (_0056_ ? _1756_ : _3429_);
	assign _3431_ = (_0146_ ? _3428_ : _3430_);
	assign _3432_ = ~_1025_;
	assign _3433_ = (_4387_ ? _0035_ : _0100_);
	assign _3434_ = (_0127_ ? _3432_ : _3433_);
	assign _3435_ = (_4389_ ? _4433_ : _4372_);
	assign _3437_ = (_4387_ ? _0489_ : _3435_);
	assign _3438_ = (_4389_ ? _4427_ : _0259_);
	assign _3439_ = (_4423_ ? _2053_ : _3438_);
	assign _3440_ = (_0127_ ? _3437_ : _3439_);
	assign _3441_ = (_0146_ ? _3434_ : _3440_);
	assign _3442_ = (\mchip.pong.game.vga.pix_ind [0] ? _3441_ : _3431_);
	assign _3443_ = (_1103_ ? _3426_ : _3442_);
	assign _3444_ = (_0044_ ? _3410_ : _3443_);
	assign _3445_ = (_0088_ ? _3384_ : _3444_);
	assign _3446_ = _0330_ | _0056_;
	assign _3448_ = ~_0332_;
	assign _3449_ = (_0146_ ? _3446_ : _3448_);
	assign _3450_ = ~_0116_;
	assign _3451_ = ~_0335_;
	assign _3452_ = (_0146_ ? _3451_ : _3450_);
	assign _3453_ = (\mchip.pong.game.vga.pix_ind [0] ? _3452_ : _3449_);
	assign _3454_ = ~_1041_;
	assign _3455_ = (_0056_ ? _0143_ : _3454_);
	assign _3456_ = ~_1038_;
	assign _3457_ = (_4387_ ? _0403_ : _0903_);
	assign _3459_ = (_0127_ ? _3456_ : _3457_);
	assign _3460_ = (_0159_ ? _3455_ : _3459_);
	assign _3461_ = ~_1047_;
	assign _3462_ = ~_2484_;
	assign _3463_ = (_4423_ ? _0102_ : _3462_);
	assign _3464_ = (_0056_ ? _0140_ : _3463_);
	assign _3465_ = (_0146_ ? _3461_ : _3464_);
	assign _3466_ = (\mchip.pong.game.vga.pix_ind [0] ? _3465_ : _3460_);
	assign _3467_ = (_1103_ ? _3453_ : _3466_);
	assign _3468_ = ~_0309_;
	assign _3470_ = (_0127_ ? _0058_ : _1548_);
	assign _3471_ = (_0146_ ? _3468_ : _3470_);
	assign _3472_ = ~_0316_;
	assign _3473_ = (_0146_ ? _0047_ : _3472_);
	assign _3474_ = (\mchip.pong.game.vga.pix_ind [0] ? _3473_ : _3471_);
	assign _3475_ = ~_0319_;
	assign _3476_ = _0320_ | _0056_;
	assign _3477_ = (_0146_ ? _3476_ : _3475_);
	assign _3478_ = ~_0326_;
	assign _3479_ = _0323_ | _0056_;
	assign _3481_ = (_0146_ ? _3479_ : _3478_);
	assign _3482_ = (\mchip.pong.game.vga.pix_ind [0] ? _3481_ : _3477_);
	assign _3483_ = (_1103_ ? _3474_ : _3482_);
	assign _3484_ = (_0044_ ? _3467_ : _3483_);
	assign _3485_ = _0088_ & ~_3484_;
	assign _3486_ = _2976_ & ~_3485_;
	assign _3487_ = (_4368_ ? _3445_ : _3486_);
	assign _3488_ = (_4367_ ? _3343_ : _3487_);
	assign _3489_ = (_1058_ ? _3488_ : _2988_);
	assign _3490_ = (_0723_ ? _3250_ : _3489_);
	assign _3492_ = (_1061_ ? _2988_ : _3490_);
	assign \mchip.pong.VGA_R2  = _1264_ & ~_3492_;
	assign _3493_ = _1103_ & ~_1530_;
	assign _3494_ = _0063_ & ~_1539_;
	assign _3495_ = _3494_ | _3493_;
	assign _3496_ = _1551_ | _1546_;
	assign _3497_ = _4442_ & ~_1559_;
	assign _3498_ = \mchip.pong.game.vga.pix_ind [0] & ~_1564_;
	assign _3499_ = _3498_ | _3497_;
	assign _3500_ = (_1103_ ? _3496_ : _3499_);
	assign _3502_ = (_0044_ ? _3495_ : _3500_);
	assign _3503_ = ~(_1586_ & _0044_);
	assign _3504_ = _1595_ & ~_0044_;
	assign _3505_ = _3503_ & ~_3504_;
	assign _3506_ = (_0088_ ? _3502_ : _3505_);
	assign _3507_ = _0044_ & ~_1598_;
	assign _3508_ = (_1103_ ? _0218_ : _1604_);
	assign _3509_ = _3508_ & ~_0044_;
	assign _3510_ = _3509_ | _3507_;
	assign _3511_ = (_0044_ ? _1616_ : _1610_);
	assign _3513_ = (_0088_ ? _3510_ : _3511_);
	assign _3514_ = (_4368_ ? _3506_ : _3513_);
	assign _3515_ = _0088_ | ~_1673_;
	assign _3516_ = _1703_ & _0088_;
	assign _3517_ = _3515_ & ~_3516_;
	assign _3518_ = (_0044_ ? _1627_ : _1624_);
	assign _3519_ = _3518_ & ~_0152_;
	assign _3520_ = _0152_ & ~_1641_;
	assign _3521_ = _3520_ | _3519_;
	assign _3522_ = (_4368_ ? _3521_ : _3517_);
	assign _3524_ = (_4367_ ? _3514_ : _3522_);
	assign _3525_ = ~_1570_;
	assign _3526_ = _1571_ | _0127_;
	assign _3527_ = (_0146_ ? _3525_ : _3526_);
	assign _3528_ = ~_1575_;
	assign _3529_ = ~_1576_;
	assign _3530_ = (_0146_ ? _3528_ : _3529_);
	assign _3531_ = (\mchip.pong.game.vga.pix_ind [0] ? _3530_ : _3527_);
	assign _3532_ = ~_1580_;
	assign _3533_ = (_0146_ ? _3532_ : _2994_);
	assign _3535_ = ~_0096_;
	assign _3536_ = ~_1583_;
	assign _3537_ = (_0146_ ? _3536_ : _3535_);
	assign _3538_ = (\mchip.pong.game.vga.pix_ind [0] ? _3537_ : _3533_);
	assign _3539_ = (_1103_ ? _3531_ : _3538_);
	assign _3540_ = (_0056_ ? _0783_ : _0166_);
	assign _3541_ = (_4423_ ? _2053_ : _0114_);
	assign _3542_ = (_0127_ ? _2014_ : _3541_);
	assign _3543_ = (_0146_ ? _3540_ : _3542_);
	assign _3544_ = ~(_0451_ & _4423_);
	assign _3546_ = (_0127_ ? _0128_ : _3544_);
	assign _3547_ = _0403_ | _4437_;
	assign _3548_ = (_4423_ ? _0792_ : _3547_);
	assign _3549_ = (_0056_ ? _0117_ : _3548_);
	assign _3550_ = (_0146_ ? _3546_ : _3549_);
	assign _3551_ = (\mchip.pong.game.vga.pix_ind [0] ? _3550_ : _3543_);
	assign _3552_ = (_0056_ ? _1651_ : _0766_);
	assign _3553_ = ~_1723_;
	assign _3554_ = (_0127_ ? _3146_ : _3553_);
	assign _3555_ = (_0146_ ? _3552_ : _3554_);
	assign _3557_ = (_0056_ ? _1569_ : _1747_);
	assign _3558_ = (_0146_ ? _1726_ : _3557_);
	assign _3559_ = (\mchip.pong.game.vga.pix_ind [0] ? _3558_ : _3555_);
	assign _3560_ = (_1103_ ? _3551_ : _3559_);
	assign _3561_ = (_0044_ ? _3539_ : _3560_);
	assign _3562_ = (_0088_ ? _3502_ : _3561_);
	assign _3563_ = ~_1740_;
	assign _3564_ = (_4423_ ? _0153_ : _1870_);
	assign _3565_ = _0056_ & ~_3564_;
	assign _3566_ = (_0146_ ? _3563_ : _3565_);
	assign _3568_ = (_0056_ ? _0727_ : _1798_);
	assign _3569_ = _0098_ & ~_2356_;
	assign _3570_ = (_0127_ ? _1738_ : _3569_);
	assign _3571_ = (_0146_ ? _3568_ : _3570_);
	assign _3572_ = (\mchip.pong.game.vga.pix_ind [0] ? _3571_ : _3566_);
	assign _3573_ = (_0127_ ? _1560_ : _1756_);
	assign _3574_ = (_0146_ ? _3568_ : _3573_);
	assign _3575_ = (_4387_ ? _0119_ : _0474_);
	assign _3576_ = (_0127_ ? _0166_ : _3575_);
	assign _3577_ = ~(_1764_ | _0127_);
	assign _3579_ = _3300_ | _3577_;
	assign _3580_ = (_0146_ ? _3576_ : _3579_);
	assign _3581_ = (\mchip.pong.game.vga.pix_ind [0] ? _3580_ : _3574_);
	assign _3582_ = (_1103_ ? _3572_ : _3581_);
	assign _3583_ = _4409_ | _4387_;
	assign _3584_ = _0056_ & ~_3583_;
	assign _3585_ = (_0146_ ? _1770_ : _3584_);
	assign _3586_ = (_0146_ ? _1777_ : _3584_);
	assign _3587_ = (\mchip.pong.game.vga.pix_ind [0] ? _3586_ : _3585_);
	assign _3589_ = ~_1784_;
	assign _3590_ = (_0056_ ? _0500_ : _3589_);
	assign _3591_ = (_0146_ ? _3590_ : _3584_);
	assign _3592_ = (_4423_ ? _0153_ : _0639_);
	assign _3593_ = _0056_ & ~_3592_;
	assign _3594_ = (_0146_ ? _3033_ : _3593_);
	assign _3595_ = (\mchip.pong.game.vga.pix_ind [0] ? _3594_ : _3591_);
	assign _3596_ = (_1103_ ? _3587_ : _3595_);
	assign _3597_ = (_0044_ ? _3582_ : _3596_);
	assign _3598_ = (_0127_ ? _0154_ : _0452_);
	assign _3600_ = ~_0435_;
	assign _3601_ = (_4412_ ? _0665_ : _3600_);
	assign _3602_ = _3601_ & ~_0127_;
	assign _3603_ = (_0146_ ? _3598_ : _3602_);
	assign _3604_ = _1806_ & ~_0056_;
	assign _3605_ = _4443_ | _4387_;
	assign _3606_ = _0056_ & ~_3605_;
	assign _3607_ = (_0146_ ? _3604_ : _3606_);
	assign _3608_ = (\mchip.pong.game.vga.pix_ind [0] ? _3607_ : _3603_);
	assign _3609_ = _4434_ | _4387_;
	assign _3611_ = _0056_ & ~_3609_;
	assign _3612_ = (_0146_ ? _1823_ : _3611_);
	assign _3613_ = (_1103_ ? _3608_ : _3612_);
	assign _3614_ = (_0127_ ? _2189_ : _1833_);
	assign _3615_ = (_0146_ ? _0155_ : _3614_);
	assign _3616_ = _4387_ & ~_0207_;
	assign _3617_ = (_0127_ ? _0154_ : _3616_);
	assign _3618_ = (_0056_ ? _0429_ : _0519_);
	assign _3619_ = (_0146_ ? _3617_ : _3618_);
	assign _3620_ = (\mchip.pong.game.vga.pix_ind [0] ? _3619_ : _3615_);
	assign _3622_ = _0435_ | _4387_;
	assign _3623_ = _0056_ & ~_3622_;
	assign _3624_ = (_0146_ ? _0155_ : _3623_);
	assign _3625_ = (_0127_ ? _0591_ : _3601_);
	assign _3626_ = (_0146_ ? _3598_ : _3625_);
	assign _3627_ = (\mchip.pong.game.vga.pix_ind [0] ? _3626_ : _3624_);
	assign _3628_ = (_1103_ ? _3620_ : _3627_);
	assign _3629_ = (_0044_ ? _3613_ : _3628_);
	assign _3630_ = (_0088_ ? _3597_ : _3629_);
	assign _3631_ = (_4368_ ? _3562_ : _3630_);
	assign _3633_ = _1996_ & _0088_;
	assign _3634_ = _3515_ & ~_3633_;
	assign _3635_ = (_0127_ ? _1806_ : _3151_);
	assign _3636_ = _1853_ | _4387_;
	assign _3637_ = _0056_ & ~_3636_;
	assign _3638_ = (_0146_ ? _3635_ : _3637_);
	assign _3639_ = (_0146_ ? _0155_ : _3637_);
	assign _3640_ = (\mchip.pong.game.vga.pix_ind [0] ? _3639_ : _3638_);
	assign _3641_ = _1889_ | _4387_;
	assign _3642_ = _0056_ & ~_3641_;
	assign _3644_ = (_0146_ ? _0155_ : _3642_);
	assign _3645_ = _4387_ & ~_0475_;
	assign _3646_ = (_0127_ ? _0154_ : _3645_);
	assign _3647_ = _4387_ & ~_1853_;
	assign _3648_ = (_0056_ ? _0429_ : _3647_);
	assign _3649_ = (_0146_ ? _3646_ : _3648_);
	assign _3650_ = (\mchip.pong.game.vga.pix_ind [0] ? _3649_ : _3644_);
	assign _3651_ = (_1103_ ? _3640_ : _3650_);
	assign _3652_ = _0054_ | _4423_;
	assign _3653_ = _0127_ & ~_3652_;
	assign _3655_ = (_0146_ ? _3653_ : _2066_);
	assign _3656_ = _3138_ & ~_0056_;
	assign _3657_ = _0056_ & ~_1912_;
	assign _3658_ = (_0146_ ? _3656_ : _3657_);
	assign _3659_ = (\mchip.pong.game.vga.pix_ind [0] ? _3658_ : _3655_);
	assign _3660_ = (_0127_ ? _3138_ : _3344_);
	assign _3661_ = _0056_ & ~_1920_;
	assign _3662_ = (_0146_ ? _3660_ : _3661_);
	assign _3663_ = _1927_ | _4387_;
	assign _3664_ = _0056_ & ~_3663_;
	assign _3666_ = (_0146_ ? _3152_ : _3664_);
	assign _3667_ = (\mchip.pong.game.vga.pix_ind [0] ? _3666_ : _3662_);
	assign _3668_ = (_1103_ ? _3659_ : _3667_);
	assign _3669_ = (_0044_ ? _3651_ : _3668_);
	assign _3670_ = _4387_ & ~_0451_;
	assign _3671_ = (_0127_ ? _1934_ : _3670_);
	assign _3672_ = (_0159_ ? _1939_ : _3671_);
	assign _3673_ = ~_1946_;
	assign _3674_ = (_0056_ ? _3670_ : _3193_);
	assign _3675_ = (_0146_ ? _3674_ : _3673_);
	assign _3677_ = (\mchip.pong.game.vga.pix_ind [0] ? _3675_ : _3672_);
	assign _3678_ = ~_1953_;
	assign _3679_ = _3193_ & ~_0056_;
	assign _3680_ = (_0159_ ? _3678_ : _3679_);
	assign _3681_ = _0127_ & ~_0742_;
	assign _3682_ = (_0056_ ? _0872_ : _3616_);
	assign _3683_ = (_0146_ ? _3681_ : _3682_);
	assign _3684_ = (\mchip.pong.game.vga.pix_ind [0] ? _3683_ : _3680_);
	assign _3685_ = (_1103_ ? _3677_ : _3684_);
	assign _3686_ = ~(_1968_ & _4442_);
	assign _3688_ = (_4387_ ? _4380_ : _0792_);
	assign _3689_ = (_0056_ ? _1971_ : _3688_);
	assign _3690_ = (_0146_ ? _3689_ : _0287_);
	assign _3691_ = \mchip.pong.game.vga.pix_ind [0] & ~_3690_;
	assign _3692_ = _3686_ & ~_3691_;
	assign _3693_ = (_0146_ ? _2006_ : _0287_);
	assign _3694_ = (_0159_ ? _1983_ : _2042_);
	assign _3695_ = (\mchip.pong.game.vga.pix_ind [0] ? _3694_ : _3693_);
	assign _3696_ = (_1103_ ? _3692_ : _3695_);
	assign _3697_ = (_0044_ ? _3685_ : _3696_);
	assign _3699_ = (_0088_ ? _3669_ : _3697_);
	assign _3700_ = (_4368_ ? _3699_ : _3634_);
	assign _3701_ = (_4367_ ? _3631_ : _3700_);
	assign _3702_ = (\mchip.pong.game.vga.pix_ind [0] ? _2004_ : _2009_);
	assign _3703_ = ~_2020_;
	assign _3704_ = (_0146_ ? _3451_ : _3703_);
	assign _3705_ = (\mchip.pong.game.vga.pix_ind [0] ? _3704_ : _2017_);
	assign _3706_ = (_1103_ ? _3702_ : _3705_);
	assign _3707_ = (_0044_ ? _3539_ : _3706_);
	assign _3708_ = (_0088_ ? _3502_ : _3707_);
	assign _3710_ = _2063_ & ~_2074_;
	assign _3711_ = (_4423_ ? _0425_ : _0391_);
	assign _3712_ = (_0056_ ? _0500_ : _3711_);
	assign _3713_ = (_0146_ ? _3712_ : _2071_);
	assign _3714_ = _0761_ & ~_0127_;
	assign _3715_ = (_0146_ ? _2037_ : _3714_);
	assign _3716_ = (\mchip.pong.game.vga.pix_ind [0] ? _3715_ : _3713_);
	assign _3717_ = ~(_0972_ | _0127_);
	assign _3718_ = (_0146_ ? _2042_ : _3717_);
	assign _3719_ = (_0146_ ? _2006_ : _3577_);
	assign _3721_ = (\mchip.pong.game.vga.pix_ind [0] ? _3719_ : _3718_);
	assign _3722_ = (_1103_ ? _3716_ : _3721_);
	assign _3723_ = (_0044_ ? _3722_ : _3710_);
	assign _3724_ = ~(_2090_ & \mchip.pong.game.vga.pix_ind [0]);
	assign _3725_ = (_4423_ ? _4389_ : _0292_);
	assign _3726_ = (_0127_ ? _0199_ : _3725_);
	assign _3727_ = (_0146_ ? _3726_ : _2081_);
	assign _3728_ = _4442_ & ~_3727_;
	assign _3729_ = _3724_ & ~_3728_;
	assign _3730_ = ~_2092_;
	assign _3732_ = (_0056_ ? _0500_ : _3730_);
	assign _3733_ = ~_2094_;
	assign _3734_ = (_0127_ ? _1850_ : _3733_);
	assign _3735_ = (_0146_ ? _3732_ : _3734_);
	assign _3736_ = ~_2098_;
	assign _3737_ = (_0056_ ? _1817_ : _3736_);
	assign _3738_ = _4420_ & ~_4423_;
	assign _3739_ = (_0056_ ? _3733_ : _3738_);
	assign _3740_ = (_0146_ ? _3737_ : _3739_);
	assign _3741_ = (\mchip.pong.game.vga.pix_ind [0] ? _3740_ : _3735_);
	assign _3743_ = (_1103_ ? _3729_ : _3741_);
	assign _3744_ = ~_2105_;
	assign _3745_ = (_0056_ ? _1532_ : _3744_);
	assign _3746_ = (_0146_ ? _3745_ : _2112_);
	assign _3747_ = ~_2108_;
	assign _3748_ = (_4387_ ? _0292_ : _0403_);
	assign _3749_ = (_0127_ ? _3747_ : _3748_);
	assign _3750_ = (_0146_ ? _3749_ : _2112_);
	assign _3751_ = (\mchip.pong.game.vga.pix_ind [0] ? _3750_ : _3746_);
	assign _3752_ = (_0159_ ? _2112_ : _3726_);
	assign _3754_ = (_4387_ ? _0292_ : _0114_);
	assign _3755_ = (_0127_ ? _0199_ : _3754_);
	assign _3756_ = (_0146_ ? _3755_ : _2112_);
	assign _3757_ = (\mchip.pong.game.vga.pix_ind [0] ? _3756_ : _3752_);
	assign _3758_ = (_1103_ ? _3751_ : _3757_);
	assign _3759_ = (_0044_ ? _3743_ : _3758_);
	assign _3760_ = (_0088_ ? _3723_ : _3759_);
	assign _3761_ = (_4368_ ? _3708_ : _3760_);
	assign _3762_ = _0127_ & ~_2123_;
	assign _3763_ = (_0159_ ? _2125_ : _3762_);
	assign _3765_ = (_0159_ ? _2125_ : _2132_);
	assign _3766_ = (\mchip.pong.game.vga.pix_ind [0] ? _3765_ : _3763_);
	assign _3767_ = (_0127_ ? _3355_ : _2080_);
	assign _3768_ = (_0146_ ? _2132_ : _3767_);
	assign _3769_ = (_0146_ ? _2132_ : _2138_);
	assign _3770_ = (\mchip.pong.game.vga.pix_ind [0] ? _3769_ : _3768_);
	assign _3771_ = (_1103_ ? _3766_ : _3770_);
	assign _3772_ = (_4387_ ? _2053_ : _0254_);
	assign _3773_ = (_0056_ ? _0875_ : _3772_);
	assign _3774_ = (_0056_ ? _3295_ : _1971_);
	assign _3776_ = (_0146_ ? _3773_ : _3774_);
	assign _3777_ = ~_2057_;
	assign _3778_ = ~_2149_;
	assign _3779_ = (_0056_ ? _0875_ : _3778_);
	assign _3780_ = (_0146_ ? _3779_ : _3777_);
	assign _3781_ = (\mchip.pong.game.vga.pix_ind [0] ? _3780_ : _3776_);
	assign _3782_ = ~_2153_;
	assign _3783_ = (_0056_ ? _0875_ : _3782_);
	assign _3784_ = (_0146_ ? _3783_ : _2066_);
	assign _3785_ = (_4387_ ? _2053_ : _0094_);
	assign _3787_ = (_0056_ ? _0875_ : _3785_);
	assign _3788_ = (_0146_ ? _3787_ : _2159_);
	assign _3789_ = (\mchip.pong.game.vga.pix_ind [0] ? _3788_ : _3784_);
	assign _3790_ = (_1103_ ? _3781_ : _3789_);
	assign _3791_ = (_0044_ ? _3771_ : _3790_);
	assign _3792_ = (_4387_ ? _0292_ : _0118_);
	assign _3793_ = (_0127_ ? _1798_ : _3792_);
	assign _3794_ = (_0127_ ? _1555_ : _3395_);
	assign _3795_ = (_0146_ ? _3793_ : _3794_);
	assign _3796_ = _0146_ | ~_2174_;
	assign _3798_ = _0146_ & ~_2070_;
	assign _3799_ = _3796_ & ~_3798_;
	assign _3800_ = (\mchip.pong.game.vga.pix_ind [0] ? _3799_ : _3795_);
	assign _3801_ = (_0056_ ? _0500_ : _0162_);
	assign _3802_ = _4423_ | ~_0093_;
	assign _3803_ = _3802_ & ~_3171_;
	assign _3804_ = (_0056_ ? _3782_ : _3803_);
	assign _3805_ = (_0146_ ? _3801_ : _3804_);
	assign _3806_ = ~_2184_;
	assign _3807_ = (_0127_ ? _0162_ : _0875_);
	assign _3809_ = (_0159_ ? _3806_ : _3807_);
	assign _3810_ = (\mchip.pong.game.vga.pix_ind [0] ? _3809_ : _3805_);
	assign _3811_ = (_1103_ ? _3800_ : _3810_);
	assign _3812_ = _0146_ | ~_2195_;
	assign _3813_ = _0127_ & ~_2191_;
	assign _3814_ = _0146_ & ~_3813_;
	assign _3815_ = _3812_ & ~_3814_;
	assign _3816_ = ~_2197_;
	assign _3817_ = (_0127_ ? _3816_ : _3792_);
	assign _3818_ = (_4387_ ? _0404_ : _2202_);
	assign _3820_ = (_4423_ ? _2053_ : _0089_);
	assign _3821_ = (_0127_ ? _3818_ : _3820_);
	assign _3822_ = (_0146_ ? _3817_ : _3821_);
	assign _3823_ = (\mchip.pong.game.vga.pix_ind [0] ? _3822_ : _3815_);
	assign _3824_ = _0146_ | ~_2211_;
	assign _3825_ = (_0056_ ? _0068_ : _1976_);
	assign _3826_ = _3825_ & ~_0159_;
	assign _3827_ = _3824_ & ~_3826_;
	assign _3828_ = ~_2213_;
	assign _3829_ = (_0056_ ? _1557_ : _3828_);
	assign _3831_ = (_4387_ ? _0035_ : _0206_);
	assign _3832_ = (_0056_ ? _1756_ : _3831_);
	assign _3833_ = (_0146_ ? _3829_ : _3832_);
	assign _3834_ = (\mchip.pong.game.vga.pix_ind [0] ? _3833_ : _3827_);
	assign _3835_ = (_1103_ ? _3823_ : _3834_);
	assign _3836_ = (_0044_ ? _3811_ : _3835_);
	assign _3837_ = (_0088_ ? _3791_ : _3836_);
	assign _3838_ = _0128_ | _0127_;
	assign _3839_ = (_0146_ ? _3479_ : _3838_);
	assign _3840_ = (_0146_ ? _3446_ : _3526_);
	assign _3842_ = (\mchip.pong.game.vga.pix_ind [0] ? _3840_ : _3839_);
	assign _3843_ = _0127_ & ~_2225_;
	assign _3844_ = (_0159_ ? _2228_ : _3843_);
	assign _3845_ = (_4423_ ? _0131_ : _2200_);
	assign _3846_ = (_0056_ ? _0330_ : _3845_);
	assign _3847_ = (_0146_ ? _2233_ : _3846_);
	assign _3848_ = (\mchip.pong.game.vga.pix_ind [0] ? _3847_ : _3844_);
	assign _3849_ = (_1103_ ? _3842_ : _3848_);
	assign _3850_ = (_0056_ ? _0052_ : _0197_);
	assign _3851_ = _0193_ | _0127_;
	assign _3853_ = (_0146_ ? _3850_ : _3851_);
	assign _3854_ = _1679_ | _0127_;
	assign _3855_ = (_0146_ ? _1541_ : _3854_);
	assign _3856_ = (\mchip.pong.game.vga.pix_ind [0] ? _3855_ : _3853_);
	assign _3857_ = _1683_ | _0056_;
	assign _3858_ = _0402_ | _0127_;
	assign _3859_ = (_0146_ ? _3857_ : _3858_);
	assign _3860_ = _0288_ | _0127_;
	assign _3861_ = (_0146_ ? _3476_ : _3860_);
	assign _3862_ = (\mchip.pong.game.vga.pix_ind [0] ? _3861_ : _3859_);
	assign _3864_ = (_1103_ ? _3856_ : _3862_);
	assign _3865_ = (_0044_ ? _3849_ : _3864_);
	assign _3866_ = _0088_ & ~_3865_;
	assign _3867_ = _3515_ & ~_3866_;
	assign _3868_ = (_4368_ ? _3837_ : _3867_);
	assign _3869_ = (_4367_ ? _3761_ : _3868_);
	assign _3870_ = (_1058_ ? _3869_ : _3524_);
	assign _3871_ = (_0723_ ? _3701_ : _3870_);
	assign _3872_ = (_1061_ ? _3524_ : _3871_);
	assign \mchip.pong.VGA_R3  = _1264_ & ~_3872_;
	assign \mchip.pong.game.right_paddle.next_coord [1] = _0927_ ^ \mchip.pong.game.right_paddle.coord [0];
	assign \mchip.pong.game.left_paddle.next_coord [1] = _0677_ ^ \mchip.pong.game.left_paddle.coord [0];
	assign _3874_ = ~(\mchip.pong.game.ball.cpath.state [3] | \mchip.pong.game.ball.cpath.state [5]);
	assign _3875_ = _3874_ ^ \mchip.pong.game.ball.dpath.ballX [2];
	assign \mchip.pong.game.ball.dpath.nextX [2] = _3875_ ^ \mchip.pong.game.ball.dpath.ballX [1];
	assign _3876_ = ~(_3874_ & \mchip.pong.game.ball.dpath.ballX [2]);
	assign _3877_ = ~(_3875_ & \mchip.pong.game.ball.dpath.ballX [1]);
	assign _3878_ = ~(_3877_ & _3876_);
	assign _3879_ = _3874_ ^ \mchip.pong.game.ball.dpath.ballX [3];
	assign \mchip.pong.game.ball.dpath.nextX [3] = _3879_ ^ _3878_;
	assign _3881_ = _3874_ & \mchip.pong.game.ball.dpath.ballX [3];
	assign _3882_ = _3879_ & _3878_;
	assign _3883_ = _3882_ | _3881_;
	assign _3884_ = _3874_ ^ \mchip.pong.game.ball.dpath.ballX [4];
	assign \mchip.pong.game.ball.dpath.nextX [4] = _3884_ ^ _3883_;
	assign _3885_ = ~(_3874_ & \mchip.pong.game.ball.dpath.ballX [4]);
	assign _3886_ = ~(_3884_ & _3881_);
	assign _3887_ = ~(_3886_ & _3885_);
	assign _3888_ = ~(_3884_ & _3879_);
	assign _3889_ = _3878_ & ~_3888_;
	assign _3891_ = _3889_ | _3887_;
	assign _3892_ = _3874_ ^ \mchip.pong.game.ball.dpath.ballX [5];
	assign \mchip.pong.game.ball.dpath.nextX [5] = _3892_ ^ _3891_;
	assign _3893_ = _3874_ & \mchip.pong.game.ball.dpath.ballX [5];
	assign _3894_ = _3892_ & _3891_;
	assign _3895_ = _3894_ | _3893_;
	assign _3896_ = _3874_ ^ \mchip.pong.game.ball.dpath.ballX [6];
	assign \mchip.pong.game.ball.dpath.nextX [6] = _3896_ ^ _3895_;
	assign _3897_ = _3874_ & ~_1085_;
	assign _3898_ = _3896_ & _3893_;
	assign _3900_ = _3898_ | _3897_;
	assign _3901_ = ~(_3896_ & _3892_);
	assign _3902_ = _3891_ & ~_3901_;
	assign _3903_ = _3902_ | _3900_;
	assign _3904_ = _3874_ ^ \mchip.pong.game.ball.dpath.ballX [7];
	assign \mchip.pong.game.ball.dpath.nextX [7] = _3904_ ^ _3903_;
	assign _3905_ = _3874_ & ~_3271_;
	assign _3906_ = _3904_ & _3903_;
	assign _3907_ = _3906_ | _3905_;
	assign _3908_ = _3874_ ^ \mchip.pong.game.ball.dpath.ballX [8];
	assign \mchip.pong.game.ball.dpath.nextX [8] = _3908_ ^ _3907_;
	assign _3910_ = _3874_ & ~_1074_;
	assign _3911_ = _3908_ & _3905_;
	assign _3912_ = _3911_ | _3910_;
	assign _3913_ = ~(_3908_ & _3904_);
	assign _3914_ = _3900_ & ~_3913_;
	assign _3915_ = _3914_ | _3912_;
	assign _3916_ = _3913_ | _3901_;
	assign _3917_ = _3891_ & ~_3916_;
	assign _3918_ = _3917_ | _3915_;
	assign _3920_ = _3874_ ^ \mchip.pong.game.ball.dpath.ballX [9];
	assign \mchip.pong.game.ball.dpath.nextX [9] = _3920_ ^ _3918_;
	assign _3921_ = _4165_ ^ \mchip.pong.game.ball.dpath.ballY [1];
	assign \mchip.pong.game.ball.dpath.nextY [1] = _3921_ ^ \mchip.pong.game.ball.dpath.ballY [0];
	assign _3922_ = _4165_ & ~_3073_;
	assign _3923_ = _3921_ & ~\mchip.pong.game.ball.dpath.nextY [0];
	assign _3924_ = _3923_ | _3922_;
	assign _3925_ = _4165_ ^ \mchip.pong.game.ball.dpath.ballY [2];
	assign \mchip.pong.game.ball.dpath.nextY [2] = _3925_ ^ _3924_;
	assign _3926_ = _4165_ & ~_3029_;
	assign _3927_ = _3925_ & _3924_;
	assign _3928_ = _3927_ | _3926_;
	assign _3929_ = _4165_ ^ \mchip.pong.game.ball.dpath.ballY [3];
	assign \mchip.pong.game.ball.dpath.nextY [3] = _3929_ ^ _3928_;
	assign _3930_ = _4165_ & ~_4393_;
	assign _3931_ = _3929_ & _3926_;
	assign _3932_ = _3931_ | _3930_;
	assign _3933_ = ~(_3929_ & _3925_);
	assign _3934_ = _3924_ & ~_3933_;
	assign _3935_ = _3934_ | _3932_;
	assign _3937_ = _4165_ ^ \mchip.pong.game.ball.dpath.ballY [4];
	assign \mchip.pong.game.ball.dpath.nextY [4] = _3937_ ^ _3935_;
	assign _3938_ = _4165_ & ~_2625_;
	assign _3939_ = _3937_ & _3935_;
	assign _3940_ = _3939_ | _3938_;
	assign _3941_ = _4165_ ^ \mchip.pong.game.ball.dpath.ballY [5];
	assign \mchip.pong.game.ball.dpath.nextY [5] = _3941_ ^ _3940_;
	assign _3942_ = _4165_ & ~_2658_;
	assign _3943_ = _3941_ & _3938_;
	assign _3944_ = _3943_ | _3942_;
	assign _3946_ = ~(_3941_ & _3937_);
	assign _3947_ = _3935_ & ~_3946_;
	assign _3948_ = _3947_ | _3944_;
	assign _3949_ = _4165_ ^ \mchip.pong.game.ball.dpath.ballY [6];
	assign \mchip.pong.game.ball.dpath.nextY [6] = _3949_ ^ _3948_;
	assign _3950_ = _4165_ & ~_1739_;
	assign _3951_ = _3949_ & _3948_;
	assign _3952_ = _3951_ | _3950_;
	assign _3953_ = _4165_ ^ \mchip.pong.game.ball.dpath.ballY [7];
	assign \mchip.pong.game.ball.dpath.nextY [7] = _3953_ ^ _3952_;
	assign _3955_ = _4165_ & ~_2877_;
	assign _3956_ = _3953_ & _3950_;
	assign _3957_ = _3956_ | _3955_;
	assign _3958_ = ~(_3953_ & _3949_);
	assign _3959_ = _3944_ & ~_3958_;
	assign _3960_ = _3959_ | _3957_;
	assign _3961_ = _3958_ | _3946_;
	assign _3962_ = _3935_ & ~_3961_;
	assign _3963_ = _3962_ | _3960_;
	assign _3964_ = _4165_ ^ \mchip.pong.game.ball.dpath.ballY [8];
	assign \mchip.pong.game.ball.dpath.nextY [8] = _3964_ ^ _3963_;
	always @(posedge io_in[12])
		if (_0010_)
			\mchip.pong.game.vga.pclk_ctr  <= 1'h0;
		else
			\mchip.pong.game.vga.pclk_ctr  <= _4446_;
	always @(posedge io_in[12]) \mchip.pong.game.ball.cpath.state [0] <= _0000_;
	always @(posedge io_in[12]) \mchip.pong.game.ball.cpath.state [1] <= _0001_;
	always @(posedge io_in[12]) \mchip.pong.game.ball.cpath.state [2] <= _0002_;
	always @(posedge io_in[12]) \mchip.pong.game.ball.cpath.state [3] <= _0003_;
	always @(posedge io_in[12]) \mchip.pong.game.ball.cpath.state [4] <= _0004_;
	always @(posedge io_in[12]) \mchip.pong.game.ball.cpath.state [5] <= _0005_;
	always @(posedge io_in[12]) \mchip.pong.game.ball.cpath.state [6] <= _0006_;
	always @(posedge io_in[12]) \mchip.pong.game.ball.cpath.state [7] <= _0007_;
	always @(posedge io_in[12]) \mchip.pong.game.ball.cpath.state [8] <= _0008_;
	always @(posedge io_in[12]) \mchip.pong.sync.o_out [0] <= \mchip.pong.sync.sync [0];
	always @(posedge io_in[12]) \mchip.pong.sync.o_out [1] <= \mchip.pong.sync.sync [1];
	always @(posedge io_in[12]) \mchip.pong.sync.o_out [2] <= \mchip.pong.sync.sync [2];
	always @(posedge io_in[12]) \mchip.pong.sync.o_out [3] <= \mchip.pong.sync.sync [3];
	always @(posedge io_in[12]) \mchip.pong.sync.o_out [4] <= \mchip.pong.sync.sync [4];
	always @(posedge io_in[12]) \mchip.pong.sync.o_out [5] <= \mchip.pong.sync.sync [5];
	always @(posedge io_in[12]) \mchip.pong.sync.o_out [6] <= \mchip.pong.sync.sync [6];
	always @(posedge io_in[12]) \mchip.pong.sync.o_out [7] <= \mchip.pong.sync.sync [7];
	always @(posedge io_in[12]) \mchip.pong.sync.sync [0] <= io_in[6];
	always @(posedge io_in[12]) \mchip.pong.sync.sync [1] <= io_in[7];
	always @(posedge io_in[12]) \mchip.pong.sync.sync [2] <= io_in[4];
	always @(posedge io_in[12]) \mchip.pong.sync.sync [3] <= io_in[5];
	always @(posedge io_in[12]) \mchip.pong.sync.sync [4] <= io_in[0];
	always @(posedge io_in[12]) \mchip.pong.sync.sync [5] <= io_in[1];
	always @(posedge io_in[12]) \mchip.pong.sync.sync [6] <= io_in[2];
	always @(posedge io_in[12]) \mchip.pong.sync.sync [7] <= io_in[3];
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [0] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [0] <= _0023_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [1] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [1] <= _0024_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [2] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [2] <= _0025_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [3] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [3] <= _0026_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [4] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [4] <= _0027_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [5] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [5] <= _0028_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [6] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [6] <= _0029_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [7] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [7] <= _0030_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [8] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [8] <= _0031_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.pix_ind [9] <= 1'h0;
		else if (!\mchip.pong.game.vga.pclk_ctr )
			\mchip.pong.game.vga.pix_ind [9] <= _0032_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [0] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [0] <= _0013_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [1] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [1] <= _0014_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [2] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [2] <= _0015_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [3] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [3] <= _0016_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [4] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [4] <= _0017_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [5] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [5] <= _0018_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [6] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [6] <= _0019_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [7] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [7] <= _0020_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [8] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [8] <= _0021_;
	always @(posedge io_in[12])
		if (\mchip.pong.sync.o_out [2])
			\mchip.pong.game.vga.line_ind [9] <= 1'h0;
		else if (_0009_)
			\mchip.pong.game.vga.line_ind [9] <= _0022_;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.right_paddle.coord [0] <= 1'h0;
		else if (_0012_)
			\mchip.pong.game.right_paddle.coord [0] <= \mchip.pong.game.right_paddle.next_coord [0];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.right_paddle.coord [1] <= 1'h0;
		else if (_0012_)
			\mchip.pong.game.right_paddle.coord [1] <= \mchip.pong.game.right_paddle.next_coord [1];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.right_paddle.coord [2] <= 1'h0;
		else if (_0012_)
			\mchip.pong.game.right_paddle.coord [2] <= \mchip.pong.game.right_paddle.next_coord [2];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.right_paddle.coord [3] <= 1'h0;
		else if (_0012_)
			\mchip.pong.game.right_paddle.coord [3] <= \mchip.pong.game.right_paddle.next_coord [3];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.right_paddle.coord [4] <= 1'h0;
		else if (_0012_)
			\mchip.pong.game.right_paddle.coord [4] <= \mchip.pong.game.right_paddle.next_coord [4];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.right_paddle.coord [5] <= 1'h0;
		else if (_0012_)
			\mchip.pong.game.right_paddle.coord [5] <= \mchip.pong.game.right_paddle.next_coord [5];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.right_paddle.coord [6] <= 1'h0;
		else if (_0012_)
			\mchip.pong.game.right_paddle.coord [6] <= \mchip.pong.game.right_paddle.next_coord [6];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.right_paddle.coord [7] <= 1'h0;
		else if (_0012_)
			\mchip.pong.game.right_paddle.coord [7] <= \mchip.pong.game.right_paddle.next_coord [7];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.right_paddle.coord [8] <= 1'h0;
		else if (_0012_)
			\mchip.pong.game.right_paddle.coord [8] <= \mchip.pong.game.right_paddle.next_coord [8];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.left_paddle.coord [0] <= 1'h0;
		else if (_0011_)
			\mchip.pong.game.left_paddle.coord [0] <= \mchip.pong.game.left_paddle.next_coord [0];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.left_paddle.coord [1] <= 1'h0;
		else if (_0011_)
			\mchip.pong.game.left_paddle.coord [1] <= \mchip.pong.game.left_paddle.next_coord [1];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.left_paddle.coord [2] <= 1'h0;
		else if (_0011_)
			\mchip.pong.game.left_paddle.coord [2] <= \mchip.pong.game.left_paddle.next_coord [2];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.left_paddle.coord [3] <= 1'h0;
		else if (_0011_)
			\mchip.pong.game.left_paddle.coord [3] <= \mchip.pong.game.left_paddle.next_coord [3];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.left_paddle.coord [4] <= 1'h0;
		else if (_0011_)
			\mchip.pong.game.left_paddle.coord [4] <= \mchip.pong.game.left_paddle.next_coord [4];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.left_paddle.coord [5] <= 1'h0;
		else if (_0011_)
			\mchip.pong.game.left_paddle.coord [5] <= \mchip.pong.game.left_paddle.next_coord [5];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.left_paddle.coord [6] <= 1'h0;
		else if (_0011_)
			\mchip.pong.game.left_paddle.coord [6] <= \mchip.pong.game.left_paddle.next_coord [6];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.left_paddle.coord [7] <= 1'h0;
		else if (_0011_)
			\mchip.pong.game.left_paddle.coord [7] <= \mchip.pong.game.left_paddle.next_coord [7];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.cpath.state [0])
			\mchip.pong.game.left_paddle.coord [8] <= 1'h0;
		else if (_0011_)
			\mchip.pong.game.left_paddle.coord [8] <= \mchip.pong.game.left_paddle.next_coord [8];
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballY [0] <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballY [0] <= \mchip.pong.game.ball.dpath.nextY [0];
		end
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballY [1] <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballY [1] <= \mchip.pong.game.ball.dpath.nextY [1];
		end
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballY [2] <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballY [2] <= \mchip.pong.game.ball.dpath.nextY [2];
		end
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballY [3] <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballY [3] <= \mchip.pong.game.ball.dpath.nextY [3];
		end
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballY [4] <= 1'h1;
			else
				\mchip.pong.game.ball.dpath.ballY [4] <= \mchip.pong.game.ball.dpath.nextY [4];
		end
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballY [5] <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballY [5] <= \mchip.pong.game.ball.dpath.nextY [5];
		end
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballY [6] <= 1'h1;
			else
				\mchip.pong.game.ball.dpath.ballY [6] <= \mchip.pong.game.ball.dpath.nextY [6];
		end
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballY [7] <= 1'h1;
			else
				\mchip.pong.game.ball.dpath.ballY [7] <= \mchip.pong.game.ball.dpath.nextY [7];
		end
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballY [8] <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballY [8] <= \mchip.pong.game.ball.dpath.nextY [8];
		end
	reg \mchip.pong.game.ball.dpath.ballX_reg[1] ;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballX_reg[1]  <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballX_reg[1]  <= \mchip.pong.game.ball.dpath.nextX [1];
		end
	assign \mchip.pong.game.ball.dpath.ballX [1] = \mchip.pong.game.ball.dpath.ballX_reg[1] ;
	reg \mchip.pong.game.ball.dpath.ballX_reg[2] ;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballX_reg[2]  <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballX_reg[2]  <= \mchip.pong.game.ball.dpath.nextX [2];
		end
	assign \mchip.pong.game.ball.dpath.ballX [2] = \mchip.pong.game.ball.dpath.ballX_reg[2] ;
	reg \mchip.pong.game.ball.dpath.ballX_reg[3] ;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballX_reg[3]  <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballX_reg[3]  <= \mchip.pong.game.ball.dpath.nextX [3];
		end
	assign \mchip.pong.game.ball.dpath.ballX [3] = \mchip.pong.game.ball.dpath.ballX_reg[3] ;
	reg \mchip.pong.game.ball.dpath.ballX_reg[4] ;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballX_reg[4]  <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballX_reg[4]  <= \mchip.pong.game.ball.dpath.nextX [4];
		end
	assign \mchip.pong.game.ball.dpath.ballX [4] = \mchip.pong.game.ball.dpath.ballX_reg[4] ;
	reg \mchip.pong.game.ball.dpath.ballX_reg[5] ;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballX_reg[5]  <= 1'h1;
			else
				\mchip.pong.game.ball.dpath.ballX_reg[5]  <= \mchip.pong.game.ball.dpath.nextX [5];
		end
	assign \mchip.pong.game.ball.dpath.ballX [5] = \mchip.pong.game.ball.dpath.ballX_reg[5] ;
	reg \mchip.pong.game.ball.dpath.ballX_reg[6] ;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballX_reg[6]  <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballX_reg[6]  <= \mchip.pong.game.ball.dpath.nextX [6];
		end
	assign \mchip.pong.game.ball.dpath.ballX [6] = \mchip.pong.game.ball.dpath.ballX_reg[6] ;
	reg \mchip.pong.game.ball.dpath.ballX_reg[7] ;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballX_reg[7]  <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballX_reg[7]  <= \mchip.pong.game.ball.dpath.nextX [7];
		end
	assign \mchip.pong.game.ball.dpath.ballX [7] = \mchip.pong.game.ball.dpath.ballX_reg[7] ;
	reg \mchip.pong.game.ball.dpath.ballX_reg[8] ;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballX_reg[8]  <= 1'h1;
			else
				\mchip.pong.game.ball.dpath.ballX_reg[8]  <= \mchip.pong.game.ball.dpath.nextX [8];
		end
	assign \mchip.pong.game.ball.dpath.ballX [8] = \mchip.pong.game.ball.dpath.ballX_reg[8] ;
	reg \mchip.pong.game.ball.dpath.ballX_reg[9] ;
	always @(posedge io_in[12])
		if (\mchip.pong.game.ball.dpath.en_pos_reg ) begin
			if (_0033_)
				\mchip.pong.game.ball.dpath.ballX_reg[9]  <= 1'h0;
			else
				\mchip.pong.game.ball.dpath.ballX_reg[9]  <= \mchip.pong.game.ball.dpath.nextX [9];
		end
	assign \mchip.pong.game.ball.dpath.ballX [9] = \mchip.pong.game.ball.dpath.ballX_reg[9] ;
	assign io_out = {6'h00, \mchip.pong.VGA_R3 , \mchip.pong.VGA_R2 , \mchip.pong.VGA_G3 , \mchip.pong.VGA_G2 , \mchip.pong.VGA_B3 , \mchip.pong.VGA_B2 , \mchip.pong.VGA_VS , \mchip.pong.VGA_HS };
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {4'h0, \mchip.pong.VGA_R3 , \mchip.pong.VGA_R2 , \mchip.pong.VGA_G3 , \mchip.pong.VGA_G2 , \mchip.pong.VGA_B3 , \mchip.pong.VGA_B2 , \mchip.pong.VGA_VS , \mchip.pong.VGA_HS };
	assign \mchip.pong.VGA_B  = {\mchip.pong.VGA_B3 , \mchip.pong.VGA_B2 , 6'h00};
	assign \mchip.pong.VGA_B0  = 1'h0;
	assign \mchip.pong.VGA_B1  = 1'h0;
	assign \mchip.pong.VGA_G  = {\mchip.pong.VGA_G3 , \mchip.pong.VGA_G2 , 6'h00};
	assign \mchip.pong.VGA_G0  = 1'h0;
	assign \mchip.pong.VGA_G1  = 1'h0;
	assign \mchip.pong.VGA_R  = {\mchip.pong.VGA_R3 , \mchip.pong.VGA_R2 , 6'h00};
	assign \mchip.pong.VGA_R0  = 1'h0;
	assign \mchip.pong.VGA_R1  = 1'h0;
	assign \mchip.pong.btn_rst  = io_in[4];
	assign \mchip.pong.btn_serve  = io_in[5];
	assign \mchip.pong.cfg1  = io_in[7];
	assign \mchip.pong.cfg1_o  = \mchip.pong.sync.o_out [1];
	assign \mchip.pong.cfg2  = io_in[6];
	assign \mchip.pong.cfg2_o  = \mchip.pong.sync.o_out [0];
	assign \mchip.pong.clk_25mhz  = io_in[12];
	assign \mchip.pong.game.Cnewgame  = \mchip.pong.game.ball.cpath.state [0];
	assign \mchip.pong.game.VGA_B  = {\mchip.pong.VGA_B3 , \mchip.pong.VGA_B2 , 6'h00};
	assign \mchip.pong.game.VGA_G  = {\mchip.pong.VGA_G3 , \mchip.pong.VGA_G2 , 6'h00};
	assign \mchip.pong.game.VGA_HS  = \mchip.pong.VGA_HS ;
	assign \mchip.pong.game.VGA_R  = {\mchip.pong.VGA_R3 , \mchip.pong.VGA_R2 , 6'h00};
	assign \mchip.pong.game.VGA_VS  = \mchip.pong.VGA_VS ;
	assign \mchip.pong.game.ball.Cnewgame  = \mchip.pong.game.ball.cpath.state [0];
	assign \mchip.pong.game.ball.ballX  = {\mchip.pong.game.ball.dpath.ballX [9:1], 1'h0};
	assign \mchip.pong.game.ball.ballY  = \mchip.pong.game.ball.dpath.ballY ;
	assign \mchip.pong.game.ball.clock  = io_in[12];
	assign \mchip.pong.game.ball.cpath.Cnewgame  = \mchip.pong.game.ball.cpath.state [0];
	assign \mchip.pong.game.ball.cpath.clock  = io_in[12];
	assign \mchip.pong.game.ball.cpath.reset  = \mchip.pong.sync.o_out [2];
	assign \mchip.pong.game.ball.cpath.serve_input  = \mchip.pong.sync.o_out [3];
	assign \mchip.pong.game.ball.dpath.Cnewgame  = \mchip.pong.game.ball.cpath.state [0];
	assign \mchip.pong.game.ball.dpath.ballX [0] = 1'h0;
	assign \mchip.pong.game.ball.dpath.clock  = io_in[12];
	assign \mchip.pong.game.ball.dpath.nextX [0] = 1'h0;
	assign \mchip.pong.game.ball.dpath.paddleLY  = \mchip.pong.game.left_paddle.coord ;
	assign \mchip.pong.game.ball.dpath.paddleRY  = \mchip.pong.game.right_paddle.coord ;
	assign \mchip.pong.game.ball.paddleLY  = \mchip.pong.game.left_paddle.coord ;
	assign \mchip.pong.game.ball.paddleRY  = \mchip.pong.game.right_paddle.coord ;
	assign \mchip.pong.game.ball.reset  = \mchip.pong.sync.o_out [2];
	assign \mchip.pong.game.ball.serve_input  = \mchip.pong.sync.o_out [3];
	assign \mchip.pong.game.ballX  = {\mchip.pong.game.ball.dpath.ballX [9:1], 1'h0};
	assign \mchip.pong.game.ballY  = \mchip.pong.game.ball.dpath.ballY ;
	assign \mchip.pong.game.cfg1  = \mchip.pong.sync.o_out [1];
	assign \mchip.pong.game.cfg2  = \mchip.pong.sync.o_out [0];
	assign \mchip.pong.game.clock  = io_in[12];
	assign \mchip.pong.game.left_movedir  = \mchip.pong.sync.o_out [7];
	assign \mchip.pong.game.left_paddle.Cnewgame  = \mchip.pong.game.ball.cpath.state [0];
	assign \mchip.pong.game.left_paddle.clock  = io_in[12];
	assign \mchip.pong.game.left_paddle.movedir_input  = \mchip.pong.sync.o_out [7];
	assign \mchip.pong.game.paddleLY  = \mchip.pong.game.left_paddle.coord ;
	assign \mchip.pong.game.paddleRY  = \mchip.pong.game.right_paddle.coord ;
	assign \mchip.pong.game.renderer.ball.color  = 24'h000000;
	assign \mchip.pong.game.renderer.ball1.color  = 24'h000000;
	assign \mchip.pong.game.renderer.ball2.color  = 24'h000000;
	assign \mchip.pong.game.renderer.ballX  = {\mchip.pong.game.ball.dpath.ballX [9:1], 1'h0};
	assign \mchip.pong.game.renderer.ballY  = \mchip.pong.game.ball.dpath.ballY ;
	assign \mchip.pong.game.renderer.ballrom_out  = 24'h000000;
	assign \mchip.pong.game.renderer.ballrom_out0  = 24'h000000;
	assign \mchip.pong.game.renderer.ballrom_out1  = 24'h000000;
	assign \mchip.pong.game.renderer.ballrom_out2  = 24'h000000;
	assign \mchip.pong.game.renderer.cfg1  = \mchip.pong.sync.o_out [1];
	assign \mchip.pong.game.renderer.cfg2  = \mchip.pong.sync.o_out [0];
	assign \mchip.pong.game.renderer.paddleLY  = \mchip.pong.game.left_paddle.coord ;
	assign \mchip.pong.game.renderer.paddleRY  = \mchip.pong.game.right_paddle.coord ;
	assign \mchip.pong.game.renderer.vga_b  = {\mchip.pong.VGA_B3 , \mchip.pong.VGA_B2 , 6'h00};
	assign \mchip.pong.game.renderer.vga_col  = {6'h00, \mchip.pong.game.vga.pix_ind [3:0]};
	assign \mchip.pong.game.renderer.vga_g  = {\mchip.pong.VGA_G3 , \mchip.pong.VGA_G2 , 6'h00};
	assign \mchip.pong.game.renderer.vga_r  = {\mchip.pong.VGA_R3 , \mchip.pong.VGA_R2 , 6'h00};
	assign \mchip.pong.game.reset  = \mchip.pong.sync.o_out [2];
	assign \mchip.pong.game.right_movedir  = \mchip.pong.sync.o_out [5];
	assign \mchip.pong.game.right_paddle.Cnewgame  = \mchip.pong.game.ball.cpath.state [0];
	assign \mchip.pong.game.right_paddle.clock  = io_in[12];
	assign \mchip.pong.game.right_paddle.movedir_input  = \mchip.pong.sync.o_out [5];
	assign \mchip.pong.game.score.Cnewgame  = \mchip.pong.game.ball.cpath.state [0];
	assign \mchip.pong.game.score.clock  = io_in[12];
	assign \mchip.pong.game.score.lscore_adder.B  = 16'h0001;
	assign \mchip.pong.game.score.lscore_adder.add0.B  = 4'h1;
	assign \mchip.pong.game.score.lscore_adder.add0.Cin  = 1'h0;
	assign \mchip.pong.game.score.lscore_adder.add1.B  = 4'h0;
	assign \mchip.pong.game.score.lscore_adder.add2.B  = 4'h0;
	assign \mchip.pong.game.score.lscore_adder.add3.B  = 4'h0;
	assign \mchip.pong.game.score.rscore_adder.B  = 16'h0001;
	assign \mchip.pong.game.score.rscore_adder.add0.B  = 4'h1;
	assign \mchip.pong.game.score.rscore_adder.add0.Cin  = 1'h0;
	assign \mchip.pong.game.score.rscore_adder.add1.B  = 4'h0;
	assign \mchip.pong.game.score.rscore_adder.add2.B  = 4'h0;
	assign \mchip.pong.game.score.rscore_adder.add3.B  = 4'h0;
	assign \mchip.pong.game.serve_input  = \mchip.pong.sync.o_out [3];
	assign \mchip.pong.game.tick.clock  = io_in[12];
	assign \mchip.pong.game.tick.col  = {6'h00, \mchip.pong.game.vga.pix_ind [3:0]};
	assign \mchip.pong.game.vga.HS  = \mchip.pong.VGA_HS ;
	assign \mchip.pong.game.vga.VS  = \mchip.pong.VGA_VS ;
	assign \mchip.pong.game.vga.clock  = io_in[12];
	assign \mchip.pong.game.vga.col  = {6'h00, \mchip.pong.game.vga.pix_ind [3:0]};
	assign \mchip.pong.game.vga.reset  = \mchip.pong.sync.o_out [2];
	assign \mchip.pong.game.vga_col  = {6'h00, \mchip.pong.game.vga.pix_ind [3:0]};
	assign \mchip.pong.left_down  = \mchip.pong.sync.o_out [6];
	assign \mchip.pong.left_up  = \mchip.pong.sync.o_out [7];
	assign \mchip.pong.right_down  = \mchip.pong.sync.o_out [4];
	assign \mchip.pong.right_up  = \mchip.pong.sync.o_out [5];
	assign \mchip.pong.rst  = \mchip.pong.sync.o_out [2];
	assign \mchip.pong.serve  = \mchip.pong.sync.o_out [3];
	assign \mchip.pong.sync.i_clk  = io_in[12];
	assign \mchip.pong.sync.i_in  = {io_in[3:0], io_in[5:4], io_in[7:6]};
	assign \mchip.pong.sync.i_rst  = 1'h0;
	assign \mchip.reset  = io_in[13];
endmodule
module d07_demo_vgarunner (
	io_in,
	io_out
);
	wire [6:0] _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire _2025_;
	wire _2026_;
	wire _2027_;
	wire _2028_;
	wire _2029_;
	wire _2030_;
	wire _2031_;
	wire _2032_;
	wire _2033_;
	wire _2034_;
	wire _2035_;
	wire _2036_;
	wire _2037_;
	wire _2038_;
	wire _2039_;
	wire _2040_;
	wire _2041_;
	wire _2042_;
	wire _2043_;
	wire _2044_;
	wire _2045_;
	wire _2046_;
	wire _2047_;
	wire _2048_;
	wire _2049_;
	wire _2050_;
	wire _2051_;
	wire _2052_;
	wire _2053_;
	wire _2054_;
	wire _2055_;
	wire _2056_;
	wire _2057_;
	wire _2058_;
	wire _2059_;
	wire _2060_;
	wire _2061_;
	wire _2062_;
	wire _2063_;
	wire _2064_;
	wire _2065_;
	wire _2066_;
	wire _2067_;
	wire _2068_;
	wire _2069_;
	wire _2070_;
	wire _2071_;
	wire _2072_;
	wire _2073_;
	wire _2074_;
	wire _2075_;
	wire _2076_;
	wire _2077_;
	wire _2078_;
	wire _2079_;
	wire _2080_;
	wire _2081_;
	wire _2082_;
	wire _2083_;
	wire _2084_;
	wire _2085_;
	wire _2086_;
	wire _2087_;
	wire _2088_;
	wire _2089_;
	wire _2090_;
	wire _2091_;
	wire _2092_;
	wire _2093_;
	wire _2094_;
	wire _2095_;
	wire _2096_;
	wire _2097_;
	wire _2098_;
	wire _2099_;
	wire _2100_;
	wire _2101_;
	wire _2102_;
	wire _2103_;
	wire _2104_;
	wire _2105_;
	wire _2106_;
	wire _2107_;
	wire _2108_;
	wire _2109_;
	wire _2110_;
	wire _2111_;
	wire _2112_;
	wire _2113_;
	wire _2114_;
	wire _2115_;
	wire _2116_;
	wire _2117_;
	wire _2118_;
	wire _2119_;
	wire _2120_;
	wire _2121_;
	wire _2122_;
	wire _2123_;
	wire _2124_;
	wire _2125_;
	wire _2126_;
	wire _2127_;
	wire _2128_;
	wire _2129_;
	wire _2130_;
	wire _2131_;
	wire _2132_;
	wire _2133_;
	wire _2134_;
	wire _2135_;
	wire _2136_;
	wire _2137_;
	wire _2138_;
	wire _2139_;
	wire _2140_;
	wire _2141_;
	wire _2142_;
	wire _2143_;
	wire _2144_;
	wire _2145_;
	wire _2146_;
	wire _2147_;
	wire _2148_;
	wire _2149_;
	wire _2150_;
	wire _2151_;
	wire _2152_;
	wire _2153_;
	wire _2154_;
	wire _2155_;
	wire _2156_;
	wire _2157_;
	wire _2158_;
	wire _2159_;
	wire _2160_;
	wire _2161_;
	wire _2162_;
	wire _2163_;
	wire _2164_;
	wire _2165_;
	wire _2166_;
	wire _2167_;
	wire _2168_;
	wire _2169_;
	wire _2170_;
	wire _2171_;
	wire _2172_;
	wire _2173_;
	wire _2174_;
	wire _2175_;
	wire _2176_;
	wire _2177_;
	wire _2178_;
	wire _2179_;
	wire _2180_;
	wire _2181_;
	wire _2182_;
	wire _2183_;
	wire _2184_;
	wire _2185_;
	wire _2186_;
	wire _2187_;
	wire _2188_;
	wire _2189_;
	wire _2190_;
	wire _2191_;
	wire _2192_;
	wire _2193_;
	wire _2194_;
	wire _2195_;
	wire _2196_;
	wire _2197_;
	wire _2198_;
	wire _2199_;
	wire _2200_;
	wire _2201_;
	wire _2202_;
	wire _2203_;
	wire _2204_;
	wire _2205_;
	wire _2206_;
	wire _2207_;
	wire _2208_;
	wire _2209_;
	wire _2210_;
	wire _2211_;
	wire _2212_;
	wire _2213_;
	wire _2214_;
	wire _2215_;
	wire _2216_;
	wire _2217_;
	wire _2218_;
	wire _2219_;
	wire _2220_;
	wire _2221_;
	wire _2222_;
	wire _2223_;
	wire _2224_;
	wire _2225_;
	wire _2226_;
	wire _2227_;
	wire _2228_;
	wire _2229_;
	wire _2230_;
	wire _2231_;
	wire _2232_;
	wire _2233_;
	wire _2234_;
	wire _2235_;
	wire _2236_;
	wire _2237_;
	wire _2238_;
	wire _2239_;
	wire _2240_;
	wire _2241_;
	wire _2242_;
	wire _2243_;
	wire _2244_;
	wire _2245_;
	wire _2246_;
	wire _2247_;
	wire _2248_;
	wire _2249_;
	wire _2250_;
	wire _2251_;
	wire _2252_;
	wire _2253_;
	wire _2254_;
	wire _2255_;
	wire _2256_;
	wire _2257_;
	wire _2258_;
	wire _2259_;
	wire _2260_;
	wire _2261_;
	wire _2262_;
	wire _2263_;
	wire _2264_;
	wire _2265_;
	wire _2266_;
	wire _2267_;
	wire _2268_;
	wire _2269_;
	wire _2270_;
	wire _2271_;
	wire _2272_;
	wire _2273_;
	wire _2274_;
	wire _2275_;
	wire _2276_;
	wire _2277_;
	wire _2278_;
	wire _2279_;
	wire _2280_;
	wire _2281_;
	wire _2282_;
	wire _2283_;
	wire _2284_;
	wire _2285_;
	wire _2286_;
	wire _2287_;
	wire _2288_;
	wire _2289_;
	wire _2290_;
	wire _2291_;
	wire _2292_;
	wire _2293_;
	wire _2294_;
	wire _2295_;
	wire _2296_;
	wire _2297_;
	wire _2298_;
	wire _2299_;
	wire _2300_;
	wire _2301_;
	wire _2302_;
	wire _2303_;
	wire _2304_;
	wire _2305_;
	wire _2306_;
	wire _2307_;
	wire _2308_;
	wire _2309_;
	wire _2310_;
	wire _2311_;
	wire _2312_;
	wire _2313_;
	wire _2314_;
	wire _2315_;
	wire _2316_;
	wire _2317_;
	wire _2318_;
	wire _2319_;
	wire _2320_;
	wire _2321_;
	wire _2322_;
	wire _2323_;
	wire _2324_;
	wire _2325_;
	wire _2326_;
	wire _2327_;
	wire _2328_;
	wire _2329_;
	wire _2330_;
	wire _2331_;
	wire _2332_;
	wire _2333_;
	wire _2334_;
	wire _2335_;
	wire _2336_;
	wire _2337_;
	wire _2338_;
	wire _2339_;
	wire _2340_;
	wire _2341_;
	wire _2342_;
	wire _2343_;
	wire _2344_;
	wire _2345_;
	wire _2346_;
	wire _2347_;
	wire _2348_;
	wire _2349_;
	wire _2350_;
	wire _2351_;
	wire _2352_;
	wire _2353_;
	wire _2354_;
	wire _2355_;
	wire _2356_;
	wire _2357_;
	wire _2358_;
	wire _2359_;
	wire _2360_;
	wire _2361_;
	wire _2362_;
	wire _2363_;
	wire _2364_;
	wire _2365_;
	wire _2366_;
	wire _2367_;
	wire _2368_;
	wire _2369_;
	wire _2370_;
	wire _2371_;
	wire _2372_;
	wire _2373_;
	wire _2374_;
	wire _2375_;
	wire _2376_;
	wire _2377_;
	wire _2378_;
	wire _2379_;
	wire _2380_;
	wire _2381_;
	wire _2382_;
	wire _2383_;
	wire _2384_;
	wire _2385_;
	wire _2386_;
	wire _2387_;
	wire _2388_;
	wire _2389_;
	wire _2390_;
	wire _2391_;
	wire _2392_;
	wire _2393_;
	wire _2394_;
	wire _2395_;
	wire _2396_;
	wire _2397_;
	wire _2398_;
	wire _2399_;
	wire _2400_;
	wire _2401_;
	wire _2402_;
	wire _2403_;
	wire _2404_;
	wire _2405_;
	wire _2406_;
	wire _2407_;
	wire _2408_;
	wire _2409_;
	wire _2410_;
	wire _2411_;
	wire _2412_;
	wire _2413_;
	wire _2414_;
	wire _2415_;
	wire _2416_;
	wire _2417_;
	wire _2418_;
	wire _2419_;
	wire _2420_;
	wire _2421_;
	wire _2422_;
	wire _2423_;
	wire _2424_;
	wire _2425_;
	wire _2426_;
	wire _2427_;
	wire _2428_;
	wire _2429_;
	wire _2430_;
	wire _2431_;
	wire _2432_;
	wire _2433_;
	wire _2434_;
	wire _2435_;
	wire _2436_;
	wire _2437_;
	wire _2438_;
	wire _2439_;
	wire _2440_;
	wire _2441_;
	wire _2442_;
	wire _2443_;
	wire _2444_;
	wire _2445_;
	wire _2446_;
	wire _2447_;
	wire _2448_;
	wire _2449_;
	wire _2450_;
	wire _2451_;
	wire _2452_;
	wire _2453_;
	wire _2454_;
	wire _2455_;
	wire _2456_;
	wire _2457_;
	wire _2458_;
	wire _2459_;
	wire _2460_;
	wire _2461_;
	wire _2462_;
	wire _2463_;
	wire _2464_;
	wire _2465_;
	wire _2466_;
	wire _2467_;
	wire _2468_;
	wire _2469_;
	wire _2470_;
	wire _2471_;
	wire _2472_;
	wire _2473_;
	wire _2474_;
	wire _2475_;
	wire _2476_;
	wire _2477_;
	wire _2478_;
	wire _2479_;
	wire _2480_;
	wire _2481_;
	wire _2482_;
	wire _2483_;
	wire _2484_;
	wire _2485_;
	wire _2486_;
	wire _2487_;
	wire _2488_;
	wire _2489_;
	wire _2490_;
	wire _2491_;
	wire _2492_;
	wire _2493_;
	wire _2494_;
	wire _2495_;
	wire _2496_;
	wire _2497_;
	wire _2498_;
	wire _2499_;
	wire _2500_;
	wire _2501_;
	wire _2502_;
	wire _2503_;
	wire _2504_;
	wire _2505_;
	wire _2506_;
	wire _2507_;
	wire _2508_;
	wire _2509_;
	wire _2510_;
	wire _2511_;
	wire _2512_;
	wire _2513_;
	wire _2514_;
	wire _2515_;
	wire _2516_;
	wire _2517_;
	wire _2518_;
	wire _2519_;
	wire _2520_;
	wire _2521_;
	wire _2522_;
	wire _2523_;
	wire _2524_;
	wire _2525_;
	wire _2526_;
	wire _2527_;
	wire _2528_;
	wire _2529_;
	wire _2530_;
	wire _2531_;
	wire _2532_;
	wire _2533_;
	wire _2534_;
	wire _2535_;
	wire _2536_;
	wire _2537_;
	wire _2538_;
	wire _2539_;
	wire _2540_;
	wire _2541_;
	wire _2542_;
	wire _2543_;
	wire _2544_;
	wire _2545_;
	wire _2546_;
	wire _2547_;
	wire _2548_;
	wire _2549_;
	wire _2550_;
	wire _2551_;
	wire _2552_;
	wire _2553_;
	wire _2554_;
	wire _2555_;
	wire _2556_;
	wire _2557_;
	wire _2558_;
	wire _2559_;
	wire _2560_;
	wire _2561_;
	wire _2562_;
	wire _2563_;
	wire _2564_;
	wire _2565_;
	wire _2566_;
	wire _2567_;
	wire _2568_;
	wire _2569_;
	wire _2570_;
	wire _2571_;
	wire _2572_;
	wire _2573_;
	wire _2574_;
	wire _2575_;
	wire _2576_;
	wire _2577_;
	wire _2578_;
	wire _2579_;
	wire _2580_;
	wire _2581_;
	wire _2582_;
	wire _2583_;
	wire _2584_;
	wire _2585_;
	wire _2586_;
	wire _2587_;
	wire _2588_;
	wire _2589_;
	wire _2590_;
	wire _2591_;
	wire _2592_;
	wire _2593_;
	wire _2594_;
	wire _2595_;
	wire _2596_;
	wire _2597_;
	wire _2598_;
	wire _2599_;
	wire _2600_;
	wire _2601_;
	wire _2602_;
	wire _2603_;
	wire _2604_;
	wire _2605_;
	wire _2606_;
	wire _2607_;
	wire _2608_;
	wire _2609_;
	wire _2610_;
	wire _2611_;
	wire _2612_;
	wire _2613_;
	wire _2614_;
	wire _2615_;
	wire _2616_;
	wire _2617_;
	wire _2618_;
	wire _2619_;
	wire _2620_;
	wire _2621_;
	wire _2622_;
	wire _2623_;
	wire _2624_;
	wire _2625_;
	wire _2626_;
	wire _2627_;
	wire _2628_;
	wire _2629_;
	wire _2630_;
	wire _2631_;
	wire _2632_;
	wire _2633_;
	wire _2634_;
	wire _2635_;
	wire _2636_;
	wire _2637_;
	wire _2638_;
	wire _2639_;
	wire _2640_;
	wire _2641_;
	wire _2642_;
	wire _2643_;
	wire _2644_;
	wire _2645_;
	wire _2646_;
	wire _2647_;
	wire _2648_;
	wire _2649_;
	wire _2650_;
	wire _2651_;
	wire _2652_;
	wire _2653_;
	wire _2654_;
	wire _2655_;
	wire _2656_;
	wire _2657_;
	wire _2658_;
	wire _2659_;
	wire _2660_;
	wire _2661_;
	wire _2662_;
	wire _2663_;
	wire _2664_;
	wire _2665_;
	wire _2666_;
	wire _2667_;
	wire _2668_;
	wire _2669_;
	wire _2670_;
	wire _2671_;
	wire _2672_;
	wire _2673_;
	wire _2674_;
	wire _2675_;
	wire _2676_;
	wire _2677_;
	wire _2678_;
	wire _2679_;
	wire _2680_;
	wire _2681_;
	wire _2682_;
	wire _2683_;
	wire _2684_;
	wire _2685_;
	wire _2686_;
	wire _2687_;
	wire _2688_;
	wire _2689_;
	wire _2690_;
	wire _2691_;
	wire _2692_;
	wire _2693_;
	wire _2694_;
	wire _2695_;
	wire _2696_;
	wire _2697_;
	wire _2698_;
	wire _2699_;
	wire _2700_;
	wire _2701_;
	wire _2702_;
	wire _2703_;
	wire _2704_;
	wire _2705_;
	wire _2706_;
	wire _2707_;
	wire _2708_;
	wire _2709_;
	wire _2710_;
	wire _2711_;
	wire _2712_;
	wire _2713_;
	wire _2714_;
	wire _2715_;
	wire _2716_;
	wire _2717_;
	wire _2718_;
	wire _2719_;
	wire _2720_;
	wire _2721_;
	wire _2722_;
	wire _2723_;
	wire _2724_;
	wire _2725_;
	wire _2726_;
	wire _2727_;
	wire _2728_;
	wire _2729_;
	wire _2730_;
	wire _2731_;
	wire _2732_;
	wire _2733_;
	wire _2734_;
	wire _2735_;
	wire _2736_;
	wire _2737_;
	wire _2738_;
	wire _2739_;
	wire _2740_;
	wire _2741_;
	wire _2742_;
	wire _2743_;
	wire _2744_;
	wire _2745_;
	wire _2746_;
	wire _2747_;
	wire _2748_;
	wire _2749_;
	wire _2750_;
	wire _2751_;
	wire _2752_;
	wire _2753_;
	wire _2754_;
	wire _2755_;
	wire _2756_;
	wire _2757_;
	wire _2758_;
	wire _2759_;
	wire _2760_;
	wire _2761_;
	wire _2762_;
	wire _2763_;
	wire _2764_;
	wire _2765_;
	wire _2766_;
	wire _2767_;
	wire _2768_;
	wire _2769_;
	wire _2770_;
	wire _2771_;
	wire _2772_;
	wire _2773_;
	wire _2774_;
	wire _2775_;
	wire _2776_;
	wire _2777_;
	wire _2778_;
	wire _2779_;
	wire _2780_;
	wire _2781_;
	wire _2782_;
	wire _2783_;
	wire _2784_;
	wire _2785_;
	wire _2786_;
	wire _2787_;
	wire _2788_;
	wire _2789_;
	wire _2790_;
	wire _2791_;
	wire _2792_;
	wire _2793_;
	wire _2794_;
	wire _2795_;
	wire _2796_;
	wire _2797_;
	wire _2798_;
	wire _2799_;
	wire _2800_;
	wire _2801_;
	wire _2802_;
	wire _2803_;
	wire _2804_;
	wire _2805_;
	wire _2806_;
	wire _2807_;
	wire _2808_;
	wire _2809_;
	wire _2810_;
	wire _2811_;
	wire _2812_;
	wire _2813_;
	wire _2814_;
	wire _2815_;
	wire _2816_;
	wire _2817_;
	wire _2818_;
	wire _2819_;
	wire _2820_;
	wire _2821_;
	wire _2822_;
	wire _2823_;
	wire _2824_;
	wire _2825_;
	wire _2826_;
	wire _2827_;
	wire _2828_;
	wire _2829_;
	wire _2830_;
	wire _2831_;
	wire _2832_;
	wire _2833_;
	wire _2834_;
	wire _2835_;
	wire _2836_;
	wire _2837_;
	wire _2838_;
	wire _2839_;
	wire _2840_;
	wire _2841_;
	wire _2842_;
	wire _2843_;
	wire _2844_;
	wire _2845_;
	wire _2846_;
	wire _2847_;
	wire _2848_;
	wire _2849_;
	wire _2850_;
	wire _2851_;
	wire _2852_;
	wire _2853_;
	wire _2854_;
	wire _2855_;
	wire _2856_;
	wire _2857_;
	wire _2858_;
	wire _2859_;
	wire _2860_;
	wire _2861_;
	wire _2862_;
	wire _2863_;
	wire _2864_;
	wire _2865_;
	wire _2866_;
	wire _2867_;
	wire _2868_;
	wire _2869_;
	wire _2870_;
	wire _2871_;
	wire _2872_;
	wire _2873_;
	wire _2874_;
	wire _2875_;
	wire _2876_;
	wire _2877_;
	wire _2878_;
	wire _2879_;
	wire _2880_;
	wire _2881_;
	wire _2882_;
	wire _2883_;
	wire _2884_;
	wire _2885_;
	wire _2886_;
	wire _2887_;
	wire _2888_;
	wire _2889_;
	wire _2890_;
	wire _2891_;
	wire _2892_;
	wire _2893_;
	wire _2894_;
	wire _2895_;
	wire _2896_;
	wire _2897_;
	wire _2898_;
	wire _2899_;
	wire _2900_;
	wire _2901_;
	wire _2902_;
	wire _2903_;
	wire _2904_;
	wire _2905_;
	wire _2906_;
	wire _2907_;
	wire _2908_;
	wire _2909_;
	wire _2910_;
	wire _2911_;
	wire _2912_;
	wire _2913_;
	wire _2914_;
	wire _2915_;
	wire _2916_;
	wire _2917_;
	wire _2918_;
	wire _2919_;
	wire _2920_;
	wire _2921_;
	wire _2922_;
	wire _2923_;
	wire _2924_;
	wire _2925_;
	wire _2926_;
	wire _2927_;
	wire _2928_;
	wire _2929_;
	wire _2930_;
	wire _2931_;
	wire _2932_;
	wire _2933_;
	wire _2934_;
	wire _2935_;
	wire _2936_;
	wire _2937_;
	wire _2938_;
	wire _2939_;
	wire _2940_;
	wire _2941_;
	wire _2942_;
	wire _2943_;
	wire _2944_;
	wire _2945_;
	wire _2946_;
	wire _2947_;
	wire _2948_;
	wire _2949_;
	wire _2950_;
	wire _2951_;
	wire _2952_;
	wire _2953_;
	wire _2954_;
	wire _2955_;
	wire _2956_;
	wire _2957_;
	wire _2958_;
	wire _2959_;
	wire _2960_;
	wire _2961_;
	wire _2962_;
	wire _2963_;
	wire _2964_;
	wire _2965_;
	wire _2966_;
	wire _2967_;
	wire _2968_;
	wire _2969_;
	wire _2970_;
	wire _2971_;
	wire _2972_;
	wire _2973_;
	wire _2974_;
	wire _2975_;
	wire _2976_;
	wire _2977_;
	wire _2978_;
	wire _2979_;
	wire _2980_;
	wire _2981_;
	wire _2982_;
	wire _2983_;
	wire _2984_;
	wire _2985_;
	wire _2986_;
	wire _2987_;
	wire _2988_;
	wire _2989_;
	wire _2990_;
	wire _2991_;
	wire _2992_;
	wire _2993_;
	wire _2994_;
	wire _2995_;
	wire _2996_;
	wire _2997_;
	wire _2998_;
	wire _2999_;
	wire _3000_;
	wire _3001_;
	wire _3002_;
	wire _3003_;
	wire _3004_;
	wire _3005_;
	wire _3006_;
	wire _3007_;
	wire _3008_;
	wire _3009_;
	wire _3010_;
	wire _3011_;
	wire _3012_;
	wire _3013_;
	wire _3014_;
	wire _3015_;
	wire _3016_;
	wire _3017_;
	wire _3018_;
	wire _3019_;
	wire _3020_;
	wire _3021_;
	wire _3022_;
	wire _3023_;
	wire _3024_;
	wire _3025_;
	wire _3026_;
	wire _3027_;
	wire _3028_;
	wire _3029_;
	wire _3030_;
	wire _3031_;
	wire _3032_;
	wire _3033_;
	wire _3034_;
	wire _3035_;
	wire _3036_;
	wire _3037_;
	wire _3038_;
	wire _3039_;
	wire _3040_;
	wire _3041_;
	wire _3042_;
	wire _3043_;
	wire _3044_;
	wire _3045_;
	wire _3046_;
	wire _3047_;
	wire _3048_;
	wire _3049_;
	wire _3050_;
	wire _3051_;
	wire _3052_;
	wire _3053_;
	wire _3054_;
	wire _3055_;
	wire _3056_;
	wire _3057_;
	wire _3058_;
	wire _3059_;
	wire _3060_;
	wire _3061_;
	wire _3062_;
	wire _3063_;
	wire _3064_;
	wire _3065_;
	wire _3066_;
	wire _3067_;
	wire _3068_;
	wire _3069_;
	wire _3070_;
	wire _3071_;
	wire _3072_;
	wire _3073_;
	wire _3074_;
	wire _3075_;
	wire _3076_;
	wire _3077_;
	wire _3078_;
	wire _3079_;
	wire _3080_;
	wire _3081_;
	wire _3082_;
	wire _3083_;
	wire _3084_;
	wire _3085_;
	wire _3086_;
	wire _3087_;
	wire _3088_;
	wire _3089_;
	wire _3090_;
	wire _3091_;
	wire _3092_;
	wire _3093_;
	wire _3094_;
	wire _3095_;
	wire _3096_;
	wire _3097_;
	wire _3098_;
	wire _3099_;
	wire _3100_;
	wire _3101_;
	wire _3102_;
	wire _3103_;
	wire _3104_;
	wire _3105_;
	wire _3106_;
	wire _3107_;
	wire _3108_;
	wire _3109_;
	wire _3110_;
	wire _3111_;
	wire _3112_;
	wire _3113_;
	wire _3114_;
	wire _3115_;
	wire _3116_;
	wire _3117_;
	wire _3118_;
	wire _3119_;
	wire _3120_;
	wire _3121_;
	wire _3122_;
	wire _3123_;
	wire _3124_;
	wire _3125_;
	wire _3126_;
	wire _3127_;
	wire _3128_;
	wire _3129_;
	wire _3130_;
	wire _3131_;
	wire _3132_;
	wire _3133_;
	wire _3134_;
	wire _3135_;
	wire _3136_;
	wire _3137_;
	wire _3138_;
	wire _3139_;
	wire _3140_;
	wire _3141_;
	wire _3142_;
	wire _3143_;
	wire _3144_;
	wire _3145_;
	wire _3146_;
	wire _3147_;
	wire _3148_;
	wire _3149_;
	wire _3150_;
	wire _3151_;
	wire _3152_;
	wire _3153_;
	wire _3154_;
	wire _3155_;
	wire _3156_;
	wire _3157_;
	wire _3158_;
	wire _3159_;
	wire _3160_;
	wire _3161_;
	wire _3162_;
	wire _3163_;
	wire _3164_;
	wire _3165_;
	wire _3166_;
	wire _3167_;
	wire _3168_;
	wire _3169_;
	wire _3170_;
	wire _3171_;
	wire _3172_;
	wire _3173_;
	wire _3174_;
	wire _3175_;
	wire _3176_;
	wire _3177_;
	wire _3178_;
	wire _3179_;
	wire _3180_;
	wire _3181_;
	wire _3182_;
	wire _3183_;
	wire _3184_;
	wire _3185_;
	wire _3186_;
	wire _3187_;
	wire _3188_;
	wire _3189_;
	wire _3190_;
	wire _3191_;
	wire _3192_;
	wire _3193_;
	wire _3194_;
	wire _3195_;
	wire _3196_;
	wire _3197_;
	wire _3198_;
	wire _3199_;
	wire _3200_;
	wire _3201_;
	wire _3202_;
	wire _3203_;
	wire _3204_;
	wire _3205_;
	wire _3206_;
	wire _3207_;
	wire _3208_;
	wire _3209_;
	wire _3210_;
	wire _3211_;
	wire _3212_;
	wire _3213_;
	wire _3214_;
	wire _3215_;
	wire _3216_;
	wire _3217_;
	wire _3218_;
	wire _3219_;
	wire _3220_;
	wire _3221_;
	wire _3222_;
	wire _3223_;
	wire _3224_;
	wire _3225_;
	wire _3226_;
	wire _3227_;
	wire _3228_;
	wire _3229_;
	wire _3230_;
	wire _3231_;
	wire _3232_;
	wire _3233_;
	wire _3234_;
	wire _3235_;
	wire _3236_;
	wire _3237_;
	wire _3238_;
	wire _3239_;
	wire _3240_;
	wire _3241_;
	wire _3242_;
	wire _3243_;
	wire _3244_;
	wire _3245_;
	wire _3246_;
	wire _3247_;
	wire _3248_;
	wire _3249_;
	wire _3250_;
	wire _3251_;
	wire _3252_;
	wire _3253_;
	wire _3254_;
	wire _3255_;
	wire _3256_;
	wire _3257_;
	wire _3258_;
	wire _3259_;
	wire _3260_;
	wire _3261_;
	wire _3262_;
	wire _3263_;
	wire _3264_;
	wire _3265_;
	wire _3266_;
	wire _3267_;
	wire _3268_;
	wire _3269_;
	wire _3270_;
	wire _3271_;
	wire _3272_;
	wire _3273_;
	wire _3274_;
	wire _3275_;
	wire _3276_;
	wire _3277_;
	wire _3278_;
	wire _3279_;
	wire _3280_;
	wire _3281_;
	wire _3282_;
	wire _3283_;
	wire _3284_;
	wire _3285_;
	wire _3286_;
	wire _3287_;
	wire _3288_;
	wire _3289_;
	wire _3290_;
	wire _3291_;
	wire _3292_;
	wire _3293_;
	wire _3294_;
	wire _3295_;
	wire _3296_;
	wire _3297_;
	wire _3298_;
	wire _3299_;
	wire _3300_;
	wire _3301_;
	wire _3302_;
	wire _3303_;
	wire _3304_;
	wire _3305_;
	wire _3306_;
	wire _3307_;
	wire _3308_;
	wire _3309_;
	wire _3310_;
	wire _3311_;
	wire _3312_;
	wire _3313_;
	wire _3314_;
	wire _3315_;
	wire _3316_;
	wire _3317_;
	wire _3318_;
	wire _3319_;
	wire _3320_;
	wire _3321_;
	wire _3322_;
	wire _3323_;
	wire _3324_;
	wire _3325_;
	wire _3326_;
	wire _3327_;
	wire _3328_;
	wire _3329_;
	wire _3330_;
	wire _3331_;
	wire _3332_;
	wire _3333_;
	wire _3334_;
	wire _3335_;
	wire _3336_;
	wire _3337_;
	wire _3338_;
	wire _3339_;
	wire _3340_;
	wire _3341_;
	wire _3342_;
	wire _3343_;
	wire _3344_;
	wire _3345_;
	wire _3346_;
	wire _3347_;
	wire _3348_;
	wire _3349_;
	wire _3350_;
	wire _3351_;
	wire _3352_;
	wire _3353_;
	wire _3354_;
	wire _3355_;
	wire _3356_;
	wire _3357_;
	wire _3358_;
	wire _3359_;
	wire _3360_;
	wire _3361_;
	wire _3362_;
	wire _3363_;
	wire _3364_;
	wire _3365_;
	wire _3366_;
	wire _3367_;
	wire _3368_;
	wire _3369_;
	wire _3370_;
	wire _3371_;
	wire _3372_;
	wire _3373_;
	wire _3374_;
	wire _3375_;
	wire _3376_;
	wire _3377_;
	wire _3378_;
	wire _3379_;
	wire _3380_;
	wire _3381_;
	wire _3382_;
	wire _3383_;
	wire _3384_;
	wire _3385_;
	wire _3386_;
	wire _3387_;
	wire _3388_;
	wire _3389_;
	wire _3390_;
	wire _3391_;
	wire _3392_;
	wire _3393_;
	wire _3394_;
	wire _3395_;
	wire _3396_;
	wire _3397_;
	wire _3398_;
	wire _3399_;
	wire _3400_;
	wire _3401_;
	wire _3402_;
	wire _3403_;
	wire _3404_;
	wire _3405_;
	wire _3406_;
	wire _3407_;
	wire _3408_;
	wire _3409_;
	wire _3410_;
	wire _3411_;
	wire _3412_;
	wire _3413_;
	wire _3414_;
	wire _3415_;
	wire _3416_;
	wire _3417_;
	wire _3418_;
	wire _3419_;
	wire _3420_;
	wire _3421_;
	wire _3422_;
	wire _3423_;
	wire _3424_;
	wire _3425_;
	wire _3426_;
	wire _3427_;
	wire _3428_;
	wire _3429_;
	wire _3430_;
	wire _3431_;
	wire _3432_;
	wire _3433_;
	wire _3434_;
	wire _3435_;
	wire _3436_;
	wire _3437_;
	wire _3438_;
	wire _3439_;
	wire _3440_;
	wire _3441_;
	wire _3442_;
	wire _3443_;
	wire _3444_;
	wire _3445_;
	wire _3446_;
	wire _3447_;
	wire _3448_;
	wire _3449_;
	wire _3450_;
	wire _3451_;
	wire _3452_;
	wire _3453_;
	wire _3454_;
	wire _3455_;
	wire _3456_;
	wire _3457_;
	wire _3458_;
	wire _3459_;
	wire _3460_;
	wire _3461_;
	wire _3462_;
	wire _3463_;
	wire _3464_;
	wire _3465_;
	wire _3466_;
	wire _3467_;
	wire _3468_;
	wire _3469_;
	wire _3470_;
	wire _3471_;
	wire _3472_;
	wire _3473_;
	wire _3474_;
	wire _3475_;
	wire _3476_;
	wire _3477_;
	wire _3478_;
	wire _3479_;
	wire _3480_;
	wire _3481_;
	wire _3482_;
	wire _3483_;
	wire _3484_;
	wire _3485_;
	wire _3486_;
	wire _3487_;
	wire _3488_;
	wire _3489_;
	wire _3490_;
	wire _3491_;
	wire _3492_;
	wire _3493_;
	wire _3494_;
	wire _3495_;
	wire _3496_;
	wire _3497_;
	wire _3498_;
	wire _3499_;
	wire _3500_;
	wire _3501_;
	wire _3502_;
	wire _3503_;
	wire _3504_;
	wire _3505_;
	wire _3506_;
	wire _3507_;
	wire _3508_;
	wire _3509_;
	wire _3510_;
	wire _3511_;
	wire _3512_;
	wire _3513_;
	wire _3514_;
	wire _3515_;
	wire _3516_;
	wire _3517_;
	wire _3518_;
	wire _3519_;
	wire _3520_;
	wire _3521_;
	wire _3522_;
	wire _3523_;
	wire _3524_;
	wire _3525_;
	wire _3526_;
	wire _3527_;
	wire _3528_;
	wire _3529_;
	wire _3530_;
	wire _3531_;
	wire _3532_;
	wire _3533_;
	wire _3534_;
	wire _3535_;
	wire _3536_;
	wire _3537_;
	wire _3538_;
	wire _3539_;
	wire _3540_;
	wire _3541_;
	wire _3542_;
	wire _3543_;
	wire _3544_;
	wire _3545_;
	wire _3546_;
	wire _3547_;
	wire _3548_;
	wire _3549_;
	wire _3550_;
	wire _3551_;
	wire _3552_;
	wire _3553_;
	wire _3554_;
	wire _3555_;
	wire _3556_;
	wire _3557_;
	wire _3558_;
	wire _3559_;
	wire _3560_;
	wire _3561_;
	wire _3562_;
	wire _3563_;
	wire _3564_;
	wire _3565_;
	wire _3566_;
	wire _3567_;
	wire _3568_;
	wire _3569_;
	wire _3570_;
	wire _3571_;
	wire _3572_;
	wire _3573_;
	wire _3574_;
	wire _3575_;
	wire _3576_;
	wire _3577_;
	wire _3578_;
	wire _3579_;
	wire _3580_;
	wire _3581_;
	wire _3582_;
	wire _3583_;
	wire _3584_;
	wire _3585_;
	wire _3586_;
	wire _3587_;
	wire _3588_;
	wire _3589_;
	wire _3590_;
	wire _3591_;
	wire _3592_;
	wire _3593_;
	wire _3594_;
	wire _3595_;
	wire _3596_;
	wire _3597_;
	wire _3598_;
	wire _3599_;
	wire _3600_;
	wire _3601_;
	wire _3602_;
	wire _3603_;
	wire _3604_;
	wire _3605_;
	wire _3606_;
	wire _3607_;
	wire _3608_;
	wire _3609_;
	wire _3610_;
	wire _3611_;
	wire _3612_;
	wire _3613_;
	wire _3614_;
	wire _3615_;
	wire _3616_;
	wire _3617_;
	wire _3618_;
	wire _3619_;
	wire [9:0] _3620_;
	wire [19:0] _3621_;
	wire [31:0] _3622_;
	wire [19:0] _3623_;
	wire [31:0] _3624_;
	wire [9:0] _3625_;
	wire [10:0] _3626_;
	wire [10:0] _3627_;
	wire [17:0] _3628_;
	wire _3629_;
	wire _3630_;
	wire _3631_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [2:0] \mchip.game2.cactus_select ;
	reg [2:0] \mchip.game2.cactus_select_last ;
	reg [2:0] \mchip.game2.cactus_type ;
	wire \mchip.game2.clk ;
	wire \mchip.game2.dbg_pixel ;
	wire [15:0] \mchip.game2.dbg_score ;
	wire [10:0] \mchip.game2.dbg_scrolladdr ;
	wire [23:0] \mchip.game2.dbg_speed ;
	wire \mchip.game2.debug_in ;
	wire \mchip.game2.dinosprite_inst.clk ;
	reg [24:0] \mchip.game2.dinosprite_inst.ctr ;
	reg \mchip.game2.dinosprite_inst.sprite ;
	wire \mchip.game2.dinosprite_inst.sys_rst ;
	wire \mchip.game2.dinosprite_num ;
	reg \mchip.game2.game_over ;
	wire [9:0] \mchip.game2.haddr ;
	wire \mchip.game2.halt_in ;
	wire \mchip.game2.jump_in ;
	wire [6:0] \mchip.game2.jump_pos ;
	wire \mchip.game2.jumping_inst.clk ;
	reg [23:0] \mchip.game2.jumping_inst.ctr ;
	reg [8:0] \mchip.game2.jumping_inst.frame ;
	reg \mchip.game2.jumping_inst.in_air ;
	wire \mchip.game2.jumping_inst.jump ;
	reg [6:0] \mchip.game2.jumping_inst.jump_pos ;
	wire [23:0] \mchip.game2.jumping_inst.speed ;
	wire \mchip.game2.jumping_inst.sys_rst ;
	reg [19:0] \mchip.game2.no_jump_ctr ;
	wire [4:0] \mchip.game2.random ;
	reg [2:0] \mchip.game2.rendering_inst.cactus_select ;
	wire [2:0] \mchip.game2.rendering_inst.cactus_type ;
	wire \mchip.game2.rendering_inst.clk ;
	wire \mchip.game2.rendering_inst.dinosprite_num ;
	wire \mchip.game2.rendering_inst.game_over ;
	wire [9:0] \mchip.game2.rendering_inst.haddr ;
	wire [6:0] \mchip.game2.rendering_inst.jump_pos ;
	reg [4:0] \mchip.game2.rendering_inst.layers ;
	wire \mchip.game2.rendering_inst.pixel ;
	wire \mchip.game2.rendering_inst.score_pixel ;
	wire [10:0] \mchip.game2.rendering_inst.scrolladdr ;
	wire \mchip.game2.rendering_inst.sys_rst ;
	wire [9:0] \mchip.game2.rendering_inst.vaddr ;
	wire \mchip.game2.rng_inst.clk ;
	wire \mchip.game2.rng_inst.entropy_in ;
	reg [4:0] \mchip.game2.rng_inst.out ;
	wire \mchip.game2.rng_inst.sys_rst ;
	wire \mchip.game2.score_inst.clk ;
	reg [21:0] \mchip.game2.score_inst.ctr ;
	wire [9:0] \mchip.game2.score_inst.haddr ;
	reg \mchip.game2.score_inst.pixel ;
	reg [3:0] \mchip.game2.score_inst.score[0] ;
	reg [3:0] \mchip.game2.score_inst.score[1] ;
	reg [3:0] \mchip.game2.score_inst.score[2] ;
	reg [3:0] \mchip.game2.score_inst.score[3] ;
	wire [15:0] \mchip.game2.score_inst.score_out ;
	reg [3:0] \mchip.game2.score_inst.score_saved[0] ;
	reg [3:0] \mchip.game2.score_inst.score_saved[1] ;
	reg [3:0] \mchip.game2.score_inst.score_saved[2] ;
	reg [3:0] \mchip.game2.score_inst.score_saved[3] ;
	wire \mchip.game2.score_inst.sys_rst ;
	wire [9:0] \mchip.game2.score_inst.vaddr ;
	wire [15:0] \mchip.game2.score_out ;
	wire \mchip.game2.score_pixel ;
	wire \mchip.game2.scroll_inst.clk ;
	reg [17:0] \mchip.game2.scroll_inst.ctr ;
	wire [7:0] \mchip.game2.scroll_inst.move_amt ;
	reg [10:0] \mchip.game2.scroll_inst.pos ;
	wire [23:0] \mchip.game2.scroll_inst.speed ;
	wire [7:0] \mchip.game2.scroll_inst.speed_change ;
	wire \mchip.game2.scroll_inst.sys_rst ;
	reg [17:0] \mchip.game2.scroll_inst.tick_time ;
	wire [10:0] \mchip.game2.scrolladdr ;
	wire [23:0] \mchip.game2.speed ;
	reg [31:0] \mchip.game2.start_ctr ;
	wire \mchip.game2.sys_rst ;
	wire [9:0] \mchip.game2.vaddr ;
	wire [3:0] \mchip.game2.vga_blue ;
	wire [3:0] \mchip.game2.vga_green ;
	wire \mchip.game2.vga_hsync ;
	wire \mchip.game2.vga_inst.clk ;
	reg [9:0] \mchip.game2.vga_inst.haddr ;
	reg \mchip.game2.vga_inst.hsync ;
	wire \mchip.game2.vga_inst.sys_rst ;
	reg [9:0] \mchip.game2.vga_inst.vaddr ;
	reg \mchip.game2.vga_inst.vsync ;
	wire \mchip.game2.vga_pixel ;
	wire [3:0] \mchip.game2.vga_red ;
	wire \mchip.game2.vga_vsync ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _3171_ = io_in[11] & io_in[7];
	assign _3628_[0] = _3171_ ^ \mchip.game2.scroll_inst.tick_time [0];
	assign _3620_[0] = ~\mchip.game2.vga_inst.haddr [0];
	assign _3172_ = ~(\mchip.game2.vga_inst.haddr [8] & \mchip.game2.vga_inst.haddr [7]);
	assign _3173_ = \mchip.game2.vga_inst.haddr [8] & ~\mchip.game2.vga_inst.haddr [7];
	assign _3174_ = ~(\mchip.game2.vga_inst.haddr [6] | \mchip.game2.vga_inst.haddr [5]);
	assign _3175_ = _3173_ & ~_3174_;
	assign _3176_ = _3172_ & ~_3175_;
	assign _3177_ = \mchip.game2.vga_inst.haddr [9] & ~_3176_;
	assign _3178_ = \mchip.game2.vga_inst.haddr [5] & ~\mchip.game2.vga_inst.haddr [4];
	assign _3179_ = \mchip.game2.vga_inst.haddr [1] | \mchip.game2.vga_inst.haddr [0];
	assign _3180_ = _3178_ & ~_3179_;
	assign _3181_ = \mchip.game2.vga_inst.haddr [9] & \mchip.game2.vga_inst.haddr [8];
	assign _3182_ = ~(\mchip.game2.vga_inst.haddr [6] | \mchip.game2.vga_inst.haddr [7]);
	assign _3183_ = ~(_3182_ & _3181_);
	assign _3184_ = _3180_ & ~_3183_;
	assign _3185_ = ~(\mchip.game2.vga_inst.haddr [2] | \mchip.game2.vga_inst.haddr [3]);
	assign _3186_ = ~_3185_;
	assign _3187_ = _3184_ & ~_3186_;
	assign _0023_ = _3187_ | _3177_;
	assign _3188_ = ~(\mchip.game2.vga_inst.vaddr [8] | \mchip.game2.vga_inst.vaddr [9]);
	assign _3189_ = \mchip.game2.vga_inst.vaddr [1] & ~\mchip.game2.vga_inst.vaddr [0];
	assign _3190_ = \mchip.game2.vga_inst.vaddr [3] & ~\mchip.game2.vga_inst.vaddr [2];
	assign _3191_ = ~(_3190_ & _3189_);
	assign _3192_ = \mchip.game2.vga_inst.vaddr [6] & \mchip.game2.vga_inst.vaddr [7];
	assign _3193_ = \mchip.game2.vga_inst.vaddr [4] & \mchip.game2.vga_inst.vaddr [5];
	assign _3194_ = _3193_ & _3192_;
	assign _3195_ = _3191_ | ~_3194_;
	assign _3196_ = _3188_ & ~_3195_;
	assign _3197_ = ~_3188_;
	assign _3198_ = \mchip.game2.vga_inst.vaddr [0] & \mchip.game2.vga_inst.vaddr [1];
	assign _3199_ = _3190_ & ~_3198_;
	assign _3200_ = \mchip.game2.vga_inst.vaddr [3] & ~_3199_;
	assign _3201_ = _3194_ & ~_3200_;
	assign _3202_ = _3194_ & ~_3201_;
	assign _3203_ = _3202_ | _3197_;
	assign _3204_ = _3203_ | _3196_;
	assign _3205_ = _3192_ & _3188_;
	assign _3206_ = \mchip.game2.vga_inst.vaddr [2] & \mchip.game2.vga_inst.vaddr [3];
	assign _3207_ = ~(\mchip.game2.vga_inst.vaddr [4] | \mchip.game2.vga_inst.vaddr [5]);
	assign _3208_ = _3206_ | ~_3207_;
	assign _3209_ = _3205_ & ~_3208_;
	assign _3210_ = _3188_ & ~_3192_;
	assign _3211_ = _3210_ | _3209_;
	assign _3212_ = _3211_ | _3204_;
	assign _3213_ = \mchip.game2.vga_inst.vaddr [8] & ~\mchip.game2.vga_inst.vaddr [9];
	assign _3214_ = ~\mchip.game2.vga_inst.vaddr [5];
	assign _3215_ = _3192_ & ~_3214_;
	assign _3216_ = \mchip.game2.vga_inst.vaddr [4] | ~\mchip.game2.vga_inst.vaddr [5];
	assign _3217_ = _3216_ | ~_3192_;
	assign _3218_ = \mchip.game2.vga_inst.vaddr [2] | \mchip.game2.vga_inst.vaddr [3];
	assign _3219_ = ~(\mchip.game2.vga_inst.vaddr [0] | \mchip.game2.vga_inst.vaddr [1]);
	assign _3220_ = _3218_ | ~_3219_;
	assign _3221_ = ~(_3220_ | _3217_);
	assign _3222_ = _3215_ & ~_3221_;
	assign _3223_ = _3213_ & ~_3222_;
	assign _3224_ = _3223_ | _3188_;
	assign _3225_ = _3221_ & _3213_;
	assign _3226_ = _3224_ & ~_3225_;
	assign _3227_ = ~(\mchip.game2.vga_inst.haddr [8] | \mchip.game2.vga_inst.haddr [7]);
	assign _3228_ = \mchip.game2.vga_inst.haddr [9] & ~_3227_;
	assign _3229_ = _3226_ & ~_3228_;
	assign _3230_ = _3212_ | ~_3229_;
	assign _3231_ = io_in[13] | ~\mchip.game2.rendering_inst.cactus_select [0];
	assign _0015_ = _3231_ | _3230_;
	assign _3232_ = _3177_ & ~_3187_;
	assign _3233_ = _3232_ | io_in[13];
	assign _0013_ = _3233_ | _3187_;
	assign _3234_ = ~(\mchip.game2.start_ctr [24] | \mchip.game2.start_ctr [25]);
	assign _3235_ = \mchip.game2.start_ctr [26] | \mchip.game2.start_ctr [27];
	assign _3236_ = _3234_ & ~_3235_;
	assign _3237_ = \mchip.game2.start_ctr [29] | \mchip.game2.start_ctr [28];
	assign _3238_ = \mchip.game2.start_ctr [30] | \mchip.game2.start_ctr [31];
	assign _3239_ = _3238_ | _3237_;
	assign _3240_ = _3236_ & ~_3239_;
	assign _3241_ = \mchip.game2.start_ctr [25] | ~\mchip.game2.start_ctr [24];
	assign _3242_ = _3241_ | _3235_;
	assign _3243_ = ~(_3242_ | _3239_);
	assign _3244_ = \mchip.game2.start_ctr [22] & \mchip.game2.start_ctr [23];
	assign _3245_ = \mchip.game2.start_ctr [20] | \mchip.game2.start_ctr [21];
	assign _3246_ = _3244_ & ~_3245_;
	assign _3247_ = \mchip.game2.start_ctr [19] & ~\mchip.game2.start_ctr [18];
	assign _3248_ = \mchip.game2.start_ctr [17] | \mchip.game2.start_ctr [16];
	assign _3249_ = _3247_ & ~_3248_;
	assign _3250_ = \mchip.game2.start_ctr [19] & ~_3249_;
	assign _3251_ = _3246_ & ~_3250_;
	assign _3252_ = _3244_ & ~_3251_;
	assign _3253_ = _3243_ & ~_3252_;
	assign _3254_ = ~(_3253_ | _3240_);
	assign _3255_ = ~(\mchip.game2.start_ctr [15] & \mchip.game2.start_ctr [14]);
	assign _3256_ = \mchip.game2.start_ctr [12] | \mchip.game2.start_ctr [13];
	assign _3257_ = ~(_3256_ | _3255_);
	assign _3258_ = \mchip.game2.start_ctr [9] & \mchip.game2.start_ctr [8];
	assign _3259_ = \mchip.game2.start_ctr [10] | \mchip.game2.start_ctr [11];
	assign _3260_ = _3259_ | _3258_;
	assign _3261_ = _3257_ & ~_3260_;
	assign _3262_ = _3261_ | _3255_;
	assign _3263_ = \mchip.game2.start_ctr [7] & ~\mchip.game2.start_ctr [6];
	assign _3264_ = \mchip.game2.start_ctr [5] | \mchip.game2.start_ctr [4];
	assign _3265_ = _3263_ & ~_3264_;
	assign _3266_ = \mchip.game2.start_ctr [0] | \mchip.game2.start_ctr [1];
	assign _3267_ = \mchip.game2.start_ctr [2] | \mchip.game2.start_ctr [3];
	assign _3268_ = _3267_ | _3266_;
	assign _3269_ = _3265_ & ~_3268_;
	assign _3270_ = _3269_ | ~\mchip.game2.start_ctr [7];
	assign _3271_ = _3258_ & ~_3259_;
	assign _3272_ = ~(_3271_ & _3257_);
	assign _3273_ = _3270_ & ~_3272_;
	assign _3274_ = ~(_3273_ | _3262_);
	assign _3275_ = \mchip.game2.start_ctr [16] & ~\mchip.game2.start_ctr [17];
	assign _3276_ = _3275_ & _3247_;
	assign _3277_ = ~(_3276_ & _3246_);
	assign _3278_ = _3243_ & ~_3277_;
	assign _3279_ = _3278_ & ~_3274_;
	assign _3280_ = _3254_ & ~_3279_;
	assign _3281_ = _3272_ | ~_3269_;
	assign _3282_ = _3278_ & ~_3281_;
	assign _0162_ = ~(_3282_ | _3280_);
	assign _3283_ = ~(\mchip.game2.game_over  | io_in[1]);
	assign _0163_ = _3283_ & ~_0162_;
	assign _3284_ = \mchip.game2.score_inst.ctr [17] & ~\mchip.game2.score_inst.ctr [16];
	assign _3285_ = \mchip.game2.score_inst.ctr [19] | ~\mchip.game2.score_inst.ctr [18];
	assign _3286_ = _3285_ | ~_3284_;
	assign _3287_ = \mchip.game2.score_inst.ctr [20] | ~\mchip.game2.score_inst.ctr [21];
	assign _3288_ = _3287_ | _3286_;
	assign _3289_ = \mchip.game2.score_inst.ctr [13] & ~\mchip.game2.score_inst.ctr [12];
	assign _3290_ = \mchip.game2.score_inst.ctr [15] | ~\mchip.game2.score_inst.ctr [14];
	assign _3291_ = _3290_ | ~_3289_;
	assign _3292_ = \mchip.game2.score_inst.ctr [8] & ~\mchip.game2.score_inst.ctr [9];
	assign _3293_ = \mchip.game2.score_inst.ctr [10] | ~\mchip.game2.score_inst.ctr [11];
	assign _3294_ = _3293_ | ~_3292_;
	assign _3295_ = _3294_ | _3291_;
	assign _3296_ = ~(\mchip.game2.score_inst.ctr [4] & \mchip.game2.score_inst.ctr [5]);
	assign _3297_ = ~(\mchip.game2.score_inst.ctr [6] & \mchip.game2.score_inst.ctr [7]);
	assign _3298_ = _3297_ | _3296_;
	assign _3299_ = \mchip.game2.score_inst.ctr [0] | \mchip.game2.score_inst.ctr [1];
	assign _3300_ = ~(\mchip.game2.score_inst.ctr [2] & \mchip.game2.score_inst.ctr [3]);
	assign _3301_ = _3300_ | _3299_;
	assign _3302_ = _3301_ | _3298_;
	assign _3303_ = _3302_ | _3295_;
	assign _3304_ = _3303_ | _3288_;
	assign _3305_ = ~(_3287_ | _3285_);
	assign _3306_ = ~(\mchip.game2.score_inst.ctr [17] & \mchip.game2.score_inst.ctr [16]);
	assign _3307_ = ~\mchip.game2.score_inst.ctr [15];
	assign _3308_ = _3284_ & ~_3307_;
	assign _3309_ = _3306_ & ~_3308_;
	assign _3310_ = _3284_ & ~_3290_;
	assign _3311_ = ~(\mchip.game2.score_inst.ctr [12] & \mchip.game2.score_inst.ctr [13]);
	assign _3312_ = ~(\mchip.game2.score_inst.ctr [11] & \mchip.game2.score_inst.ctr [10]);
	assign _3313_ = _3289_ & ~_3312_;
	assign _3314_ = _3311_ & ~_3313_;
	assign _3315_ = _3310_ & ~_3314_;
	assign _3316_ = _3309_ & ~_3315_;
	assign _3317_ = _3293_ | ~_3289_;
	assign _3318_ = _3310_ & ~_3317_;
	assign _3319_ = ~\mchip.game2.score_inst.ctr [9];
	assign _3320_ = _3292_ & ~_3297_;
	assign _3321_ = _3300_ | _3296_;
	assign _3322_ = _3320_ & ~_3321_;
	assign _3323_ = _3319_ & ~_3322_;
	assign _3324_ = _3318_ & ~_3323_;
	assign _3325_ = _3316_ & ~_3324_;
	assign _3326_ = _3305_ & ~_3325_;
	assign _3327_ = \mchip.game2.score_inst.ctr [19] & ~_3287_;
	assign _3328_ = \mchip.game2.score_inst.ctr [20] & \mchip.game2.score_inst.ctr [21];
	assign _3329_ = _3328_ | _3327_;
	assign _3330_ = _3329_ | _3326_;
	assign _3331_ = _3304_ & ~_3330_;
	assign _0006_ = _0163_ & ~_3331_;
	assign _3332_ = \mchip.game2.score_inst.score[1] [1] & \mchip.game2.score_inst.score[1] [0];
	assign _3333_ = _3332_ & \mchip.game2.score_inst.score[1] [2];
	assign _3334_ = ~(_3333_ ^ \mchip.game2.score_inst.score[1] [3]);
	assign _3335_ = ~_3334_;
	assign _3336_ = \mchip.game2.score_inst.score[1] [0] | ~\mchip.game2.score_inst.score[1] [1];
	assign _3337_ = _3332_ ^ \mchip.game2.score_inst.score[1] [2];
	assign _3338_ = _3337_ | _3334_;
	assign _3339_ = _3336_ & ~_3338_;
	assign _3340_ = _3335_ & ~_3339_;
	assign _3341_ = ~(\mchip.game2.score_inst.score[1] [3] & \mchip.game2.score_inst.score[1] [2]);
	assign _3342_ = _3332_ & ~_3341_;
	assign _3343_ = _3342_ | _3340_;
	assign _3344_ = \mchip.game2.score_inst.score[1] [1] | ~\mchip.game2.score_inst.score[1] [0];
	assign _3345_ = _3344_ | _3338_;
	assign _3346_ = ~(_3345_ | _3342_);
	assign _3347_ = _3346_ | _3343_;
	assign _3348_ = \mchip.game2.score_inst.score[0] [1] & \mchip.game2.score_inst.score[0] [0];
	assign _3349_ = _3348_ & \mchip.game2.score_inst.score[0] [2];
	assign _3350_ = ~(_3349_ ^ \mchip.game2.score_inst.score[0] [3]);
	assign _3351_ = \mchip.game2.score_inst.score[0] [0] | ~\mchip.game2.score_inst.score[0] [1];
	assign _3352_ = _3348_ ^ \mchip.game2.score_inst.score[0] [2];
	assign _3353_ = _3352_ | _3350_;
	assign _3354_ = _3353_ | ~_3351_;
	assign _3355_ = _3354_ & ~_3350_;
	assign _3356_ = ~(\mchip.game2.score_inst.score[0] [3] & \mchip.game2.score_inst.score[0] [2]);
	assign _3357_ = _3348_ & ~_3356_;
	assign _3358_ = ~(_3357_ | _3355_);
	assign _3359_ = \mchip.game2.score_inst.score[0] [1] | ~\mchip.game2.score_inst.score[0] [0];
	assign _3360_ = _3359_ | _3353_;
	assign _3361_ = ~(_3360_ | _3357_);
	assign _3362_ = _3358_ & ~_3361_;
	assign _3363_ = _3362_ | ~_3347_;
	assign _0004_ = _0006_ & ~_3363_;
	assign _3364_ = \mchip.game2.score_inst.score[2] [1] & \mchip.game2.score_inst.score[2] [0];
	assign _3365_ = _3364_ & \mchip.game2.score_inst.score[2] [2];
	assign _3366_ = ~(_3365_ ^ \mchip.game2.score_inst.score[2] [3]);
	assign _3367_ = ~_3366_;
	assign _3368_ = \mchip.game2.score_inst.score[2] [0] | ~\mchip.game2.score_inst.score[2] [1];
	assign _3369_ = _3364_ ^ \mchip.game2.score_inst.score[2] [2];
	assign _3370_ = _3369_ | _3366_;
	assign _3371_ = _3368_ & ~_3370_;
	assign _3372_ = _3367_ & ~_3371_;
	assign _3373_ = ~(\mchip.game2.score_inst.score[2] [3] & \mchip.game2.score_inst.score[2] [2]);
	assign _3374_ = _3364_ & ~_3373_;
	assign _3375_ = _3374_ | _3372_;
	assign _3376_ = \mchip.game2.score_inst.score[2] [1] | ~\mchip.game2.score_inst.score[2] [0];
	assign _3377_ = _3376_ | _3370_;
	assign _3378_ = ~(_3377_ | _3374_);
	assign _3379_ = _3378_ | _3375_;
	assign _0003_ = _3379_ & _0004_;
	assign _3380_ = ~(\mchip.game2.rendering_inst.cactus_select [1] & \mchip.game2.cactus_type [1]);
	assign _3381_ = \mchip.game2.scroll_inst.pos [8] & \mchip.game2.vga_inst.haddr [8];
	assign _3382_ = \mchip.game2.scroll_inst.pos [7] & \mchip.game2.vga_inst.haddr [7];
	assign _3383_ = \mchip.game2.scroll_inst.pos [6] & \mchip.game2.vga_inst.haddr [6];
	assign _3384_ = \mchip.game2.scroll_inst.pos [7] ^ \mchip.game2.vga_inst.haddr [7];
	assign _3385_ = _3384_ & _3383_;
	assign _3386_ = _3385_ | _3382_;
	assign _3387_ = \mchip.game2.scroll_inst.pos [5] & \mchip.game2.vga_inst.haddr [5];
	assign _3388_ = \mchip.game2.scroll_inst.pos [4] & \mchip.game2.vga_inst.haddr [4];
	assign _3389_ = \mchip.game2.scroll_inst.pos [5] | \mchip.game2.vga_inst.haddr [5];
	assign _3390_ = _3389_ & ~_3387_;
	assign _3391_ = _3390_ & _3388_;
	assign _3392_ = ~(_3391_ | _3387_);
	assign _3393_ = \mchip.game2.scroll_inst.pos [6] ^ \mchip.game2.vga_inst.haddr [6];
	assign _3394_ = ~(_3393_ & _3384_);
	assign _3395_ = ~(_3394_ | _3392_);
	assign _3396_ = _3395_ | _3386_;
	assign _3397_ = \mchip.game2.scroll_inst.pos [3] & \mchip.game2.vga_inst.haddr [3];
	assign _3398_ = \mchip.game2.scroll_inst.pos [2] & \mchip.game2.vga_inst.haddr [2];
	assign _3399_ = ~_3398_;
	assign _3400_ = ~(\mchip.game2.scroll_inst.pos [3] | \mchip.game2.vga_inst.haddr [3]);
	assign _3401_ = ~(_3400_ | _3397_);
	assign _3402_ = _3401_ & ~_3399_;
	assign _3403_ = _3402_ | _3397_;
	assign _3404_ = \mchip.game2.scroll_inst.pos [1] & \mchip.game2.vga_inst.haddr [1];
	assign _3405_ = \mchip.game2.scroll_inst.pos [0] & \mchip.game2.vga_inst.haddr [0];
	assign _3406_ = ~(\mchip.game2.scroll_inst.pos [1] | \mchip.game2.vga_inst.haddr [1]);
	assign _3407_ = _3406_ | _3404_;
	assign _3408_ = _3405_ & ~_3407_;
	assign _3409_ = _3408_ | _3404_;
	assign _3410_ = ~(\mchip.game2.scroll_inst.pos [2] | \mchip.game2.vga_inst.haddr [2]);
	assign _3411_ = ~(_3410_ | _3398_);
	assign _3412_ = ~(_3411_ & _3401_);
	assign _3413_ = _3409_ & ~_3412_;
	assign _3414_ = _3413_ | _3403_;
	assign _3415_ = ~(\mchip.game2.scroll_inst.pos [4] | \mchip.game2.vga_inst.haddr [4]);
	assign _3416_ = ~(_3415_ | _3388_);
	assign _3417_ = ~(_3416_ & _3390_);
	assign _3418_ = _3417_ | _3394_;
	assign _3419_ = _3414_ & ~_3418_;
	assign _3420_ = _3419_ | _3396_;
	assign _3421_ = \mchip.game2.scroll_inst.pos [8] ^ \mchip.game2.vga_inst.haddr [8];
	assign _3422_ = _3421_ & _3420_;
	assign _3423_ = ~(_3422_ | _3381_);
	assign _3424_ = \mchip.game2.scroll_inst.pos [9] ^ \mchip.game2.vga_inst.haddr [9];
	assign _3425_ = ~_3424_;
	assign _3426_ = _3425_ ^ _3423_;
	assign _3427_ = \mchip.game2.scroll_inst.pos [9] & \mchip.game2.vga_inst.haddr [9];
	assign _3428_ = _3424_ & _3381_;
	assign _3429_ = _3428_ | _3427_;
	assign _3430_ = ~(_3424_ & _3421_);
	assign _3431_ = _3420_ & ~_3430_;
	assign _3432_ = _3431_ | _3429_;
	assign _3433_ = _3432_ | _3426_;
	assign _3434_ = _3421_ ^ _3420_;
	assign _3435_ = _3411_ ^ _3409_;
	assign _3436_ = ~(_3407_ ^ _3405_);
	assign _3437_ = ~_3436_;
	assign _3438_ = _3437_ & ~_3435_;
	assign _3439_ = _3411_ & _3409_;
	assign _3440_ = _3399_ & ~_3439_;
	assign _3441_ = ~(_3440_ ^ _3401_);
	assign _3442_ = _3416_ ^ _3414_;
	assign _3443_ = ~(_3442_ & _3441_);
	assign _3444_ = ~(_3443_ | _3438_);
	assign _3445_ = ~(_3416_ & _3414_);
	assign _3446_ = _3445_ & ~_3388_;
	assign _3447_ = ~(_3446_ ^ _3390_);
	assign _3448_ = _3414_ & ~_3417_;
	assign _3449_ = _3392_ & ~_3448_;
	assign _3450_ = ~(_3449_ ^ _3393_);
	assign _3451_ = ~(_3450_ & _3447_);
	assign _3452_ = _3449_ | ~_3393_;
	assign _3453_ = _3452_ & ~_3383_;
	assign _3454_ = _3453_ ^ _3384_;
	assign _3455_ = _3454_ | _3434_;
	assign _3456_ = _3455_ | _3451_;
	assign _3457_ = _3444_ & ~_3456_;
	assign _3458_ = _3457_ | _3434_;
	assign _3459_ = ~(_3458_ | _3433_);
	assign _3460_ = _3447_ ^ _3444_;
	assign _3461_ = _3441_ & ~_3438_;
	assign _3462_ = _3461_ ^ _3442_;
	assign _3463_ = _3462_ & ~_3460_;
	assign _3464_ = _3444_ & ~_3451_;
	assign _3465_ = _3464_ ^ _3454_;
	assign _3466_ = _3447_ & _3444_;
	assign _3467_ = _3466_ ^ _3450_;
	assign _3468_ = ~(_3467_ | _3465_);
	assign _3469_ = ~(_3468_ & _3463_);
	assign _3470_ = \mchip.game2.scroll_inst.pos [0] ^ \mchip.game2.vga_inst.haddr [0];
	assign _3471_ = ~_3470_;
	assign _3472_ = _3471_ | _3436_;
	assign _3473_ = _3437_ ^ _3435_;
	assign _3474_ = _3438_ & ~_3441_;
	assign _3475_ = ~(_3474_ | _3461_);
	assign _3476_ = _3473_ | ~_3475_;
	assign _3477_ = _3476_ | _3472_;
	assign _3478_ = ~(_3477_ | _3469_);
	assign _3479_ = ~_3426_;
	assign _3480_ = _3479_ & ~_3458_;
	assign _3481_ = _3480_ ^ _3432_;
	assign _3482_ = _3481_ | _3459_;
	assign _3483_ = ~(_3458_ ^ _3479_);
	assign _3484_ = ~_3434_;
	assign _3485_ = _3464_ & ~_3454_;
	assign _3486_ = _3485_ ^ _3484_;
	assign _3487_ = _3486_ | _3483_;
	assign _3488_ = _3487_ | _3482_;
	assign _3489_ = ~(_3488_ | _3459_);
	assign _3490_ = ~(_3489_ & _3478_);
	assign _3491_ = ~(_3490_ | _3459_);
	assign _3492_ = ~_3483_;
	assign _3493_ = _3465_ & ~_3487_;
	assign _3494_ = _3492_ & ~_3493_;
	assign _3495_ = _3468_ & ~_3487_;
	assign _3496_ = _3462_ | _3460_;
	assign _3497_ = _3475_ & _3473_;
	assign _3498_ = _3463_ & ~_3497_;
	assign _3499_ = _3496_ & ~_3498_;
	assign _3500_ = _3495_ & ~_3499_;
	assign _3501_ = _3494_ & ~_3500_;
	assign _3502_ = _3501_ | _3482_;
	assign _3503_ = _3502_ | _3459_;
	assign _3504_ = _3503_ | _3491_;
	assign _3505_ = _3492_ | _3482_;
	assign _3506_ = _3505_ | _3459_;
	assign _3507_ = _3468_ & ~_3496_;
	assign _3508_ = ~(_3471_ & _3436_);
	assign _3509_ = _3475_ | _3473_;
	assign _3510_ = _3509_ | _3508_;
	assign _3511_ = _3510_ | ~_3507_;
	assign _3512_ = _3511_ & ~_3465_;
	assign _3513_ = _3489_ & ~_3512_;
	assign _3514_ = _3506_ & ~_3513_;
	assign _3515_ = ~(_3514_ | _3459_);
	assign _3516_ = _3515_ | _3504_;
	assign _3517_ = _3516_ | io_in[13];
	assign _3518_ = _3517_ | _3380_;
	assign _0014_ = _3518_ | _3230_;
	assign _0005_ = _0006_ & ~_3362_;
	assign _3519_ = ~(\mchip.game2.scroll_inst.tick_time [16] ^ \mchip.game2.scroll_inst.ctr [16]);
	assign _3520_ = \mchip.game2.scroll_inst.tick_time [17] ^ \mchip.game2.scroll_inst.ctr [17];
	assign _3521_ = _3519_ & ~_3520_;
	assign _3522_ = ~(\mchip.game2.scroll_inst.tick_time [8] ^ \mchip.game2.scroll_inst.ctr [8]);
	assign _3523_ = \mchip.game2.scroll_inst.tick_time [9] ^ \mchip.game2.scroll_inst.ctr [9];
	assign _3524_ = _3522_ & ~_3523_;
	assign _3525_ = ~(\mchip.game2.scroll_inst.tick_time [11] ^ \mchip.game2.scroll_inst.ctr [11]);
	assign _3526_ = \mchip.game2.scroll_inst.tick_time [10] ^ \mchip.game2.scroll_inst.ctr [10];
	assign _3527_ = _3526_ | ~_3525_;
	assign _3528_ = _3524_ & ~_3527_;
	assign _3529_ = ~(\mchip.game2.scroll_inst.tick_time [15] ^ \mchip.game2.scroll_inst.ctr [15]);
	assign _3530_ = \mchip.game2.scroll_inst.tick_time [14] ^ \mchip.game2.scroll_inst.ctr [14];
	assign _3531_ = _3529_ & ~_3530_;
	assign _3532_ = \mchip.game2.scroll_inst.tick_time [12] ^ \mchip.game2.scroll_inst.ctr [12];
	assign _3533_ = \mchip.game2.scroll_inst.tick_time [13] ^ \mchip.game2.scroll_inst.ctr [13];
	assign _3534_ = _3533_ | _3532_;
	assign _3535_ = _3534_ | ~_3531_;
	assign _3536_ = _3528_ & ~_3535_;
	assign _3537_ = ~(\mchip.game2.scroll_inst.tick_time [4] ^ \mchip.game2.scroll_inst.ctr [4]);
	assign _3538_ = \mchip.game2.scroll_inst.tick_time [5] ^ \mchip.game2.scroll_inst.ctr [5];
	assign _3539_ = _3537_ & ~_3538_;
	assign _3540_ = ~(\mchip.game2.scroll_inst.tick_time [7] ^ \mchip.game2.scroll_inst.ctr [7]);
	assign _3541_ = \mchip.game2.scroll_inst.tick_time [6] ^ \mchip.game2.scroll_inst.ctr [6];
	assign _3542_ = _3541_ | ~_3540_;
	assign _3543_ = _3539_ & ~_3542_;
	assign _3544_ = ~(\mchip.game2.scroll_inst.ctr [2] ^ \mchip.game2.scroll_inst.tick_time [2]);
	assign _3545_ = \mchip.game2.scroll_inst.ctr [3] ^ \mchip.game2.scroll_inst.tick_time [3];
	assign _3546_ = _3544_ & ~_3545_;
	assign _3547_ = ~(\mchip.game2.scroll_inst.ctr [1] ^ \mchip.game2.scroll_inst.tick_time [1]);
	assign _3548_ = ~(\mchip.game2.scroll_inst.ctr [0] ^ \mchip.game2.scroll_inst.tick_time [0]);
	assign _3549_ = _3548_ & _3547_;
	assign _3550_ = _3549_ & _3546_;
	assign _3551_ = _3550_ & _3543_;
	assign _3552_ = ~(_3551_ & _3536_);
	assign _3553_ = _3552_ | ~_3521_;
	assign _3554_ = \mchip.game2.scroll_inst.ctr [17] | ~\mchip.game2.scroll_inst.tick_time [17];
	assign _3555_ = \mchip.game2.scroll_inst.tick_time [16] & ~\mchip.game2.scroll_inst.ctr [16];
	assign _3556_ = _3555_ & ~_3520_;
	assign _3557_ = _3554_ & ~_3556_;
	assign _3558_ = \mchip.game2.scroll_inst.ctr [15] | ~\mchip.game2.scroll_inst.tick_time [15];
	assign _3559_ = \mchip.game2.scroll_inst.ctr [14] | ~\mchip.game2.scroll_inst.tick_time [14];
	assign _3560_ = _3529_ & ~_3559_;
	assign _3561_ = _3558_ & ~_3560_;
	assign _3562_ = \mchip.game2.scroll_inst.ctr [13] | ~\mchip.game2.scroll_inst.tick_time [13];
	assign _3563_ = \mchip.game2.scroll_inst.tick_time [12] & ~\mchip.game2.scroll_inst.ctr [12];
	assign _3564_ = _3563_ & ~_3533_;
	assign _3565_ = _3562_ & ~_3564_;
	assign _3566_ = _3531_ & ~_3565_;
	assign _3567_ = _3561_ & ~_3566_;
	assign _3568_ = \mchip.game2.scroll_inst.ctr [11] | ~\mchip.game2.scroll_inst.tick_time [11];
	assign _3569_ = \mchip.game2.scroll_inst.ctr [10] | ~\mchip.game2.scroll_inst.tick_time [10];
	assign _3570_ = _3525_ & ~_3569_;
	assign _3571_ = _3568_ & ~_3570_;
	assign _3572_ = \mchip.game2.scroll_inst.ctr [9] | ~\mchip.game2.scroll_inst.tick_time [9];
	assign _3573_ = \mchip.game2.scroll_inst.tick_time [8] & ~\mchip.game2.scroll_inst.ctr [8];
	assign _3574_ = _3573_ & ~_3523_;
	assign _3575_ = _3572_ & ~_3574_;
	assign _3576_ = ~(_3575_ | _3527_);
	assign _3577_ = _3571_ & ~_3576_;
	assign _3578_ = ~(_3577_ | _3535_);
	assign _3579_ = _3567_ & ~_3578_;
	assign _3580_ = \mchip.game2.scroll_inst.ctr [7] | ~\mchip.game2.scroll_inst.tick_time [7];
	assign _3581_ = \mchip.game2.scroll_inst.ctr [6] | ~\mchip.game2.scroll_inst.tick_time [6];
	assign _3582_ = _3540_ & ~_3581_;
	assign _3583_ = _3580_ & ~_3582_;
	assign _3584_ = \mchip.game2.scroll_inst.ctr [5] | ~\mchip.game2.scroll_inst.tick_time [5];
	assign _3585_ = \mchip.game2.scroll_inst.tick_time [4] & ~\mchip.game2.scroll_inst.ctr [4];
	assign _3586_ = _3585_ & ~_3538_;
	assign _3587_ = _3584_ & ~_3586_;
	assign _3588_ = ~(_3587_ | _3542_);
	assign _3589_ = _3583_ & ~_3588_;
	assign _3590_ = \mchip.game2.scroll_inst.ctr [3] | ~\mchip.game2.scroll_inst.tick_time [3];
	assign _3591_ = \mchip.game2.scroll_inst.tick_time [2] & ~\mchip.game2.scroll_inst.ctr [2];
	assign _3592_ = _3591_ & ~_3545_;
	assign _3593_ = _3590_ & ~_3592_;
	assign _3594_ = \mchip.game2.scroll_inst.ctr [1] | ~\mchip.game2.scroll_inst.tick_time [1];
	assign _3595_ = \mchip.game2.scroll_inst.ctr [0] & ~\mchip.game2.scroll_inst.tick_time [0];
	assign _3596_ = _3547_ & ~_3595_;
	assign _3597_ = _3594_ & ~_3596_;
	assign _3598_ = _3546_ & ~_3597_;
	assign _3599_ = _3593_ & ~_3598_;
	assign _3600_ = _3543_ & ~_3599_;
	assign _3601_ = _3589_ & ~_3600_;
	assign _3602_ = _3536_ & ~_3601_;
	assign _3603_ = _3579_ & ~_3602_;
	assign _3604_ = _3521_ & ~_3603_;
	assign _3605_ = _3557_ & ~_3604_;
	assign _3606_ = _3553_ & ~_3605_;
	assign _0002_ = _0163_ & ~_3606_;
	assign _3607_ = ~\mchip.game2.game_over ;
	assign _3608_ = \mchip.game2.start_ctr [22] | ~_0162_;
	assign _3609_ = _3607_ & ~_3608_;
	assign _3610_ = ~\mchip.game2.vga_inst.vaddr [7];
	assign _3611_ = ~(\mchip.game2.jumping_inst.jump_pos [6] & \mchip.game2.vga_inst.vaddr [6]);
	assign _3612_ = _3611_ | _3610_;
	assign _3613_ = \mchip.game2.jumping_inst.jump_pos [6] ^ \mchip.game2.vga_inst.vaddr [6];
	assign _3614_ = _3613_ & ~_3610_;
	assign _3615_ = ~(\mchip.game2.jumping_inst.jump_pos [5] & \mchip.game2.vga_inst.vaddr [5]);
	assign _3616_ = \mchip.game2.jumping_inst.jump_pos [4] & \mchip.game2.vga_inst.vaddr [4];
	assign _3617_ = ~_3616_;
	assign _3618_ = \mchip.game2.jumping_inst.jump_pos [5] | \mchip.game2.vga_inst.vaddr [5];
	assign _3619_ = _3618_ & _3615_;
	assign _0164_ = _3619_ & ~_3617_;
	assign _0165_ = _3615_ & ~_0164_;
	assign _0166_ = _3614_ & ~_0165_;
	assign _0167_ = _3612_ & ~_0166_;
	assign _0168_ = \mchip.game2.jumping_inst.jump_pos [4] ^ \mchip.game2.vga_inst.vaddr [4];
	assign _0169_ = ~_0168_;
	assign _0170_ = _3619_ & ~_0169_;
	assign _0171_ = _0170_ & _3614_;
	assign _0172_ = \mchip.game2.jumping_inst.jump_pos [3] & \mchip.game2.vga_inst.vaddr [3];
	assign _0173_ = \mchip.game2.jumping_inst.jump_pos [2] & \mchip.game2.vga_inst.vaddr [2];
	assign _0174_ = \mchip.game2.jumping_inst.jump_pos [3] ^ \mchip.game2.vga_inst.vaddr [3];
	assign _0175_ = ~(_0174_ & _0173_);
	assign _0176_ = _0175_ & ~_0172_;
	assign _0177_ = ~(\mchip.game2.jumping_inst.jump_pos [2] | \mchip.game2.vga_inst.vaddr [2]);
	assign _0178_ = ~(_0177_ | _0173_);
	assign _0179_ = _0178_ & _0174_;
	assign _0180_ = ~(\mchip.game2.jumping_inst.jump_pos [0] & \mchip.game2.vga_inst.vaddr [0]);
	assign _0181_ = ~(\mchip.game2.jumping_inst.jump_pos [1] ^ \mchip.game2.vga_inst.vaddr [1]);
	assign _0182_ = _0181_ | _0180_;
	assign _0183_ = \mchip.game2.jumping_inst.jump_pos [1] & \mchip.game2.vga_inst.vaddr [1];
	assign _0184_ = _0182_ & ~_0183_;
	assign _0185_ = _0179_ & ~_0184_;
	assign _0186_ = _0176_ & ~_0185_;
	assign _0187_ = _0171_ & ~_0186_;
	assign _0188_ = _0167_ & ~_0187_;
	assign _0189_ = \mchip.game2.vga_inst.vaddr [8] & \mchip.game2.vga_inst.vaddr [9];
	assign _0190_ = _0188_ | ~_0189_;
	assign _0191_ = ~\mchip.game2.vga_inst.vaddr [8];
	assign _0192_ = _0188_ ^ _0191_;
	assign _0193_ = \mchip.game2.vga_inst.vaddr [8] & ~_0188_;
	assign _0194_ = _0193_ ^ \mchip.game2.vga_inst.vaddr [9];
	assign _0195_ = _0194_ | _0192_;
	assign _0196_ = _0190_ & ~_0195_;
	assign _0197_ = _0184_ | ~_0178_;
	assign _0198_ = _0197_ & ~_0173_;
	assign _0199_ = _0198_ ^ _0174_;
	assign _0200_ = _0184_ ^ _0178_;
	assign _0201_ = _0200_ & ~_0199_;
	assign _0202_ = \mchip.game2.jumping_inst.jump_pos [0] ^ \mchip.game2.vga_inst.vaddr [0];
	assign _0203_ = _0181_ ^ _0180_;
	assign _0204_ = _0203_ | _0202_;
	assign _0205_ = _0201_ & ~_0204_;
	assign _0206_ = _0170_ & ~_0186_;
	assign _0207_ = _0165_ & ~_0206_;
	assign _0208_ = _3613_ & ~_0207_;
	assign _0209_ = _3611_ & ~_0208_;
	assign _0210_ = _0209_ ^ \mchip.game2.vga_inst.vaddr [7];
	assign _0211_ = ~(_0207_ ^ _3613_);
	assign _0212_ = _0210_ | ~_0211_;
	assign _0213_ = _0186_ ^ _0169_;
	assign _0214_ = ~(_0186_ | _0169_);
	assign _0215_ = _3617_ & ~_0214_;
	assign _0216_ = ~(_0215_ ^ _3619_);
	assign _0217_ = ~(_0216_ & _0213_);
	assign _0218_ = _0217_ | _0212_;
	assign _0219_ = _0218_ | ~_0205_;
	assign _0220_ = _0196_ & ~_0219_;
	assign _0221_ = ~(_0205_ | _0199_);
	assign _0222_ = _0221_ | _0218_;
	assign _0223_ = _0218_ | ~_0222_;
	assign _0224_ = ~(_0223_ & _0196_);
	assign _0225_ = _0224_ | _0220_;
	assign _0226_ = _0195_ | ~_0210_;
	assign _0227_ = _0211_ | _0210_;
	assign _0228_ = ~(_0227_ | _0195_);
	assign _0229_ = _0216_ | _0213_;
	assign _0230_ = _0213_ & ~_0216_;
	assign _0231_ = ~(_0200_ | _0199_);
	assign _0232_ = _0230_ & ~_0231_;
	assign _0233_ = _0229_ & ~_0232_;
	assign _0234_ = _0228_ & ~_0233_;
	assign _0235_ = _0226_ & ~_0234_;
	assign _0236_ = _0190_ & ~_0235_;
	assign _0237_ = ~(\mchip.game2.vga_inst.haddr [9] | \mchip.game2.vga_inst.haddr [8]);
	assign _0238_ = \mchip.game2.vga_inst.haddr [7] | ~\mchip.game2.vga_inst.haddr [6];
	assign _0239_ = ~(\mchip.game2.vga_inst.haddr [4] | \mchip.game2.vga_inst.haddr [5]);
	assign _0240_ = _0238_ | ~_0239_;
	assign _0241_ = \mchip.game2.vga_inst.haddr [1] & \mchip.game2.vga_inst.haddr [0];
	assign _0242_ = \mchip.game2.vga_inst.haddr [2] | ~\mchip.game2.vga_inst.haddr [3];
	assign _0243_ = _0242_ | ~_0241_;
	assign _0244_ = _0243_ | _0240_;
	assign _0245_ = _0237_ & ~_0244_;
	assign _0246_ = ~(_0237_ & _3182_);
	assign _0247_ = _0237_ & ~_0238_;
	assign _0248_ = ~(\mchip.game2.vga_inst.haddr [2] & \mchip.game2.vga_inst.haddr [3]);
	assign _0249_ = ~(_0248_ & _0239_);
	assign _0250_ = _0247_ & ~_0249_;
	assign _0251_ = _0246_ & ~_0250_;
	assign _0252_ = _0251_ | _0245_;
	assign _0253_ = _0241_ & ~_0248_;
	assign _0254_ = \mchip.game2.vga_inst.haddr [5] | ~\mchip.game2.vga_inst.haddr [4];
	assign _0255_ = _0254_ | ~_3182_;
	assign _0256_ = _0255_ | _0253_;
	assign _0257_ = _0239_ & _3182_;
	assign _0258_ = _0256_ & ~_0257_;
	assign _0259_ = _0237_ & ~_0258_;
	assign _0260_ = _0259_ | _0252_;
	assign _0261_ = _0260_ | _0236_;
	assign _0262_ = _0261_ | _0225_;
	assign _0263_ = _0262_ | _3609_;
	assign _0264_ = io_in[13] | ~_3229_;
	assign _0018_ = _0264_ | _0263_;
	assign _0265_ = ~(\mchip.game2.scroll_inst.pos [8] | \mchip.game2.scroll_inst.pos [9]);
	assign _0266_ = \mchip.game2.scroll_inst.pos [8] & ~\mchip.game2.scroll_inst.pos [9];
	assign _0267_ = \mchip.game2.scroll_inst.pos [6] & \mchip.game2.scroll_inst.pos [7];
	assign _0268_ = \mchip.game2.scroll_inst.pos [4] | \mchip.game2.scroll_inst.pos [5];
	assign _0269_ = _0267_ & ~_0268_;
	assign _0270_ = \mchip.game2.scroll_inst.pos [0] & \mchip.game2.scroll_inst.pos [1];
	assign _0271_ = \mchip.game2.scroll_inst.pos [2] | \mchip.game2.scroll_inst.pos [3];
	assign _0272_ = _0271_ | _0270_;
	assign _0273_ = _0269_ & ~_0272_;
	assign _0274_ = _0267_ & ~_0273_;
	assign _0275_ = _0266_ & ~_0274_;
	assign _0276_ = ~(_0275_ | _0265_);
	assign _0277_ = \mchip.game2.scroll_inst.pos [0] | ~\mchip.game2.scroll_inst.pos [1];
	assign _0278_ = ~(_0277_ | _0271_);
	assign _0279_ = ~(_0278_ & _0269_);
	assign _0280_ = _0266_ & ~_0279_;
	assign _0281_ = ~(_0280_ | _0276_);
	assign _0282_ = ~(\mchip.game2.scroll_inst.pos [0] | \mchip.game2.scroll_inst.pos [1]);
	assign _0283_ = ~(\mchip.game2.scroll_inst.pos [2] & \mchip.game2.scroll_inst.pos [3]);
	assign _0284_ = _0282_ & ~_0283_;
	assign _0285_ = ~(_0284_ & _0269_);
	assign _0286_ = _0266_ & ~_0285_;
	assign _0287_ = ~(_0283_ | _0282_);
	assign _0288_ = _0269_ & ~_0287_;
	assign _0289_ = _0267_ & ~_0288_;
	assign _0290_ = _0289_ | ~_0266_;
	assign _0291_ = _0290_ & ~_0265_;
	assign _0292_ = _0291_ | _0286_;
	assign _0090_ = ~(_0292_ | _0281_);
	assign _0293_ = \mchip.game2.scroll_inst.pos [4] & ~\mchip.game2.scroll_inst.pos [5];
	assign _0294_ = \mchip.game2.scroll_inst.pos [7] | ~\mchip.game2.scroll_inst.pos [6];
	assign _0295_ = _0293_ & ~_0294_;
	assign _0296_ = \mchip.game2.scroll_inst.pos [1] | ~\mchip.game2.scroll_inst.pos [0];
	assign _0297_ = ~(_0296_ | _0283_);
	assign _0298_ = ~(_0297_ & _0295_);
	assign _0299_ = ~(_0265_ & \mchip.game2.scroll_inst.pos [10]);
	assign _0300_ = _0299_ | _0298_;
	assign _0301_ = ~\mchip.game2.scroll_inst.pos [10];
	assign _0302_ = \mchip.game2.scroll_inst.pos [5] & ~_0294_;
	assign _0303_ = _0302_ | \mchip.game2.scroll_inst.pos [7];
	assign _0304_ = _0283_ | _0282_;
	assign _0305_ = _0295_ & ~_0304_;
	assign _0306_ = _0305_ | _0303_;
	assign _0307_ = _0265_ & ~_0306_;
	assign _0308_ = _0307_ | _0301_;
	assign _0309_ = _0308_ | ~_0300_;
	assign _0310_ = _0309_ & ~_0090_;
	assign _0007_ = _3229_ & ~_0310_;
	assign _0311_ = \mchip.game2.rendering_inst.layers [3] | \mchip.game2.rendering_inst.layers [4];
	assign _0312_ = \mchip.game2.rendering_inst.layers [1] | \mchip.game2.rendering_inst.layers [2];
	assign _0313_ = \mchip.game2.score_inst.pixel  | \mchip.game2.rendering_inst.layers [0];
	assign _0314_ = _0313_ | _0312_;
	assign \mchip.game2.dbg_pixel  = _0314_ | _0311_;
	assign _0315_ = io_in[13] | ~\mchip.game2.rendering_inst.cactus_select [2];
	assign _0016_ = _0315_ | _3230_;
	assign _0316_ = \mchip.game2.scroll_inst.pos [6] | \mchip.game2.scroll_inst.pos [7];
	assign _0317_ = _0316_ | _0268_;
	assign _0318_ = \mchip.game2.scroll_inst.pos [3] | ~\mchip.game2.scroll_inst.pos [2];
	assign _0319_ = _0282_ & ~_0318_;
	assign _0320_ = _0317_ | ~_0319_;
	assign _0321_ = _0266_ & ~_0320_;
	assign _0322_ = _0271_ & ~_0319_;
	assign _0323_ = _0322_ | _0317_;
	assign _0324_ = _0266_ & ~_0323_;
	assign _0325_ = ~(_0324_ | _0265_);
	assign _0326_ = ~(_0325_ | _0321_);
	assign _0327_ = ~(\mchip.game2.scroll_inst.pos [4] & \mchip.game2.scroll_inst.pos [5]);
	assign _0328_ = _0267_ & ~_0327_;
	assign _0329_ = \mchip.game2.scroll_inst.pos [2] | ~\mchip.game2.scroll_inst.pos [3];
	assign _0330_ = ~(_0329_ | _0270_);
	assign _0331_ = \mchip.game2.scroll_inst.pos [3] & ~_0330_;
	assign _0332_ = _0328_ & ~_0331_;
	assign _0333_ = _0328_ & ~_0332_;
	assign _0334_ = _0265_ & ~_0333_;
	assign _0335_ = _0329_ | _0277_;
	assign _0336_ = _0335_ | ~_0328_;
	assign _0337_ = _0265_ & ~_0336_;
	assign _0338_ = _0334_ & ~_0337_;
	assign _0089_ = _0326_ & ~_0338_;
	assign _0339_ = ~\mchip.game2.jumping_inst.in_air ;
	assign _0011_ = _0163_ & ~_0339_;
	assign _0340_ = io_in[0] & \mchip.game2.game_over ;
	assign _0341_ = ~(\mchip.game2.no_jump_ctr [19] | \mchip.game2.no_jump_ctr [18]);
	assign _0342_ = \mchip.game2.no_jump_ctr [17] | ~\mchip.game2.no_jump_ctr [16];
	assign _0343_ = _0341_ & ~_0342_;
	assign _0344_ = \mchip.game2.no_jump_ctr [15] & ~\mchip.game2.no_jump_ctr [14];
	assign _0345_ = \mchip.game2.no_jump_ctr [12] | \mchip.game2.no_jump_ctr [13];
	assign _0346_ = _0344_ & ~_0345_;
	assign _0347_ = \mchip.game2.no_jump_ctr [10] | \mchip.game2.no_jump_ctr [11];
	assign _0348_ = \mchip.game2.no_jump_ctr [11] | ~\mchip.game2.no_jump_ctr [10];
	assign _0349_ = ~(_0348_ | \mchip.game2.no_jump_ctr [9]);
	assign _0350_ = _0347_ & ~_0349_;
	assign _0351_ = _0346_ & ~_0350_;
	assign _0352_ = \mchip.game2.no_jump_ctr [15] & ~_0351_;
	assign _0353_ = \mchip.game2.no_jump_ctr [8] | ~\mchip.game2.no_jump_ctr [9];
	assign _0354_ = _0353_ | _0348_;
	assign _0355_ = _0346_ & ~_0354_;
	assign _0356_ = \mchip.game2.no_jump_ctr [7] & ~\mchip.game2.no_jump_ctr [6];
	assign _0357_ = _0356_ & ~\mchip.game2.no_jump_ctr [5];
	assign _0358_ = \mchip.game2.no_jump_ctr [7] & ~_0357_;
	assign _0359_ = \mchip.game2.no_jump_ctr [4] | ~\mchip.game2.no_jump_ctr [5];
	assign _0360_ = _0356_ & ~_0359_;
	assign _0361_ = \mchip.game2.no_jump_ctr [0] | \mchip.game2.no_jump_ctr [1];
	assign _0362_ = \mchip.game2.no_jump_ctr [2] | \mchip.game2.no_jump_ctr [3];
	assign _0363_ = _0362_ | _0361_;
	assign _0364_ = _0360_ & ~_0363_;
	assign _0365_ = _0358_ & ~_0364_;
	assign _0366_ = _0355_ & ~_0365_;
	assign _0367_ = _0352_ & ~_0366_;
	assign _0368_ = _0343_ & ~_0367_;
	assign _0369_ = \mchip.game2.no_jump_ctr [16] | \mchip.game2.no_jump_ctr [17];
	assign _0370_ = _0341_ & ~_0369_;
	assign _0371_ = _0370_ | _0368_;
	assign _0372_ = _0340_ & ~_0371_;
	assign _0373_ = \mchip.game2.rendering_inst.layers [3] | \mchip.game2.rendering_inst.layers [1];
	assign _0374_ = _0373_ | \mchip.game2.rendering_inst.layers [4];
	assign _0375_ = _0374_ & \mchip.game2.rendering_inst.layers [0];
	assign _0376_ = _0375_ & ~io_in[2];
	assign _0001_ = _0376_ | _0372_;
	assign _0377_ = \mchip.game2.scroll_inst.pos [8] & \mchip.game2.scroll_inst.pos [9];
	assign _0378_ = ~_0377_;
	assign _0379_ = ~(_0318_ | _0296_);
	assign _0380_ = \mchip.game2.scroll_inst.pos [6] | ~\mchip.game2.scroll_inst.pos [7];
	assign _0381_ = _0293_ & ~_0380_;
	assign _0382_ = ~(_0381_ & _0379_);
	assign _0383_ = _0382_ | _0378_;
	assign _0384_ = \mchip.game2.scroll_inst.pos [5] & ~_0380_;
	assign _0385_ = ~(_0384_ | _0267_);
	assign _0386_ = _0318_ | _0282_;
	assign _0387_ = _0386_ & ~\mchip.game2.scroll_inst.pos [3];
	assign _0388_ = _0381_ & ~_0387_;
	assign _0389_ = _0385_ & ~_0388_;
	assign _0390_ = _0389_ | _0378_;
	assign _0391_ = _0390_ | ~_0383_;
	assign _0392_ = _0391_ & ~_0089_;
	assign _0008_ = _3229_ & ~_0392_;
	assign _0019_ = io_in[0] | io_in[13];
	assign _0393_ = _0331_ | _0317_;
	assign _0394_ = _0265_ & ~_0393_;
	assign _0395_ = _0335_ | _0317_;
	assign _0396_ = _0265_ & ~_0395_;
	assign _0088_ = _0394_ & ~_0396_;
	assign _0397_ = _3198_ & _3190_;
	assign _0398_ = ~(_0397_ & _3194_);
	assign _0399_ = _3188_ & ~_0398_;
	assign _0400_ = _3206_ & _3193_;
	assign _0401_ = _0400_ | ~_3205_;
	assign _0402_ = _0401_ & ~_3210_;
	assign _0403_ = _0402_ | _0399_;
	assign _0404_ = \mchip.game2.vga_inst.vaddr [3] | ~\mchip.game2.vga_inst.vaddr [2];
	assign _0405_ = _3219_ & ~_0404_;
	assign _0406_ = _3218_ & ~_0405_;
	assign _0407_ = _3194_ & ~_0406_;
	assign _0408_ = _3194_ & ~_0407_;
	assign _0409_ = _3188_ & ~_0408_;
	assign _0410_ = _0409_ | _0403_;
	assign _0017_ = _0410_ | _0264_;
	assign _0411_ = \mchip.game2.dinosprite_inst.ctr [21] & ~\mchip.game2.dinosprite_inst.ctr [20];
	assign _0412_ = \mchip.game2.dinosprite_inst.ctr [22] | \mchip.game2.dinosprite_inst.ctr [23];
	assign _0413_ = _0411_ & ~_0412_;
	assign _0414_ = \mchip.game2.dinosprite_inst.ctr [16] & ~\mchip.game2.dinosprite_inst.ctr [17];
	assign _0415_ = \mchip.game2.dinosprite_inst.ctr [18] & \mchip.game2.dinosprite_inst.ctr [19];
	assign _0416_ = ~(_0415_ & _0414_);
	assign _0417_ = _0416_ | ~_0413_;
	assign _0418_ = _0417_ | \mchip.game2.dinosprite_inst.ctr [24];
	assign _0419_ = \mchip.game2.dinosprite_inst.ctr [9] & ~\mchip.game2.dinosprite_inst.ctr [8];
	assign _0420_ = \mchip.game2.dinosprite_inst.ctr [11] | ~\mchip.game2.dinosprite_inst.ctr [10];
	assign _0421_ = _0419_ & ~_0420_;
	assign _0422_ = \mchip.game2.dinosprite_inst.ctr [12] | \mchip.game2.dinosprite_inst.ctr [13];
	assign _0423_ = ~(\mchip.game2.dinosprite_inst.ctr [14] & \mchip.game2.dinosprite_inst.ctr [15]);
	assign _0424_ = _0423_ | _0422_;
	assign _0425_ = _0421_ & ~_0424_;
	assign _0426_ = ~(\mchip.game2.dinosprite_inst.ctr [0] | \mchip.game2.dinosprite_inst.ctr [1]);
	assign _0427_ = \mchip.game2.dinosprite_inst.ctr [2] | \mchip.game2.dinosprite_inst.ctr [3];
	assign _0428_ = _0426_ & ~_0427_;
	assign _0429_ = ~(\mchip.game2.dinosprite_inst.ctr [4] | \mchip.game2.dinosprite_inst.ctr [5]);
	assign _0430_ = \mchip.game2.dinosprite_inst.ctr [6] & \mchip.game2.dinosprite_inst.ctr [7];
	assign _0431_ = ~(_0430_ & _0429_);
	assign _0432_ = _0428_ & ~_0431_;
	assign _0433_ = ~(_0432_ & _0425_);
	assign _0434_ = _0433_ | _0418_;
	assign _0435_ = _0412_ | \mchip.game2.dinosprite_inst.ctr [21];
	assign _0436_ = ~(\mchip.game2.dinosprite_inst.ctr [17] | \mchip.game2.dinosprite_inst.ctr [16]);
	assign _0437_ = _0415_ & ~_0436_;
	assign _0438_ = _0413_ & ~_0437_;
	assign _0439_ = _0435_ & ~_0438_;
	assign _0440_ = \mchip.game2.dinosprite_inst.ctr [10] | \mchip.game2.dinosprite_inst.ctr [11];
	assign _0441_ = ~\mchip.game2.dinosprite_inst.ctr [9];
	assign _0442_ = _0441_ & ~_0420_;
	assign _0443_ = _0440_ & ~_0442_;
	assign _0444_ = ~(_0443_ | _0424_);
	assign _0445_ = ~(_0444_ | _0423_);
	assign _0446_ = _0430_ & ~_0432_;
	assign _0447_ = _0425_ & ~_0446_;
	assign _0448_ = _0445_ & ~_0447_;
	assign _0449_ = ~(_0448_ | _0417_);
	assign _0450_ = _0439_ & ~_0449_;
	assign _0451_ = _0450_ | \mchip.game2.dinosprite_inst.ctr [24];
	assign _0452_ = _0434_ & ~_0451_;
	assign _0012_ = _0163_ & ~_0452_;
	assign _0020_ = _0372_ | io_in[13];
	assign _0453_ = \mchip.game2.scroll_inst.pos [9] & ~\mchip.game2.scroll_inst.pos [8];
	assign _0454_ = _0270_ & ~_0329_;
	assign _0455_ = _0454_ & _0381_;
	assign _0456_ = ~(_0455_ & _0453_);
	assign _0457_ = _0283_ & ~_0454_;
	assign _0458_ = _0381_ & ~_0457_;
	assign _0459_ = _0385_ & ~_0458_;
	assign _0460_ = _0453_ & ~_0459_;
	assign _0461_ = _0378_ & ~_0460_;
	assign _0462_ = _0461_ | ~_0456_;
	assign _0463_ = _0462_ & ~_0088_;
	assign _0009_ = _3229_ & ~_0463_;
	assign _0464_ = \mchip.game2.jumping_inst.ctr [22] | \mchip.game2.jumping_inst.ctr [23];
	assign _0465_ = \mchip.game2.jumping_inst.ctr [20] | \mchip.game2.jumping_inst.ctr [21];
	assign _0466_ = _0465_ | _0464_;
	assign _0467_ = \mchip.game2.jumping_inst.ctr [18] | \mchip.game2.jumping_inst.ctr [19];
	assign _0468_ = ~(\mchip.game2.jumping_inst.ctr [16] & \mchip.game2.jumping_inst.ctr [17]);
	assign _0469_ = _0468_ | _0467_;
	assign _0470_ = _0469_ | _0466_;
	assign _0471_ = ~(\mchip.game2.jumping_inst.ctr [14] & \mchip.game2.jumping_inst.ctr [15]);
	assign _0472_ = \mchip.game2.jumping_inst.ctr [13] | ~\mchip.game2.jumping_inst.ctr [12];
	assign _0473_ = _0472_ | _0471_;
	assign _0474_ = \mchip.game2.jumping_inst.ctr [10] | \mchip.game2.jumping_inst.ctr [11];
	assign _0475_ = \mchip.game2.jumping_inst.ctr [8] | \mchip.game2.jumping_inst.ctr [9];
	assign _0476_ = _0475_ | _0474_;
	assign _0477_ = _0476_ | _0473_;
	assign _0478_ = \mchip.game2.jumping_inst.ctr [6] | ~\mchip.game2.jumping_inst.ctr [7];
	assign _0479_ = \mchip.game2.jumping_inst.ctr [5] | ~\mchip.game2.jumping_inst.ctr [4];
	assign _0480_ = _0479_ | _0478_;
	assign _0481_ = \mchip.game2.jumping_inst.ctr [2] | \mchip.game2.jumping_inst.ctr [3];
	assign _0482_ = \mchip.game2.jumping_inst.ctr [0] | \mchip.game2.jumping_inst.ctr [1];
	assign _0483_ = _0482_ | _0481_;
	assign _0484_ = _0483_ | _0480_;
	assign _0485_ = _0484_ | _0477_;
	assign _0486_ = _0485_ | _0470_;
	assign _0487_ = _0486_ | _0339_;
	assign _0010_ = _0163_ & ~_0487_;
	assign _0024_ = \mchip.game2.rendering_inst.cactus_select [2] & ~\mchip.game2.cactus_select_last [2];
	assign _0025_ = \mchip.game2.rendering_inst.cactus_select [1] & ~\mchip.game2.cactus_select_last [1];
	assign _0026_ = \mchip.game2.rendering_inst.cactus_select [0] & ~\mchip.game2.cactus_select_last [0];
	assign _0488_ = \mchip.game2.vga_inst.vaddr [5] | ~\mchip.game2.vga_inst.vaddr [4];
	assign _0489_ = \mchip.game2.vga_inst.vaddr [6] | \mchip.game2.vga_inst.vaddr [7];
	assign _0490_ = _0489_ | _0488_;
	assign _0491_ = _0490_ | _0406_;
	assign _0492_ = _3207_ & ~_0489_;
	assign _0493_ = _0491_ & ~_0492_;
	assign _0494_ = _0493_ | _3197_;
	assign _0495_ = \mchip.game2.vga_inst.vaddr [6] & ~\mchip.game2.vga_inst.vaddr [7];
	assign _0496_ = ~(_0495_ & _3207_);
	assign _0497_ = \mchip.game2.vga_inst.vaddr [0] & ~\mchip.game2.vga_inst.vaddr [1];
	assign _0498_ = ~(_0497_ & _3190_);
	assign _0499_ = _0498_ | _0496_;
	assign _0500_ = _3188_ & ~_0499_;
	assign _0501_ = ~\mchip.game2.vga_inst.vaddr [6];
	assign _0502_ = ~(\mchip.game2.vga_inst.vaddr [7] | \mchip.game2.vga_inst.vaddr [8]);
	assign _0503_ = ~(_0502_ & _0501_);
	assign _0504_ = \mchip.game2.vga_inst.vaddr [5] | ~\mchip.game2.vga_inst.vaddr [6];
	assign _0505_ = _0502_ & ~_0504_;
	assign _0506_ = \mchip.game2.vga_inst.vaddr [3] | \mchip.game2.vga_inst.vaddr [4];
	assign _0507_ = \mchip.game2.vga_inst.vaddr [3] & ~\mchip.game2.vga_inst.vaddr [4];
	assign _0508_ = \mchip.game2.vga_inst.vaddr [1] | \mchip.game2.vga_inst.vaddr [2];
	assign _0509_ = _0507_ & ~_0508_;
	assign _0510_ = _0506_ & ~_0509_;
	assign _0511_ = _0505_ & ~_0510_;
	assign _0512_ = _0503_ & ~_0511_;
	assign _0513_ = _0512_ | \mchip.game2.vga_inst.vaddr [9];
	assign _0514_ = _0513_ | _0500_;
	assign _0092_ = _0494_ & ~_0514_;
	assign _0515_ = ~(_0497_ | _3189_);
	assign _0516_ = ~\mchip.game2.vga_inst.vaddr [2];
	assign _0517_ = _3198_ ^ _0516_;
	assign _0518_ = _0517_ | ~_0515_;
	assign _0519_ = ~\mchip.game2.vga_inst.vaddr [3];
	assign _0520_ = _0516_ & ~_3198_;
	assign _0521_ = _0520_ ^ _0519_;
	assign _0522_ = _3198_ | \mchip.game2.vga_inst.vaddr [2];
	assign _0523_ = (_0521_ ? _0518_ : _0522_);
	assign _0524_ = ~(_0397_ | _3206_);
	assign _0525_ = _0524_ ^ \mchip.game2.vga_inst.vaddr [4];
	assign _0526_ = _0523_ | ~_0525_;
	assign _0527_ = _0524_ & ~\mchip.game2.vga_inst.vaddr [4];
	assign _0528_ = _0527_ ^ \mchip.game2.vga_inst.vaddr [5];
	assign _0529_ = _0528_ | _0526_;
	assign _0530_ = _0517_ & ~_0515_;
	assign _0531_ = _0530_ & _0521_;
	assign _0532_ = ~_0531_;
	assign _0533_ = (_0528_ ? _0532_ : _0526_);
	assign _0534_ = (_3470_ ? _0529_ : _0533_);
	assign _0535_ = ~_3189_;
	assign _0536_ = _0517_ & ~_0535_;
	assign _0537_ = ~(_0536_ | _0521_);
	assign _0538_ = _0530_ | _0521_;
	assign _0539_ = (_0525_ ? _0537_ : _0538_);
	assign _0540_ = _0528_ | ~_0539_;
	assign _0541_ = _3198_ & ~\mchip.game2.vga_inst.vaddr [2];
	assign _0542_ = _0521_ & ~_0541_;
	assign _0543_ = (_0525_ ? _0542_ : _0537_);
	assign _0544_ = _0543_ | _0528_;
	assign _0545_ = (_3470_ ? _0540_ : _0544_);
	assign _0546_ = (_3436_ ? _0534_ : _0545_);
	assign _0547_ = _0546_ | _3467_;
	assign _0548_ = _0547_ | _3473_;
	assign _0549_ = _0521_ | _0518_;
	assign _0550_ = _0549_ | _0525_;
	assign _0551_ = ~(_0550_ | _0528_);
	assign _0552_ = _0551_ | _3467_;
	assign _0553_ = ~_0525_;
	assign _0554_ = ~_0521_;
	assign _0555_ = _0535_ & ~_0517_;
	assign _0556_ = _0555_ | _0536_;
	assign _0557_ = _0556_ | _0554_;
	assign _0558_ = _0557_ | _0553_;
	assign _0559_ = _0558_ | _0528_;
	assign _0560_ = _0559_ | _3467_;
	assign _0561_ = (_3470_ ? _0552_ : _0560_);
	assign _0562_ = _0521_ | ~_0541_;
	assign _0563_ = ~(_0562_ | _0525_);
	assign _0564_ = _0563_ & ~_0528_;
	assign _0565_ = _0564_ | _3467_;
	assign _0566_ = (_3470_ ? _0552_ : _0565_);
	assign _0567_ = (_3436_ ? _0561_ : _0566_);
	assign _0568_ = ~_0528_;
	assign _0569_ = _0521_ & ~_0555_;
	assign _0570_ = ~_0569_;
	assign _0571_ = ~_0517_;
	assign _0572_ = _0521_ & ~_0571_;
	assign _0573_ = (_0525_ ? _0570_ : _0572_);
	assign _0574_ = ~(_0573_ & _0568_);
	assign _0575_ = _0574_ | _3467_;
	assign _0576_ = _0575_ | ~_3470_;
	assign _0577_ = _0521_ & ~_0522_;
	assign _0578_ = (_0525_ ? _0577_ : _0570_);
	assign _0579_ = _0578_ | _0528_;
	assign _0580_ = _0579_ | _3467_;
	assign _0581_ = (_3470_ ? _0560_ : _0580_);
	assign _0582_ = (_3436_ ? _0576_ : _0581_);
	assign _0583_ = (_3473_ ? _0567_ : _0582_);
	assign _0584_ = (_3475_ ? _0548_ : _0583_);
	assign _0585_ = ~(_0584_ | _3462_);
	assign _3631_ = _0585_ & ~_3460_;
	assign _0586_ = _3219_ ^ _0516_;
	assign _0587_ = _3189_ & ~_0586_;
	assign _0588_ = _0587_ & ~_3470_;
	assign _0589_ = (_0586_ ? \mchip.game2.vga_inst.vaddr [0] : _3189_);
	assign _0590_ = ~\mchip.game2.vga_inst.vaddr [0];
	assign _0591_ = (_0586_ ? _0590_ : _3189_);
	assign _0592_ = (_3470_ ? _0589_ : _0591_);
	assign _0593_ = (_3436_ ? _0588_ : _0592_);
	assign _0594_ = (_3470_ ? _0591_ : _0587_);
	assign _0595_ = (_3436_ ? _0594_ : _0587_);
	assign _0596_ = (_3435_ ? _0593_ : _0595_);
	assign _0597_ = _0590_ & ~_0586_;
	assign _0598_ = (_3470_ ? _0587_ : _0597_);
	assign _0599_ = (_3436_ ? _0598_ : _0587_);
	assign _0600_ = (_3470_ ? _0587_ : _0589_);
	assign _0601_ = (_3436_ ? _0587_ : _0600_);
	assign _0602_ = (_3435_ ? _0599_ : _0601_);
	assign _0603_ = (_3441_ ? _0596_ : _0602_);
	assign _0604_ = (_3436_ ? _0587_ : _0598_);
	assign _0605_ = (_3435_ ? _0587_ : _0604_);
	assign _0606_ = (_3470_ ? _0589_ : _0587_);
	assign _0607_ = (_3436_ ? _0606_ : _0594_);
	assign _0608_ = (_3435_ ? _0587_ : _0607_);
	assign _0609_ = (_3441_ ? _0605_ : _0608_);
	assign _0610_ = (_3442_ ? _0603_ : _0609_);
	assign _0611_ = (_3470_ ? _0597_ : _0587_);
	assign _0612_ = (_3436_ ? _0611_ : _0597_);
	assign _0613_ = (_3435_ ? _0612_ : _0587_);
	assign _0614_ = (_3441_ ? _0605_ : _0613_);
	assign _0615_ = (_3470_ ? _0587_ : _0591_);
	assign _0616_ = (_3436_ ? _0615_ : _0611_);
	assign _0617_ = (_3435_ ? _0616_ : _0595_);
	assign _0618_ = (_3436_ ? _0591_ : _0611_);
	assign _0619_ = (_3435_ ? _0587_ : _0618_);
	assign _0620_ = (_3441_ ? _0617_ : _0619_);
	assign _0621_ = (_3442_ ? _0614_ : _0620_);
	assign _0622_ = (_3447_ ? _0610_ : _0621_);
	assign _0623_ = (_3436_ ? _0587_ : _0606_);
	assign _0624_ = (_3435_ ? _0623_ : _0601_);
	assign _0625_ = (_3441_ ? _0624_ : _0587_);
	assign _0626_ = _0497_ & ~_0586_;
	assign _0627_ = (_3470_ ? _0587_ : _0626_);
	assign _0628_ = (_0586_ ? \mchip.game2.vga_inst.vaddr [0] : _0497_);
	assign _0629_ = _3219_ | _3198_;
	assign _0630_ = ~(_0629_ | _0586_);
	assign _0631_ = (_3470_ ? _0628_ : _0630_);
	assign _0632_ = (_3436_ ? _0627_ : _0631_);
	assign _0633_ = \mchip.game2.vga_inst.vaddr [1] & \mchip.game2.vga_inst.vaddr [2];
	assign _0634_ = (_3470_ ? _0597_ : _0633_);
	assign _0635_ = (_3436_ ? _0587_ : _0634_);
	assign _0636_ = (_3435_ ? _0632_ : _0635_);
	assign _0637_ = _3198_ & ~_0586_;
	assign _0638_ = (_3470_ ? _0637_ : _0633_);
	assign _0639_ = (_3436_ ? _0637_ : _0638_);
	assign _0640_ = (_3436_ ? _0598_ : _0600_);
	assign _0641_ = (_3435_ ? _0639_ : _0640_);
	assign _0642_ = (_3441_ ? _0636_ : _0641_);
	assign _0643_ = (_3442_ ? _0625_ : _0642_);
	assign _0644_ = (_3470_ ? _0597_ : _0589_);
	assign _0645_ = (_3436_ ? _0644_ : _0587_);
	assign _0646_ = (_3435_ ? _0645_ : _0587_);
	assign _0647_ = (_3441_ ? _0587_ : _0646_);
	assign _0648_ = _0623_ & _3435_;
	assign _0649_ = _0623_ & ~_3435_;
	assign _0650_ = _0649_ | _0648_;
	assign _0651_ = (_3435_ ? _0623_ : _0604_);
	assign _0652_ = (_3441_ ? _0650_ : _0651_);
	assign _0653_ = (_3442_ ? _0647_ : _0652_);
	assign _0654_ = (_3447_ ? _0643_ : _0653_);
	assign _0655_ = (_3450_ ? _0622_ : _0654_);
	assign _0656_ = (_3436_ ? _0587_ : _0592_);
	assign _0657_ = (_3435_ ? _0656_ : _0595_);
	assign _0658_ = (_3441_ ? _0657_ : _0602_);
	assign _0659_ = (_3442_ ? _0658_ : _0609_);
	assign _0660_ = (_3447_ ? _0659_ : _0621_);
	assign _0661_ = (_3450_ ? _0660_ : _0654_);
	assign _3630_ = (_3454_ ? _0661_ : _0655_);
	assign _0028_ = ~\mchip.game2.dinosprite_inst.sprite ;
	assign _0662_ = ~\mchip.game2.vga_inst.haddr [3];
	assign _0663_ = \mchip.game2.vga_inst.haddr [2] & \mchip.game2.vga_inst.haddr [1];
	assign _0664_ = _0663_ & ~_0662_;
	assign _0665_ = _0664_ ^ \mchip.game2.vga_inst.haddr [4];
	assign _0666_ = ~\mchip.game2.vga_inst.haddr [1];
	assign _0667_ = _0172_ & _0168_;
	assign _0668_ = _0172_ ^ _0168_;
	assign _0669_ = ~_0668_;
	assign _0670_ = _0177_ | ~_0174_;
	assign _0671_ = ~(\mchip.game2.jumping_inst.jump_pos [2] ^ \mchip.game2.vga_inst.vaddr [2]);
	assign _0672_ = _0671_ & _0183_;
	assign _0673_ = ~(_0177_ ^ _0174_);
	assign _0674_ = _0673_ & _0672_;
	assign _0675_ = _0670_ & ~_0674_;
	assign _0676_ = ~(\mchip.game2.jumping_inst.jump_pos [0] | \mchip.game2.vga_inst.vaddr [0]);
	assign _0677_ = ~(_0676_ | _0181_);
	assign _0678_ = _0671_ ^ _0183_;
	assign _0679_ = ~(_0678_ & _0673_);
	assign _0680_ = _0677_ & ~_0679_;
	assign _0681_ = _0675_ & ~_0680_;
	assign _0682_ = _0681_ | _0669_;
	assign _0683_ = _0682_ & ~_0667_;
	assign _0684_ = ~(\mchip.game2.jumping_inst.jump_pos [5] ^ \mchip.game2.vga_inst.vaddr [5]);
	assign _0685_ = _0684_ ^ _3616_;
	assign _0686_ = _0685_ ^ _0683_;
	assign _0687_ = _0678_ ^ _0677_;
	assign _0688_ = _0676_ ^ _0181_;
	assign _0689_ = ~_0688_;
	assign _0690_ = _0689_ & ~_0687_;
	assign _0691_ = ~(_0678_ & _0677_);
	assign _0692_ = _0691_ & ~_0672_;
	assign _0693_ = ~(_0692_ ^ _0673_);
	assign _0694_ = _0693_ & ~_0690_;
	assign _0695_ = _0681_ ^ _0669_;
	assign _0696_ = _0694_ | ~_0695_;
	assign _0697_ = _0696_ | _0686_;
	assign _0698_ = _0684_ & _3616_;
	assign _0699_ = _0685_ & _0667_;
	assign _0700_ = ~(_0699_ | _0698_);
	assign _0701_ = ~(_0685_ & _0668_);
	assign _0702_ = ~(_0701_ | _0681_);
	assign _0703_ = _0700_ & ~_0702_;
	assign _0704_ = ~(\mchip.game2.jumping_inst.jump_pos [6] ^ \mchip.game2.vga_inst.vaddr [6]);
	assign _0705_ = _0704_ ^ _3618_;
	assign _0706_ = ~(_0705_ ^ _0703_);
	assign _0707_ = ~_0706_;
	assign _0708_ = _0697_ | ~_0707_;
	assign _0709_ = _0708_ | _0028_;
	assign _0710_ = _0028_ & ~_0708_;
	assign _0711_ = _0709_ & ~_0710_;
	assign _0712_ = ~_0687_;
	assign _0713_ = _0693_ & ~_0712_;
	assign _0714_ = _0713_ | ~_0695_;
	assign _0715_ = _0714_ | _0686_;
	assign _0716_ = _0715_ | _0706_;
	assign _0717_ = (\mchip.game2.game_over  ? _0716_ : _0711_);
	assign _0718_ = ~(\mchip.game2.vga_inst.haddr [3] & \mchip.game2.vga_inst.haddr [4]);
	assign _0719_ = _0663_ & ~_0718_;
	assign _0720_ = _3174_ & ~_0719_;
	assign _0721_ = _0720_ ^ \mchip.game2.vga_inst.haddr [7];
	assign _0722_ = _0721_ | _0717_;
	assign _0723_ = _0722_ | _0666_;
	assign _0724_ = ~(\mchip.game2.vga_inst.haddr [2] | \mchip.game2.vga_inst.haddr [1]);
	assign _0725_ = ~(_0724_ | _0663_);
	assign _0726_ = _0725_ | _0723_;
	assign _0727_ = _0663_ ^ \mchip.game2.vga_inst.haddr [3];
	assign _0728_ = _0687_ & ~_0689_;
	assign _0729_ = ~(_0728_ & _0693_);
	assign _0730_ = (_0695_ ? _0694_ : _0729_);
	assign _0731_ = _0730_ | _0686_;
	assign _0732_ = _0731_ | ~_0707_;
	assign _0733_ = _0732_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0734_ = \mchip.game2.dinosprite_inst.sprite  & ~_0732_;
	assign _0735_ = _0733_ & ~_0734_;
	assign _0736_ = (_0695_ ? _0713_ : _0729_);
	assign _0737_ = _0736_ | _0686_;
	assign _0738_ = _0737_ | ~_0707_;
	assign _0739_ = (\mchip.game2.game_over  ? _0738_ : _0735_);
	assign _0740_ = _0739_ | _0721_;
	assign _0741_ = ~(_0676_ ^ _0181_);
	assign _0742_ = _0693_ & ~_0741_;
	assign _0743_ = (_0695_ ? _0742_ : _0729_);
	assign _0744_ = _0743_ | _0686_;
	assign _0745_ = _0744_ | ~_0707_;
	assign _0746_ = _0745_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0747_ = \mchip.game2.dinosprite_inst.sprite  & ~_0745_;
	assign _0748_ = _0746_ & ~_0747_;
	assign _0749_ = _0729_ & ~_0695_;
	assign _0750_ = _0729_ | ~_0695_;
	assign _0751_ = _0749_ | ~_0750_;
	assign _0752_ = _0751_ | _0686_;
	assign _0753_ = _0752_ | ~_0707_;
	assign _0754_ = (\mchip.game2.game_over  ? _0753_ : _0748_);
	assign _0755_ = _0754_ | _0721_;
	assign _0756_ = (\mchip.game2.vga_inst.haddr [1] ? _0755_ : _0740_);
	assign _0757_ = _0689_ ^ _0687_;
	assign _0758_ = _0757_ | _0693_;
	assign _0759_ = _0758_ | _0695_;
	assign _0760_ = (_0706_ ? _0759_ : _0744_);
	assign _0761_ = _0760_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0762_ = \mchip.game2.dinosprite_inst.sprite  & ~_0760_;
	assign _0763_ = _0761_ & ~_0762_;
	assign _0764_ = (_0706_ ? _0759_ : _0752_);
	assign _0765_ = (\mchip.game2.game_over  ? _0764_ : _0763_);
	assign _0766_ = _0765_ | _0721_;
	assign _0767_ = (\mchip.game2.vga_inst.haddr [1] ? _0766_ : _0755_);
	assign _0768_ = (_0725_ ? _0756_ : _0767_);
	assign _0769_ = (_0727_ ? _0726_ : _0768_);
	assign _0770_ = ~(_0769_ | _0665_);
	assign _0771_ = ~\mchip.game2.vga_inst.haddr [5];
	assign _0772_ = _0719_ ^ _0771_;
	assign _0773_ = _0689_ | _0687_;
	assign _0774_ = ~(_0773_ | _0693_);
	assign _0775_ = _0695_ | ~_0774_;
	assign _0776_ = (_0706_ ? _0775_ : _0752_);
	assign _0777_ = _0776_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0778_ = \mchip.game2.dinosprite_inst.sprite  & ~_0776_;
	assign _0779_ = _0777_ & ~_0778_;
	assign _0780_ = (\mchip.game2.game_over  ? _0776_ : _0779_);
	assign _0781_ = _0695_ | _0694_;
	assign _0782_ = _0749_ | _0686_;
	assign _0783_ = (_0706_ ? _0781_ : _0782_);
	assign _0784_ = _0783_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0785_ = \mchip.game2.dinosprite_inst.sprite  & ~_0783_;
	assign _0786_ = _0784_ & ~_0785_;
	assign _0787_ = (\mchip.game2.game_over  ? _0783_ : _0786_);
	assign _0788_ = (\mchip.game2.vga_inst.haddr [1] ? _0787_ : _0780_);
	assign _0789_ = ~_0749_;
	assign _0790_ = (_0695_ ? _0774_ : _0729_);
	assign _0791_ = _0790_ | _0686_;
	assign _0792_ = (_0706_ ? _0789_ : _0791_);
	assign _0793_ = _0792_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0794_ = \mchip.game2.dinosprite_inst.sprite  & ~_0792_;
	assign _0795_ = _0793_ & ~_0794_;
	assign _0796_ = (\mchip.game2.game_over  ? _0792_ : _0795_);
	assign _0797_ = ~_0690_;
	assign _0798_ = _0693_ & ~_0797_;
	assign _0799_ = _0695_ & ~_0798_;
	assign _0800_ = (_0706_ ? _0799_ : _0782_);
	assign _0801_ = _0695_ & ~_0774_;
	assign _0802_ = (_0706_ ? _0801_ : _0782_);
	assign _0803_ = (\mchip.game2.dinosprite_inst.sprite  ? _0800_ : _0802_);
	assign _0804_ = (\mchip.game2.game_over  ? _0800_ : _0803_);
	assign _0805_ = (\mchip.game2.vga_inst.haddr [1] ? _0804_ : _0796_);
	assign _0806_ = (_0725_ ? _0788_ : _0805_);
	assign _0807_ = _0695_ & _0694_;
	assign _0808_ = ~_0695_;
	assign _0809_ = _0808_ | _0686_;
	assign _0810_ = (_0706_ ? _0807_ : _0809_);
	assign _0811_ = _0712_ & ~_0693_;
	assign _0812_ = _0695_ & ~_0811_;
	assign _0813_ = (_0706_ ? _0812_ : _0809_);
	assign _0814_ = (\mchip.game2.dinosprite_inst.sprite  ? _0810_ : _0813_);
	assign _0815_ = (\mchip.game2.game_over  ? _0810_ : _0814_);
	assign _0816_ = _0750_ | _0686_;
	assign _0817_ = (_0706_ ? _0812_ : _0816_);
	assign _0818_ = _0690_ & ~_0693_;
	assign _0819_ = _0695_ & ~_0818_;
	assign _0820_ = (_0706_ ? _0819_ : _0816_);
	assign _0821_ = (\mchip.game2.dinosprite_inst.sprite  ? _0817_ : _0820_);
	assign _0822_ = (\mchip.game2.game_over  ? _0817_ : _0821_);
	assign _0823_ = (\mchip.game2.vga_inst.haddr [1] ? _0822_ : _0815_);
	assign _0824_ = _0819_ | ~_0706_;
	assign _0825_ = _0824_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0826_ = \mchip.game2.dinosprite_inst.sprite  & ~_0824_;
	assign _0827_ = _0825_ & ~_0826_;
	assign _0828_ = (\mchip.game2.game_over  ? _0824_ : _0827_);
	assign _0829_ = _0812_ | ~_0706_;
	assign _0830_ = _0689_ & ~_0693_;
	assign _0831_ = _0830_ | ~_0695_;
	assign _0832_ = ~(_0831_ & _0706_);
	assign _0833_ = (\mchip.game2.dinosprite_inst.sprite  ? _0832_ : _0829_);
	assign _0834_ = (\mchip.game2.game_over  ? _0829_ : _0833_);
	assign _0835_ = (\mchip.game2.vga_inst.haddr [1] ? _0834_ : _0828_);
	assign _0836_ = (_0725_ ? _0823_ : _0835_);
	assign _0837_ = (_0727_ ? _0806_ : _0836_);
	assign _0838_ = ~(_0837_ | _0721_);
	assign _0839_ = (_0695_ ? _0694_ : _0818_);
	assign _0840_ = ~(_0728_ | _0693_);
	assign _0841_ = ~_0840_;
	assign _0842_ = (_0695_ ? _0841_ : _0818_);
	assign _0843_ = (\mchip.game2.dinosprite_inst.sprite  ? _0842_ : _0839_);
	assign _0844_ = (_0693_ ? _0797_ : _0728_);
	assign _0845_ = (_0695_ ? _0844_ : _0818_);
	assign _0846_ = (\mchip.game2.game_over  ? _0845_ : _0843_);
	assign _0847_ = _0846_ | _0707_;
	assign _0848_ = (_0695_ ? _0694_ : _0811_);
	assign _0849_ = _0848_ | ~_0706_;
	assign _0850_ = ~(_0811_ ^ _0695_);
	assign _0851_ = ~(_0850_ & _0706_);
	assign _0852_ = (\mchip.game2.dinosprite_inst.sprite  ? _0851_ : _0849_);
	assign _0853_ = (\mchip.game2.game_over  ? _0849_ : _0852_);
	assign _0854_ = (\mchip.game2.vga_inst.haddr [1] ? _0853_ : _0847_);
	assign _0855_ = (_0695_ ? _0818_ : _0841_);
	assign _0856_ = ~(_0855_ & _0706_);
	assign _0857_ = _0856_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0858_ = \mchip.game2.dinosprite_inst.sprite  & ~_0856_;
	assign _0859_ = _0857_ & ~_0858_;
	assign _0860_ = (\mchip.game2.game_over  ? _0856_ : _0859_);
	assign _0861_ = ~(_0840_ | _0695_);
	assign _0862_ = ~(_0861_ & _0706_);
	assign _0863_ = _0862_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0864_ = \mchip.game2.dinosprite_inst.sprite  & ~_0862_;
	assign _0865_ = _0863_ & ~_0864_;
	assign _0866_ = (\mchip.game2.game_over  ? _0862_ : _0865_);
	assign _0867_ = (\mchip.game2.vga_inst.haddr [1] ? _0866_ : _0860_);
	assign _0868_ = (_0725_ ? _0854_ : _0867_);
	assign _0869_ = ~(_0868_ | _0721_);
	assign _0870_ = (_0693_ ? _0728_ : _0712_);
	assign _0871_ = ~(_0870_ | _0695_);
	assign _0872_ = ~(_0871_ & _0706_);
	assign _0873_ = _0872_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0874_ = \mchip.game2.dinosprite_inst.sprite  & ~_0872_;
	assign _0875_ = _0873_ & ~_0874_;
	assign _0876_ = (\mchip.game2.game_over  ? _0872_ : _0875_);
	assign _0877_ = (_0693_ ? _0687_ : _0690_);
	assign _0878_ = ~(_0877_ | _0695_);
	assign _0879_ = ~(_0878_ & _0706_);
	assign _0880_ = _0879_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0881_ = \mchip.game2.dinosprite_inst.sprite  & ~_0879_;
	assign _0882_ = _0880_ & ~_0881_;
	assign _0883_ = (\mchip.game2.game_over  ? _0879_ : _0882_);
	assign _0884_ = (\mchip.game2.vga_inst.haddr [1] ? _0883_ : _0876_);
	assign _0885_ = ~(_0884_ | _0721_);
	assign _0886_ = (_0706_ ? _0781_ : _0816_);
	assign _0887_ = _0886_ | \mchip.game2.dinosprite_inst.sprite ;
	assign _0888_ = \mchip.game2.dinosprite_inst.sprite  & ~_0886_;
	assign _0889_ = _0887_ & ~_0888_;
	assign _0890_ = (\mchip.game2.game_over  ? _0886_ : _0889_);
	assign _0891_ = _0890_ | _0721_;
	assign _0892_ = _0666_ & ~_0891_;
	assign _0893_ = (_0725_ ? _0885_ : _0892_);
	assign _0894_ = (_0727_ ? _0869_ : _0893_);
	assign _0895_ = (_0665_ ? _0838_ : _0894_);
	assign _0896_ = (_0772_ ? _0770_ : _0895_);
	assign _0897_ = _0771_ & ~_0719_;
	assign _0898_ = _0897_ ^ \mchip.game2.vga_inst.haddr [6];
	assign _3629_ = _0896_ & ~_0898_;
	assign _0064_ = _0486_ & ~\mchip.game2.jumping_inst.ctr [0];
	assign _0899_ = \mchip.game2.jumping_inst.ctr [0] & \mchip.game2.jumping_inst.ctr [1];
	assign _0900_ = _0899_ | ~_0482_;
	assign _0075_ = _0486_ & ~_0900_;
	assign _0901_ = ~(_0899_ ^ \mchip.game2.jumping_inst.ctr [2]);
	assign _0080_ = _0486_ & ~_0901_;
	assign _0902_ = ~(_0899_ & \mchip.game2.jumping_inst.ctr [2]);
	assign _0903_ = _0902_ ^ \mchip.game2.jumping_inst.ctr [3];
	assign _0081_ = _0486_ & ~_0903_;
	assign _0904_ = ~(\mchip.game2.jumping_inst.ctr [2] & \mchip.game2.jumping_inst.ctr [3]);
	assign _0905_ = _0899_ & ~_0904_;
	assign _0906_ = ~(_0905_ ^ \mchip.game2.jumping_inst.ctr [4]);
	assign _0082_ = _0486_ & ~_0906_;
	assign _0907_ = ~(_0905_ & \mchip.game2.jumping_inst.ctr [4]);
	assign _0908_ = _0907_ ^ \mchip.game2.jumping_inst.ctr [5];
	assign _0083_ = _0486_ & ~_0908_;
	assign _0909_ = ~(\mchip.game2.jumping_inst.ctr [4] & \mchip.game2.jumping_inst.ctr [5]);
	assign _0910_ = _0905_ & ~_0909_;
	assign _0911_ = ~(_0910_ ^ \mchip.game2.jumping_inst.ctr [6]);
	assign _0084_ = _0486_ & ~_0911_;
	assign _0912_ = ~(_0910_ & \mchip.game2.jumping_inst.ctr [6]);
	assign _0913_ = _0912_ ^ \mchip.game2.jumping_inst.ctr [7];
	assign _0085_ = _0486_ & ~_0913_;
	assign _0914_ = ~(\mchip.game2.jumping_inst.ctr [7] & \mchip.game2.jumping_inst.ctr [6]);
	assign _0915_ = _0914_ | _0909_;
	assign _0916_ = _0905_ & ~_0915_;
	assign _0917_ = ~(_0916_ ^ \mchip.game2.jumping_inst.ctr [8]);
	assign _0086_ = _0486_ & ~_0917_;
	assign _0918_ = ~(_0916_ & \mchip.game2.jumping_inst.ctr [8]);
	assign _0919_ = _0918_ ^ \mchip.game2.jumping_inst.ctr [9];
	assign _0087_ = _0486_ & ~_0919_;
	assign _0920_ = ~(\mchip.game2.jumping_inst.ctr [8] & \mchip.game2.jumping_inst.ctr [9]);
	assign _0921_ = _0916_ & ~_0920_;
	assign _0922_ = ~(_0921_ ^ \mchip.game2.jumping_inst.ctr [10]);
	assign _0065_ = _0486_ & ~_0922_;
	assign _0923_ = ~(_0921_ & \mchip.game2.jumping_inst.ctr [10]);
	assign _0924_ = _0923_ ^ \mchip.game2.jumping_inst.ctr [11];
	assign _0066_ = _0486_ & ~_0924_;
	assign _0925_ = ~(\mchip.game2.jumping_inst.ctr [10] & \mchip.game2.jumping_inst.ctr [11]);
	assign _0926_ = _0925_ | _0920_;
	assign _0927_ = _0916_ & ~_0926_;
	assign _0928_ = ~(_0927_ ^ \mchip.game2.jumping_inst.ctr [12]);
	assign _0067_ = _0486_ & ~_0928_;
	assign _0929_ = ~(_0927_ & \mchip.game2.jumping_inst.ctr [12]);
	assign _0930_ = _0929_ ^ \mchip.game2.jumping_inst.ctr [13];
	assign _0068_ = _0486_ & ~_0930_;
	assign _0931_ = ~(\mchip.game2.jumping_inst.ctr [12] & \mchip.game2.jumping_inst.ctr [13]);
	assign _0932_ = _0927_ & ~_0931_;
	assign _0933_ = ~(_0932_ ^ \mchip.game2.jumping_inst.ctr [14]);
	assign _0069_ = _0486_ & ~_0933_;
	assign _0934_ = ~(_0932_ & \mchip.game2.jumping_inst.ctr [14]);
	assign _0935_ = _0934_ ^ \mchip.game2.jumping_inst.ctr [15];
	assign _0070_ = _0486_ & ~_0935_;
	assign _0936_ = _0931_ | _0471_;
	assign _0937_ = ~(_0936_ | _0926_);
	assign _0938_ = ~(_0937_ & _0916_);
	assign _0939_ = _0938_ ^ \mchip.game2.jumping_inst.ctr [16];
	assign _0071_ = _0486_ & ~_0939_;
	assign _0940_ = _0938_ | ~\mchip.game2.jumping_inst.ctr [16];
	assign _0941_ = _0940_ ^ \mchip.game2.jumping_inst.ctr [17];
	assign _0072_ = _0486_ & ~_0941_;
	assign _0942_ = ~(_0938_ | _0468_);
	assign _0943_ = ~(_0942_ ^ \mchip.game2.jumping_inst.ctr [18]);
	assign _0073_ = _0486_ & ~_0943_;
	assign _0944_ = ~(_0942_ & \mchip.game2.jumping_inst.ctr [18]);
	assign _0945_ = _0944_ ^ \mchip.game2.jumping_inst.ctr [19];
	assign _0074_ = _0486_ & ~_0945_;
	assign _0946_ = ~(\mchip.game2.jumping_inst.ctr [18] & \mchip.game2.jumping_inst.ctr [19]);
	assign _0947_ = _0946_ | _0468_;
	assign _0948_ = ~(_0947_ | _0938_);
	assign _0949_ = ~(_0948_ ^ \mchip.game2.jumping_inst.ctr [20]);
	assign _0076_ = _0486_ & ~_0949_;
	assign _0950_ = ~(_0948_ & \mchip.game2.jumping_inst.ctr [20]);
	assign _0951_ = _0950_ ^ \mchip.game2.jumping_inst.ctr [21];
	assign _0077_ = _0486_ & ~_0951_;
	assign _0952_ = ~(\mchip.game2.jumping_inst.ctr [20] & \mchip.game2.jumping_inst.ctr [21]);
	assign _0953_ = _0948_ & ~_0952_;
	assign _0954_ = ~(_0953_ ^ \mchip.game2.jumping_inst.ctr [22]);
	assign _0078_ = _0486_ & ~_0954_;
	assign _0955_ = ~(_0953_ & \mchip.game2.jumping_inst.ctr [22]);
	assign _0956_ = _0955_ ^ \mchip.game2.jumping_inst.ctr [23];
	assign _0079_ = _0486_ & ~_0956_;
	assign _0957_ = \mchip.game2.jumping_inst.frame [1] & \mchip.game2.jumping_inst.frame [0];
	assign _0958_ = ~(\mchip.game2.jumping_inst.frame [3] & \mchip.game2.jumping_inst.frame [2]);
	assign _0959_ = _0957_ & ~_0958_;
	assign _0960_ = _0959_ ^ \mchip.game2.jumping_inst.frame [4];
	assign _0961_ = ~\mchip.game2.jumping_inst.frame [5];
	assign _0962_ = ~\mchip.game2.jumping_inst.frame [4];
	assign _0963_ = _0959_ & ~_0962_;
	assign _0964_ = _0963_ ^ _0961_;
	assign _0965_ = _0964_ | ~_0960_;
	assign _0966_ = ~(\mchip.game2.jumping_inst.frame [4] & \mchip.game2.jumping_inst.frame [5]);
	assign _0967_ = _0959_ & ~_0966_;
	assign _0968_ = _0967_ ^ \mchip.game2.jumping_inst.frame [6];
	assign _0969_ = _0967_ & \mchip.game2.jumping_inst.frame [6];
	assign _0970_ = _0969_ ^ \mchip.game2.jumping_inst.frame [7];
	assign _0971_ = _0970_ | _0968_;
	assign _0972_ = _0971_ | ~_0965_;
	assign _0973_ = \mchip.game2.jumping_inst.frame [1] & ~\mchip.game2.jumping_inst.frame [0];
	assign _0974_ = ~_0973_;
	assign _0975_ = _0957_ ^ \mchip.game2.jumping_inst.frame [2];
	assign _0976_ = ~\mchip.game2.jumping_inst.frame [2];
	assign _0977_ = _0957_ & ~_0976_;
	assign _0978_ = _0977_ ^ \mchip.game2.jumping_inst.frame [3];
	assign _0979_ = _0978_ | _0975_;
	assign _0980_ = _0974_ & ~_0979_;
	assign _0981_ = _0971_ | _0965_;
	assign _0982_ = _0980_ & ~_0981_;
	assign _0983_ = _0972_ & ~_0982_;
	assign _0984_ = ~(\mchip.game2.jumping_inst.frame [7] & \mchip.game2.jumping_inst.frame [6]);
	assign _0985_ = _0984_ | _0966_;
	assign _0986_ = _0959_ & ~_0985_;
	assign _0987_ = _0986_ | \mchip.game2.jumping_inst.frame [8];
	assign _0988_ = _0987_ | _0983_;
	assign _0989_ = \mchip.game2.jumping_inst.frame [0] & ~\mchip.game2.jumping_inst.frame [1];
	assign _0990_ = ~_0989_;
	assign _0991_ = _0990_ | _0979_;
	assign _0992_ = _0991_ | _0981_;
	assign _0993_ = ~(_0992_ | _0987_);
	assign _0994_ = _0993_ | _0988_;
	assign _0055_ = ~(_0994_ | \mchip.game2.jumping_inst.frame [0]);
	assign _0995_ = _0989_ | _0973_;
	assign _0056_ = _0995_ & ~_0994_;
	assign _0057_ = _0975_ & ~_0994_;
	assign _0058_ = _0978_ & ~_0994_;
	assign _0059_ = _0960_ & ~_0994_;
	assign _0060_ = ~(_0994_ | _0964_);
	assign _0061_ = _0968_ & ~_0994_;
	assign _0062_ = _0970_ & ~_0994_;
	assign _0996_ = ~(_0986_ ^ \mchip.game2.jumping_inst.frame [8]);
	assign _0063_ = ~(_0996_ | _0994_);
	assign _0997_ = _0486_ | ~_0994_;
	assign _0054_ = (\mchip.game2.jumping_inst.in_air  ? _0997_ : io_in[0]);
	assign _0029_ = _0452_ & ~\mchip.game2.dinosprite_inst.ctr [0];
	assign _0998_ = \mchip.game2.dinosprite_inst.ctr [0] & \mchip.game2.dinosprite_inst.ctr [1];
	assign _0999_ = _0998_ | _0426_;
	assign _0040_ = _0452_ & ~_0999_;
	assign _1000_ = ~(_0998_ ^ \mchip.game2.dinosprite_inst.ctr [2]);
	assign _0046_ = _0452_ & ~_1000_;
	assign _1001_ = ~(_0998_ & \mchip.game2.dinosprite_inst.ctr [2]);
	assign _1002_ = _1001_ ^ \mchip.game2.dinosprite_inst.ctr [3];
	assign _0047_ = _0452_ & ~_1002_;
	assign _1003_ = ~(\mchip.game2.dinosprite_inst.ctr [2] & \mchip.game2.dinosprite_inst.ctr [3]);
	assign _1004_ = _0998_ & ~_1003_;
	assign _1005_ = ~(_1004_ ^ \mchip.game2.dinosprite_inst.ctr [4]);
	assign _0048_ = _0452_ & ~_1005_;
	assign _1006_ = ~(_1004_ & \mchip.game2.dinosprite_inst.ctr [4]);
	assign _1007_ = _1006_ ^ \mchip.game2.dinosprite_inst.ctr [5];
	assign _0049_ = _0452_ & ~_1007_;
	assign _1008_ = ~(\mchip.game2.dinosprite_inst.ctr [4] & \mchip.game2.dinosprite_inst.ctr [5]);
	assign _1009_ = _1004_ & ~_1008_;
	assign _1010_ = ~(_1009_ ^ \mchip.game2.dinosprite_inst.ctr [6]);
	assign _0050_ = _0452_ & ~_1010_;
	assign _1011_ = ~(_1009_ & \mchip.game2.dinosprite_inst.ctr [6]);
	assign _1012_ = _1011_ ^ \mchip.game2.dinosprite_inst.ctr [7];
	assign _0051_ = _0452_ & ~_1012_;
	assign _1013_ = ~\mchip.game2.dinosprite_inst.ctr [8];
	assign _1014_ = _1008_ | ~_0430_;
	assign _1015_ = _1004_ & ~_1014_;
	assign _1016_ = _1015_ ^ _1013_;
	assign _0052_ = _0452_ & ~_1016_;
	assign _1017_ = _1015_ & ~_1013_;
	assign _1018_ = _1017_ ^ _0441_;
	assign _0053_ = _0452_ & ~_1018_;
	assign _1019_ = ~(\mchip.game2.dinosprite_inst.ctr [9] & \mchip.game2.dinosprite_inst.ctr [8]);
	assign _1020_ = _1015_ & ~_1019_;
	assign _1021_ = ~(_1020_ ^ \mchip.game2.dinosprite_inst.ctr [10]);
	assign _0030_ = _0452_ & ~_1021_;
	assign _1022_ = ~(_1020_ & \mchip.game2.dinosprite_inst.ctr [10]);
	assign _1023_ = _1022_ ^ \mchip.game2.dinosprite_inst.ctr [11];
	assign _0031_ = _0452_ & ~_1023_;
	assign _1024_ = ~(\mchip.game2.dinosprite_inst.ctr [10] & \mchip.game2.dinosprite_inst.ctr [11]);
	assign _1025_ = _1024_ | _1019_;
	assign _1026_ = _1015_ & ~_1025_;
	assign _1027_ = ~(_1026_ ^ \mchip.game2.dinosprite_inst.ctr [12]);
	assign _0032_ = _0452_ & ~_1027_;
	assign _1028_ = ~(_1026_ & \mchip.game2.dinosprite_inst.ctr [12]);
	assign _1029_ = _1028_ ^ \mchip.game2.dinosprite_inst.ctr [13];
	assign _0033_ = _0452_ & ~_1029_;
	assign _1030_ = ~(\mchip.game2.dinosprite_inst.ctr [12] & \mchip.game2.dinosprite_inst.ctr [13]);
	assign _1031_ = _1026_ & ~_1030_;
	assign _1032_ = ~(_1031_ ^ \mchip.game2.dinosprite_inst.ctr [14]);
	assign _0034_ = _0452_ & ~_1032_;
	assign _1033_ = ~(_1031_ & \mchip.game2.dinosprite_inst.ctr [14]);
	assign _1034_ = _1033_ ^ \mchip.game2.dinosprite_inst.ctr [15];
	assign _0035_ = _0452_ & ~_1034_;
	assign _1035_ = _1030_ | _0423_;
	assign _1036_ = _1035_ | _1025_;
	assign _1037_ = _1015_ & ~_1036_;
	assign _1038_ = ~(_1037_ ^ \mchip.game2.dinosprite_inst.ctr [16]);
	assign _0036_ = _0452_ & ~_1038_;
	assign _1039_ = ~(_1037_ & \mchip.game2.dinosprite_inst.ctr [16]);
	assign _1040_ = _1039_ ^ \mchip.game2.dinosprite_inst.ctr [17];
	assign _0037_ = _0452_ & ~_1040_;
	assign _1041_ = ~(\mchip.game2.dinosprite_inst.ctr [17] & \mchip.game2.dinosprite_inst.ctr [16]);
	assign _1042_ = _1037_ & ~_1041_;
	assign _1043_ = ~(_1042_ ^ \mchip.game2.dinosprite_inst.ctr [18]);
	assign _0038_ = _0452_ & ~_1043_;
	assign _1044_ = ~(_1042_ & \mchip.game2.dinosprite_inst.ctr [18]);
	assign _1045_ = _1044_ ^ \mchip.game2.dinosprite_inst.ctr [19];
	assign _0039_ = _0452_ & ~_1045_;
	assign _1046_ = _1041_ | ~_0415_;
	assign _1047_ = _1037_ & ~_1046_;
	assign _1048_ = ~(_1047_ ^ \mchip.game2.dinosprite_inst.ctr [20]);
	assign _0041_ = _0452_ & ~_1048_;
	assign _1049_ = ~(_1047_ & \mchip.game2.dinosprite_inst.ctr [20]);
	assign _1050_ = _1049_ ^ \mchip.game2.dinosprite_inst.ctr [21];
	assign _0042_ = _0452_ & ~_1050_;
	assign _1051_ = ~(\mchip.game2.dinosprite_inst.ctr [21] & \mchip.game2.dinosprite_inst.ctr [20]);
	assign _1052_ = _1047_ & ~_1051_;
	assign _1053_ = ~(_1052_ ^ \mchip.game2.dinosprite_inst.ctr [22]);
	assign _0043_ = _0452_ & ~_1053_;
	assign _1054_ = ~(_1052_ & \mchip.game2.dinosprite_inst.ctr [22]);
	assign _1055_ = _1054_ ^ \mchip.game2.dinosprite_inst.ctr [23];
	assign _0044_ = _0452_ & ~_1055_;
	assign _1056_ = ~(\mchip.game2.dinosprite_inst.ctr [22] & \mchip.game2.dinosprite_inst.ctr [23]);
	assign _1057_ = _1056_ | _1051_;
	assign _1058_ = _1057_ | _1046_;
	assign _1059_ = _1058_ | ~_1037_;
	assign _1060_ = _1059_ ^ \mchip.game2.dinosprite_inst.ctr [24];
	assign _0045_ = _0452_ & ~_1060_;
	assign _0132_ = _3606_ & ~\mchip.game2.scroll_inst.ctr [0];
	assign _1061_ = ~(\mchip.game2.scroll_inst.ctr [1] ^ \mchip.game2.scroll_inst.ctr [0]);
	assign _0141_ = _3606_ & ~_1061_;
	assign _1062_ = \mchip.game2.scroll_inst.ctr [1] & \mchip.game2.scroll_inst.ctr [0];
	assign _1063_ = ~(_1062_ ^ \mchip.game2.scroll_inst.ctr [2]);
	assign _0142_ = _3606_ & ~_1063_;
	assign _1064_ = ~(_1062_ & \mchip.game2.scroll_inst.ctr [2]);
	assign _1065_ = _1064_ ^ \mchip.game2.scroll_inst.ctr [3];
	assign _0143_ = _3606_ & ~_1065_;
	assign _1066_ = ~(\mchip.game2.scroll_inst.ctr [2] & \mchip.game2.scroll_inst.ctr [3]);
	assign _1067_ = _1062_ & ~_1066_;
	assign _1068_ = ~(_1067_ ^ \mchip.game2.scroll_inst.ctr [4]);
	assign _0144_ = _3606_ & ~_1068_;
	assign _1069_ = ~(_1067_ & \mchip.game2.scroll_inst.ctr [4]);
	assign _1070_ = _1069_ ^ \mchip.game2.scroll_inst.ctr [5];
	assign _0145_ = _3606_ & ~_1070_;
	assign _1071_ = ~(\mchip.game2.scroll_inst.ctr [4] & \mchip.game2.scroll_inst.ctr [5]);
	assign _1072_ = _1067_ & ~_1071_;
	assign _1073_ = ~(_1072_ ^ \mchip.game2.scroll_inst.ctr [6]);
	assign _0146_ = _3606_ & ~_1073_;
	assign _1074_ = ~(_1072_ & \mchip.game2.scroll_inst.ctr [6]);
	assign _1075_ = _1074_ ^ \mchip.game2.scroll_inst.ctr [7];
	assign _0147_ = _3606_ & ~_1075_;
	assign _1076_ = ~(\mchip.game2.scroll_inst.ctr [6] & \mchip.game2.scroll_inst.ctr [7]);
	assign _1077_ = _1076_ | _1071_;
	assign _1078_ = _1067_ & ~_1077_;
	assign _1079_ = ~(_1078_ ^ \mchip.game2.scroll_inst.ctr [8]);
	assign _0148_ = _3606_ & ~_1079_;
	assign _1080_ = ~(_1078_ & \mchip.game2.scroll_inst.ctr [8]);
	assign _1081_ = _1080_ ^ \mchip.game2.scroll_inst.ctr [9];
	assign _0149_ = _3606_ & ~_1081_;
	assign _1082_ = ~(\mchip.game2.scroll_inst.ctr [8] & \mchip.game2.scroll_inst.ctr [9]);
	assign _1083_ = _1078_ & ~_1082_;
	assign _1084_ = ~(_1083_ ^ \mchip.game2.scroll_inst.ctr [10]);
	assign _0133_ = _3606_ & ~_1084_;
	assign _1085_ = ~(_1083_ & \mchip.game2.scroll_inst.ctr [10]);
	assign _1086_ = _1085_ ^ \mchip.game2.scroll_inst.ctr [11];
	assign _0134_ = _3606_ & ~_1086_;
	assign _1087_ = ~(\mchip.game2.scroll_inst.ctr [10] & \mchip.game2.scroll_inst.ctr [11]);
	assign _1088_ = _1087_ | _1082_;
	assign _1089_ = _1078_ & ~_1088_;
	assign _1090_ = ~(_1089_ ^ \mchip.game2.scroll_inst.ctr [12]);
	assign _0135_ = _3606_ & ~_1090_;
	assign _1091_ = ~(_1089_ & \mchip.game2.scroll_inst.ctr [12]);
	assign _1092_ = _1091_ ^ \mchip.game2.scroll_inst.ctr [13];
	assign _0136_ = _3606_ & ~_1092_;
	assign _1093_ = ~(\mchip.game2.scroll_inst.ctr [12] & \mchip.game2.scroll_inst.ctr [13]);
	assign _1094_ = _1089_ & ~_1093_;
	assign _1095_ = ~(_1094_ ^ \mchip.game2.scroll_inst.ctr [14]);
	assign _0137_ = _3606_ & ~_1095_;
	assign _1096_ = ~(_1094_ & \mchip.game2.scroll_inst.ctr [14]);
	assign _1097_ = _1096_ ^ \mchip.game2.scroll_inst.ctr [15];
	assign _0138_ = _3606_ & ~_1097_;
	assign _1098_ = ~(\mchip.game2.scroll_inst.ctr [14] & \mchip.game2.scroll_inst.ctr [15]);
	assign _1099_ = _1098_ | _1093_;
	assign _1100_ = _1099_ | _1088_;
	assign _1101_ = _1078_ & ~_1100_;
	assign _1102_ = ~(_1101_ ^ \mchip.game2.scroll_inst.ctr [16]);
	assign _0139_ = _3606_ & ~_1102_;
	assign _1103_ = ~(_1101_ & \mchip.game2.scroll_inst.ctr [16]);
	assign _1104_ = _1103_ ^ \mchip.game2.scroll_inst.ctr [17];
	assign _0140_ = _3606_ & ~_1104_;
	assign _1105_ = ~(_0497_ & _3206_);
	assign _1106_ = _0492_ & ~_1105_;
	assign _1107_ = \mchip.game2.vga_inst.vaddr [9] & ~\mchip.game2.vga_inst.vaddr [8];
	assign _1108_ = ~(_1107_ & _1106_);
	assign _1109_ = _3219_ | ~_3206_;
	assign _1110_ = _0492_ & ~_1109_;
	assign _1111_ = _0492_ & ~_1110_;
	assign _1112_ = _1107_ & ~_1111_;
	assign _1113_ = _1112_ | _0189_;
	assign _1114_ = _1108_ & ~_1113_;
	assign _0152_ = _1114_ & ~\mchip.game2.vga_inst.vaddr [0];
	assign _0153_ = _1114_ & ~_0515_;
	assign _1115_ = _3198_ & ~_0516_;
	assign _1116_ = _1115_ | _0520_;
	assign _0154_ = _1114_ & ~_1116_;
	assign _1117_ = _1115_ ^ _0519_;
	assign _0155_ = _1114_ & ~_1117_;
	assign _1118_ = ~(_3206_ & _3198_);
	assign _1119_ = _1118_ ^ \mchip.game2.vga_inst.vaddr [4];
	assign _0156_ = _1114_ & ~_1119_;
	assign _1120_ = \mchip.game2.vga_inst.vaddr [4] & ~_1118_;
	assign _1121_ = _1120_ ^ _3214_;
	assign _0157_ = _1114_ & ~_1121_;
	assign _1122_ = _3193_ & ~_1118_;
	assign _1123_ = _1122_ ^ _0501_;
	assign _0158_ = _1114_ & ~_1123_;
	assign _1124_ = _1122_ & ~_0501_;
	assign _1125_ = _1124_ ^ _3610_;
	assign _0159_ = _1114_ & ~_1125_;
	assign _1126_ = _3194_ & ~_1118_;
	assign _1127_ = _1126_ ^ _0191_;
	assign _0160_ = _1114_ & ~_1127_;
	assign _1128_ = ~(_1126_ & \mchip.game2.vga_inst.vaddr [8]);
	assign _1129_ = _1128_ ^ \mchip.game2.vga_inst.vaddr [9];
	assign _0161_ = _1114_ & ~_1129_;
	assign _0110_ = _3331_ & ~\mchip.game2.score_inst.ctr [0];
	assign _1130_ = \mchip.game2.score_inst.ctr [0] & \mchip.game2.score_inst.ctr [1];
	assign _1131_ = _1130_ | ~_3299_;
	assign _0121_ = _3331_ & ~_1131_;
	assign _1132_ = ~(_1130_ ^ \mchip.game2.score_inst.ctr [2]);
	assign _0124_ = _3331_ & ~_1132_;
	assign _1133_ = ~(_1130_ & \mchip.game2.score_inst.ctr [2]);
	assign _1134_ = _1133_ ^ \mchip.game2.score_inst.ctr [3];
	assign _0125_ = _3331_ & ~_1134_;
	assign _1135_ = _3300_ | ~_1130_;
	assign _1136_ = _1135_ ^ \mchip.game2.score_inst.ctr [4];
	assign _0126_ = _3331_ & ~_1136_;
	assign _1137_ = _1135_ | ~\mchip.game2.score_inst.ctr [4];
	assign _1138_ = _1137_ ^ \mchip.game2.score_inst.ctr [5];
	assign _0127_ = _3331_ & ~_1138_;
	assign _1139_ = ~(_1135_ | _3296_);
	assign _1140_ = ~(_1139_ ^ \mchip.game2.score_inst.ctr [6]);
	assign _0128_ = _3331_ & ~_1140_;
	assign _1141_ = ~(_1139_ & \mchip.game2.score_inst.ctr [6]);
	assign _1142_ = _1141_ ^ \mchip.game2.score_inst.ctr [7];
	assign _0129_ = _3331_ & ~_1142_;
	assign _1143_ = ~\mchip.game2.score_inst.ctr [8];
	assign _1144_ = ~(_1135_ | _3298_);
	assign _1145_ = _1144_ ^ _1143_;
	assign _0130_ = _3331_ & ~_1145_;
	assign _1146_ = _1144_ & ~_1143_;
	assign _1147_ = _1146_ ^ _3319_;
	assign _0131_ = _3331_ & ~_1147_;
	assign _1148_ = ~(\mchip.game2.score_inst.ctr [8] & \mchip.game2.score_inst.ctr [9]);
	assign _1149_ = _1144_ & ~_1148_;
	assign _1150_ = ~(_1149_ ^ \mchip.game2.score_inst.ctr [10]);
	assign _0111_ = _3331_ & ~_1150_;
	assign _1151_ = ~(_1149_ & \mchip.game2.score_inst.ctr [10]);
	assign _1152_ = _1151_ ^ \mchip.game2.score_inst.ctr [11];
	assign _0112_ = _3331_ & ~_1152_;
	assign _1153_ = _1148_ | _3312_;
	assign _1154_ = _1153_ | ~_1144_;
	assign _1155_ = _1154_ ^ \mchip.game2.score_inst.ctr [12];
	assign _0113_ = _3331_ & ~_1155_;
	assign _1156_ = _1154_ | ~\mchip.game2.score_inst.ctr [12];
	assign _1157_ = _1156_ ^ \mchip.game2.score_inst.ctr [13];
	assign _0114_ = _3331_ & ~_1157_;
	assign _1158_ = ~\mchip.game2.score_inst.ctr [14];
	assign _1159_ = ~(_1154_ | _3311_);
	assign _1160_ = _1159_ ^ _1158_;
	assign _0115_ = _3331_ & ~_1160_;
	assign _1161_ = _1159_ & ~_1158_;
	assign _1162_ = _1161_ ^ _3307_;
	assign _0116_ = _3331_ & ~_1162_;
	assign _1163_ = ~(\mchip.game2.score_inst.ctr [15] & \mchip.game2.score_inst.ctr [14]);
	assign _1164_ = _1163_ | _3311_;
	assign _1165_ = ~(_1164_ | _1153_);
	assign _1166_ = ~(_1165_ & _1144_);
	assign _1167_ = _1166_ ^ \mchip.game2.score_inst.ctr [16];
	assign _0117_ = _3331_ & ~_1167_;
	assign _1168_ = _1166_ | ~\mchip.game2.score_inst.ctr [16];
	assign _1169_ = _1168_ ^ \mchip.game2.score_inst.ctr [17];
	assign _0118_ = _3331_ & ~_1169_;
	assign _1170_ = ~(_1166_ | _3306_);
	assign _1171_ = ~(_1170_ ^ \mchip.game2.score_inst.ctr [18]);
	assign _0119_ = _3331_ & ~_1171_;
	assign _1172_ = ~(_1170_ & \mchip.game2.score_inst.ctr [18]);
	assign _1173_ = _1172_ ^ \mchip.game2.score_inst.ctr [19];
	assign _0120_ = _3331_ & ~_1173_;
	assign _1174_ = ~(\mchip.game2.score_inst.ctr [18] & \mchip.game2.score_inst.ctr [19]);
	assign _1175_ = _1174_ | _3306_;
	assign _1176_ = ~(_1175_ | _1166_);
	assign _1177_ = ~(_1176_ ^ \mchip.game2.score_inst.ctr [20]);
	assign _0122_ = _3331_ & ~_1177_;
	assign _1178_ = ~(_1176_ & \mchip.game2.score_inst.ctr [20]);
	assign _1179_ = _1178_ ^ \mchip.game2.score_inst.ctr [21];
	assign _0123_ = _3331_ & ~_1179_;
	assign _0106_ = _3362_ & ~\mchip.game2.score_inst.score[0] [0];
	assign _1180_ = _3359_ & _3351_;
	assign _0107_ = _3362_ & ~_1180_;
	assign _0108_ = _3362_ & _3352_;
	assign _0109_ = _3362_ & ~_3350_;
	assign _0102_ = ~(_3347_ | \mchip.game2.score_inst.score[1] [0]);
	assign _1181_ = _3344_ & _3336_;
	assign _0103_ = ~(_1181_ | _3347_);
	assign _0104_ = _3337_ & ~_3347_;
	assign _0105_ = _3335_ & ~_3347_;
	assign _0098_ = ~(_3379_ | \mchip.game2.score_inst.score[2] [0]);
	assign _1182_ = _3376_ & _3368_;
	assign _0099_ = ~(_1182_ | _3379_);
	assign _0100_ = _3369_ & ~_3379_;
	assign _0101_ = _3367_ & ~_3379_;
	assign _1183_ = \mchip.game2.score_inst.score[3] [0] & \mchip.game2.score_inst.score[3] [1];
	assign _1184_ = _1183_ & \mchip.game2.score_inst.score[3] [2];
	assign _1185_ = _1184_ ^ \mchip.game2.score_inst.score[3] [3];
	assign _1186_ = _1183_ ^ \mchip.game2.score_inst.score[3] [2];
	assign _1187_ = _1185_ & ~_1186_;
	assign _1188_ = \mchip.game2.score_inst.score[3] [1] & ~\mchip.game2.score_inst.score[3] [0];
	assign _1189_ = _1187_ & ~_1188_;
	assign _1190_ = _1185_ & ~_1189_;
	assign _1191_ = ~(\mchip.game2.score_inst.score[3] [3] & \mchip.game2.score_inst.score[3] [2]);
	assign _1192_ = _1183_ & ~_1191_;
	assign _1193_ = _1192_ | _1190_;
	assign _1194_ = \mchip.game2.score_inst.score[3] [0] & ~\mchip.game2.score_inst.score[3] [1];
	assign _1195_ = ~(_1194_ & _1187_);
	assign _1196_ = ~(_1195_ | _1192_);
	assign _1197_ = _1196_ | _1193_;
	assign _0094_ = ~(_1197_ | \mchip.game2.score_inst.score[3] [0]);
	assign _1198_ = ~(_1194_ | _1188_);
	assign _0095_ = ~(_1198_ | _1197_);
	assign _0096_ = _1186_ & ~_1197_;
	assign _0097_ = _1185_ & ~_1197_;
	assign _3625_[4] = _0253_ ^ \mchip.game2.vga_inst.haddr [4];
	assign _1199_ = ~\mchip.game2.vga_inst.haddr [4];
	assign _1200_ = _3179_ & ~_0248_;
	assign _1201_ = _1199_ & ~_1200_;
	assign _1202_ = _1201_ ^ \mchip.game2.vga_inst.haddr [5];
	assign _1203_ = \mchip.game2.score_inst.score_saved[3] [2] & \mchip.game2.score_inst.score_saved[3] [3];
	assign _1204_ = ~(\mchip.game2.score_inst.score_saved[3] [0] ^ \mchip.game2.score_inst.score_saved[3] [3]);
	assign _1205_ = _1204_ ^ _1203_;
	assign _1206_ = ~(\mchip.game2.score_inst.score_saved[3] [2] & \mchip.game2.score_inst.score_saved[3] [1]);
	assign _1207_ = ~(\mchip.game2.score_inst.score_saved[3] [2] ^ \mchip.game2.score_inst.score_saved[3] [3]);
	assign _1208_ = _1207_ | _1206_;
	assign _1209_ = _1207_ ^ _1206_;
	assign _1210_ = ~(\mchip.game2.score_inst.score_saved[3] [1] & \mchip.game2.score_inst.score_saved[3] [0]);
	assign _1211_ = ~(\mchip.game2.score_inst.score_saved[3] [2] ^ \mchip.game2.score_inst.score_saved[3] [1]);
	assign _1212_ = _1211_ | _1210_;
	assign _1213_ = _1209_ & ~_1212_;
	assign _1214_ = _1208_ & ~_1213_;
	assign _1215_ = ~(_1214_ | _1205_);
	assign _1216_ = _1203_ & ~_1204_;
	assign _1217_ = ~\mchip.game2.score_inst.score_saved[3] [1];
	assign _1218_ = \mchip.game2.score_inst.score_saved[3] [0] & \mchip.game2.score_inst.score_saved[3] [3];
	assign _1219_ = _1218_ ^ _1217_;
	assign _1220_ = _1219_ ^ _1216_;
	assign _1221_ = ~(_1220_ ^ _1215_);
	assign _1222_ = ~(_1221_ & _1202_);
	assign _1223_ = _1200_ ^ _1199_;
	assign _1224_ = ~_1223_;
	assign _1225_ = _1214_ ^ _1205_;
	assign _1226_ = _1225_ & ~_1224_;
	assign _1227_ = _1221_ ^ _1202_;
	assign _1228_ = ~(_1227_ & _1226_);
	assign _1229_ = ~(_1228_ & _1222_);
	assign _1230_ = _1225_ ^ _1224_;
	assign _1231_ = _1227_ & ~_1230_;
	assign _1232_ = ~\mchip.game2.vga_inst.haddr [2];
	assign _1233_ = _3179_ & ~_1232_;
	assign _1234_ = _1233_ ^ \mchip.game2.vga_inst.haddr [3];
	assign _1235_ = ~(_1212_ ^ _1209_);
	assign _1236_ = ~(_1235_ & _1234_);
	assign _1237_ = ~(_1235_ ^ _1234_);
	assign _1238_ = _1232_ & ~_3179_;
	assign _1239_ = ~(_1238_ | _1233_);
	assign _1240_ = _1211_ ^ _1210_;
	assign _1241_ = ~(_1240_ & _1239_);
	assign _1242_ = ~(_1241_ | _1237_);
	assign _1243_ = _1236_ & ~_1242_;
	assign _1244_ = _1240_ ^ _1239_;
	assign _1245_ = _1244_ & ~_1237_;
	assign _1246_ = ~(\mchip.game2.score_inst.score_saved[3] [1] ^ \mchip.game2.score_inst.score_saved[3] [0]);
	assign _3625_[1] = _3179_ & ~_0241_;
	assign _1247_ = _3625_[1] | _1246_;
	assign _1248_ = \mchip.game2.score_inst.score_saved[3] [0] & ~\mchip.game2.vga_inst.haddr [0];
	assign _1249_ = _3625_[1] ^ _1246_;
	assign _1250_ = _1249_ & _1248_;
	assign _1251_ = _1247_ & ~_1250_;
	assign _1252_ = _1245_ & ~_1251_;
	assign _1253_ = _1243_ & ~_1252_;
	assign _1254_ = _1231_ & ~_1253_;
	assign _1255_ = _1254_ | _1229_;
	assign _1256_ = ~\mchip.game2.vga_inst.haddr [6];
	assign _1257_ = _0239_ & ~_1200_;
	assign _1258_ = _1257_ ^ _1256_;
	assign _1259_ = _1216_ & ~_1219_;
	assign _1260_ = _1220_ | _1205_;
	assign _1261_ = ~(_1260_ | _1214_);
	assign _1262_ = _1261_ | _1259_;
	assign _1263_ = _1218_ & ~_1217_;
	assign _1264_ = _1263_ ^ \mchip.game2.score_inst.score_saved[3] [2];
	assign _1265_ = _1264_ ^ _1262_;
	assign _1266_ = _1265_ ^ _1258_;
	assign _1267_ = _1266_ ^ _1255_;
	assign _1268_ = ~(\mchip.game2.score_inst.score_saved[3] [0] ^ \mchip.game2.vga_inst.haddr [0]);
	assign _1269_ = ~\mchip.game2.vga_inst.haddr [8];
	assign _1270_ = \mchip.game2.vga_inst.haddr [6] & \mchip.game2.vga_inst.haddr [7];
	assign _1271_ = _0239_ | ~_1270_;
	assign _1272_ = _1270_ & _0239_;
	assign _1273_ = _1272_ & _1200_;
	assign _1274_ = _1271_ & ~_1273_;
	assign _1275_ = _1274_ ^ _1269_;
	assign _1276_ = ~_1275_;
	assign _1277_ = ~\mchip.game2.score_inst.score_saved[3] [3];
	assign _1278_ = ~(_1263_ & \mchip.game2.score_inst.score_saved[3] [2]);
	assign _1279_ = _1278_ | _1277_;
	assign _1280_ = ~(_1264_ & \mchip.game2.score_inst.score_saved[3] [3]);
	assign _1281_ = _1259_ & ~_1280_;
	assign _1282_ = _1279_ & ~_1281_;
	assign _1283_ = _1280_ | _1260_;
	assign _1284_ = ~(_1283_ | _1214_);
	assign _1285_ = _1282_ & ~_1284_;
	assign _1286_ = _1285_ | _1276_;
	assign _1287_ = \mchip.game2.vga_inst.haddr [6] & ~_1257_;
	assign _1288_ = _1287_ ^ \mchip.game2.vga_inst.haddr [7];
	assign _1289_ = ~_1288_;
	assign _1290_ = ~(_1264_ & _1262_);
	assign _1291_ = _1290_ & _1278_;
	assign _1292_ = _1291_ ^ _1277_;
	assign _1293_ = _1292_ & ~_1289_;
	assign _1294_ = _1265_ & _1258_;
	assign _1295_ = _1292_ ^ _1289_;
	assign _1296_ = _1294_ & ~_1295_;
	assign _1297_ = _1296_ | _1293_;
	assign _1298_ = _1295_ | ~_1266_;
	assign _1299_ = _1229_ & ~_1298_;
	assign _1300_ = _1299_ | _1297_;
	assign _1301_ = _1298_ | ~_1231_;
	assign _1302_ = ~(_1301_ | _1253_);
	assign _1303_ = _1302_ | _1300_;
	assign _1304_ = _1285_ ^ _1276_;
	assign _1305_ = _1304_ & _1303_;
	assign _1306_ = _1286_ & ~_1305_;
	assign _1307_ = ~\mchip.game2.vga_inst.haddr [9];
	assign _1308_ = \mchip.game2.vga_inst.haddr [8] & ~_1274_;
	assign _1309_ = _1308_ ^ _1307_;
	assign _1310_ = _1309_ ^ _1306_;
	assign _1311_ = \mchip.game2.vga_inst.vaddr [2] & ~_3219_;
	assign _1312_ = _1311_ ^ _0519_;
	assign _1313_ = _1312_ & ~_0630_;
	assign _1314_ = ~(_0404_ | _3219_);
	assign _1315_ = _0519_ & ~_1314_;
	assign _1316_ = ~(_1315_ ^ \mchip.game2.vga_inst.vaddr [4]);
	assign _1317_ = _1316_ | _1313_;
	assign _1318_ = \mchip.game2.vga_inst.vaddr [4] & ~_1315_;
	assign _1319_ = _1318_ ^ \mchip.game2.vga_inst.vaddr [5];
	assign _1320_ = _0629_ & _0586_;
	assign _1321_ = ~(_1320_ & _1312_);
	assign _1322_ = _1321_ | ~_1316_;
	assign _1323_ = (_1319_ ? _1322_ : _1317_);
	assign _1324_ = _1323_ | ~_1310_;
	assign _1325_ = _1324_ | _1268_;
	assign _1326_ = _1249_ ^ _1248_;
	assign _1327_ = _1326_ | _1325_;
	assign _1328_ = ~(_1251_ ^ _1244_);
	assign _1329_ = _3219_ | _0516_;
	assign _1330_ = ~(_1329_ & _1312_);
	assign _1331_ = _1330_ | ~_1316_;
	assign _1332_ = _0586_ & ~_0497_;
	assign _1333_ = _1332_ & _1312_;
	assign _1334_ = _1333_ | _1316_;
	assign _1335_ = (_1319_ ? _1331_ : _1334_);
	assign _1336_ = _1335_ | ~_1310_;
	assign _1337_ = (_1326_ ? _1324_ : _1336_);
	assign _1338_ = (_1328_ ? _1327_ : _1337_);
	assign _1339_ = _1244_ & ~_1251_;
	assign _1340_ = _1241_ & ~_1339_;
	assign _1341_ = _1340_ ^ _1237_;
	assign _1342_ = ~_3219_;
	assign _1343_ = (_0586_ ? _0629_ : _1342_);
	assign _1344_ = _1343_ | ~_1312_;
	assign _1345_ = _1344_ | ~_1316_;
	assign _1346_ = _0516_ & ~_3219_;
	assign _1347_ = (_1312_ ? _1332_ : _1346_);
	assign _1348_ = _1316_ | ~_1347_;
	assign _1349_ = (_1319_ ? _1345_ : _1348_);
	assign _1350_ = _1310_ & ~_1349_;
	assign _1351_ = ~_1350_;
	assign _1352_ = (_1319_ ? _1331_ : _1316_);
	assign _1353_ = _1310_ & ~_1352_;
	assign _1354_ = ~_1353_;
	assign _1355_ = ~_1346_;
	assign _1356_ = (_1312_ ? _0630_ : _1355_);
	assign _1357_ = _1356_ | _1316_;
	assign _1358_ = (_1319_ ? _1345_ : _1357_);
	assign _1359_ = _1358_ | ~_1310_;
	assign _1360_ = (_1268_ ? _1354_ : _1359_);
	assign _1361_ = (_1268_ ? _1359_ : _1351_);
	assign _1362_ = (_1326_ ? _1360_ : _1361_);
	assign _1363_ = (_1328_ ? _1362_ : _1351_);
	assign _1364_ = (_1341_ ? _1338_ : _1363_);
	assign _1365_ = _1253_ ^ _1230_;
	assign _1366_ = _3219_ & ~_0516_;
	assign _1367_ = ~_1366_;
	assign _1368_ = (_1312_ ? _1332_ : _1367_);
	assign _1369_ = _1316_ | ~_1368_;
	assign _1370_ = (_1319_ ? _1331_ : _1369_);
	assign _1371_ = _1310_ & ~_1370_;
	assign _1372_ = ~_1371_;
	assign _1373_ = ~_0586_;
	assign _1374_ = _1373_ & ~_1312_;
	assign _1375_ = _1316_ | ~_1374_;
	assign _1376_ = (_1319_ ? _1322_ : _1375_);
	assign _1377_ = _1376_ | ~_1310_;
	assign _1378_ = (_1268_ ? _1372_ : _1377_);
	assign _1379_ = (_1326_ ? _1372_ : _1378_);
	assign _1380_ = _1377_ | ~_1268_;
	assign _1381_ = _1368_ | _1316_;
	assign _1382_ = _1381_ | _1319_;
	assign _1383_ = _1382_ | ~_1310_;
	assign _1384_ = (_1326_ ? _1380_ : _1383_);
	assign _1385_ = (_1328_ ? _1379_ : _1384_);
	assign _1386_ = _1346_ & ~_1312_;
	assign _1387_ = _1386_ | _1316_;
	assign _1388_ = (_1319_ ? _1322_ : _1387_);
	assign _1389_ = _1388_ | ~_1310_;
	assign _1390_ = (_1268_ ? _1383_ : _1389_);
	assign _1391_ = (_1268_ ? _1389_ : _1354_);
	assign _1392_ = (_1326_ ? _1390_ : _1391_);
	assign _1393_ = ~_1312_;
	assign _1394_ = _1332_ | _0630_;
	assign _1395_ = (_1312_ ? _1394_ : _0586_);
	assign _1396_ = _1316_ | ~_1395_;
	assign _1397_ = (_1319_ ? _1345_ : _1396_);
	assign _1398_ = _1310_ & ~_1397_;
	assign _1399_ = ~_1398_;
	assign _1400_ = (_1328_ ? _1392_ : _1399_);
	assign _1401_ = (_1341_ ? _1385_ : _1400_);
	assign _1402_ = (_1365_ ? _1364_ : _1401_);
	assign _1403_ = ~(_1253_ | _1230_);
	assign _1404_ = _1403_ | _1226_;
	assign _1405_ = _1404_ ^ _1227_;
	assign _1406_ = ~(_1394_ | _1393_);
	assign _1407_ = _0626_ & ~_1312_;
	assign _1408_ = _1407_ | _1406_;
	assign _1409_ = _1408_ | _1316_;
	assign _1410_ = (_1319_ ? _1345_ : _1409_);
	assign _1411_ = _1310_ & ~_1410_;
	assign _1412_ = ~_1411_;
	assign _1413_ = \mchip.game2.vga_inst.vaddr [1] | ~\mchip.game2.vga_inst.vaddr [2];
	assign _1414_ = (_1312_ ? _1332_ : _1413_);
	assign _1415_ = _1316_ | ~_1414_;
	assign _1416_ = (_1319_ ? _1345_ : _1415_);
	assign _1417_ = _1310_ & ~_1416_;
	assign _1418_ = ~_1417_;
	assign _1419_ = (_1268_ ? _1412_ : _1418_);
	assign _1420_ = (_1268_ ? _1418_ : _1372_);
	assign _1421_ = (_1326_ ? _1419_ : _1420_);
	assign _1422_ = (_1268_ ? _1372_ : _1354_);
	assign _1423_ = _1347_ | _1316_;
	assign _1424_ = (_1319_ ? _1322_ : _1423_);
	assign _1425_ = _1424_ | ~_1310_;
	assign _1426_ = (_1326_ ? _1422_ : _1425_);
	assign _1427_ = (_1328_ ? _1421_ : _1426_);
	assign _1428_ = _1316_ | ~_1407_;
	assign _1429_ = (_1319_ ? _1331_ : _1428_);
	assign _1430_ = _1429_ | ~_1310_;
	assign _1431_ = _1430_ | _1268_;
	assign _1432_ = (_1326_ ? _1431_ : _1430_);
	assign _1433_ = (_1319_ ? _1331_ : _1375_);
	assign _1434_ = _1433_ | ~_1310_;
	assign _1435_ = _1367_ & ~_1312_;
	assign _1436_ = _1316_ | ~_1435_;
	assign _1437_ = (_1319_ ? _1331_ : _1436_);
	assign _1438_ = _1437_ | ~_1310_;
	assign _1439_ = _1413_ & ~_1312_;
	assign _1440_ = _1316_ | ~_1439_;
	assign _1441_ = (_1319_ ? _1345_ : _1440_);
	assign _1442_ = _1441_ | ~_1310_;
	assign _1443_ = (_1268_ ? _1438_ : _1442_);
	assign _1444_ = (_1326_ ? _1434_ : _1443_);
	assign _1445_ = (_1328_ ? _1432_ : _1444_);
	assign _1446_ = (_1341_ ? _1427_ : _1445_);
	assign _1447_ = _1374_ | _1316_;
	assign _1448_ = (_1319_ ? _1345_ : _1447_);
	assign _1449_ = _1310_ & ~_1448_;
	assign _1450_ = ~_1449_;
	assign _1451_ = (_1268_ ? _1442_ : _1450_);
	assign _1452_ = (_1326_ ? _1451_ : _1450_);
	assign _1453_ = _1435_ | _1316_;
	assign _1454_ = (_1319_ ? _1345_ : _1453_);
	assign _1455_ = _1454_ | ~_1310_;
	assign _1456_ = (_1326_ ? _1455_ : _1430_);
	assign _1457_ = (_1328_ ? _1452_ : _1456_);
	assign _1458_ = _1430_ | ~_1268_;
	assign _1459_ = (_1326_ ? _1430_ : _1458_);
	assign _1460_ = (_1268_ ? _1383_ : _1450_);
	assign _1461_ = (_1326_ ? _1383_ : _1460_);
	assign _1462_ = (_1328_ ? _1459_ : _1461_);
	assign _1463_ = (_1341_ ? _1457_ : _1462_);
	assign _1464_ = (_1365_ ? _1446_ : _1463_);
	assign _1465_ = (_1405_ ? _1402_ : _1464_);
	assign _1466_ = ~(_1465_ | _1267_);
	assign _1467_ = ~(_1266_ & _1255_);
	assign _1468_ = _1467_ & ~_1294_;
	assign _1469_ = _1468_ ^ _1295_;
	assign _1470_ = (_1326_ ? _1449_ : _1350_);
	assign _1471_ = (\mchip.game2.vga_inst.vaddr [1] ? _0516_ : \mchip.game2.vga_inst.vaddr [0]);
	assign _1472_ = (_1312_ ? _1332_ : _1471_);
	assign _1473_ = _1316_ | ~_1472_;
	assign _1474_ = (_1319_ ? _1331_ : _1473_);
	assign _1475_ = _1310_ & ~_1474_;
	assign _1476_ = (_1326_ ? _1350_ : _1475_);
	assign _1477_ = (_1328_ ? _1470_ : _1476_);
	assign _1478_ = (_1319_ ? _1322_ : _1316_);
	assign _1479_ = _1310_ & ~_1478_;
	assign _1480_ = (_1268_ ? _1475_ : _1479_);
	assign _1481_ = (_1326_ ? _1480_ : _1479_);
	assign _1482_ = ~(_1407_ | _1333_);
	assign _1483_ = _1316_ | ~_1482_;
	assign _1484_ = ~(_1483_ | _1319_);
	assign _1485_ = ~_1484_;
	assign _1486_ = _1310_ & ~_1485_;
	assign _1487_ = (_1312_ ? _1332_ : _1373_);
	assign _1488_ = _1487_ | _1316_;
	assign _1489_ = _1488_ | _1319_;
	assign _1490_ = _1310_ & ~_1489_;
	assign _1491_ = _1490_ & ~_1268_;
	assign _1492_ = (_1326_ ? _1486_ : _1491_);
	assign _1493_ = (_1328_ ? _1481_ : _1492_);
	assign _1494_ = (_1341_ ? _1477_ : _1493_);
	assign _1495_ = _1407_ | _1316_;
	assign _1496_ = (_1319_ ? _1345_ : _1495_);
	assign _1497_ = _1310_ & ~_1496_;
	assign _1498_ = (_1326_ ? _1490_ : _1497_);
	assign _1499_ = ~_1332_;
	assign _1500_ = _0586_ | _0497_;
	assign _1501_ = (_1312_ ? _1499_ : _1500_);
	assign _1502_ = _1501_ | _1316_;
	assign _1503_ = (_1319_ ? _1345_ : _1502_);
	assign _1504_ = _1310_ & ~_1503_;
	assign _1505_ = (_1268_ ? _1497_ : _1504_);
	assign _1506_ = (_1326_ ? _1505_ : _1504_);
	assign _1507_ = (_1328_ ? _1498_ : _1506_);
	assign _1508_ = (_1312_ ? _0630_ : _0586_);
	assign _1509_ = _1508_ | _1316_;
	assign _1510_ = (_1319_ ? _1331_ : _1509_);
	assign _1511_ = _1310_ & ~_1510_;
	assign _1512_ = _1395_ | _1316_;
	assign _1513_ = (_1319_ ? _1331_ : _1512_);
	assign _1514_ = _1310_ & ~_1513_;
	assign _1515_ = (_1268_ ? _1511_ : _1514_);
	assign _1516_ = (_1326_ ? _1511_ : _1515_);
	assign _1517_ = (_1328_ ? _1504_ : _1516_);
	assign _1518_ = (_1341_ ? _1507_ : _1517_);
	assign _1519_ = (_1365_ ? _1494_ : _1518_);
	assign _1520_ = ~_1268_;
	assign _1521_ = _1514_ & ~_1520_;
	assign _1522_ = (_1312_ ? _0630_ : _1366_);
	assign _1523_ = _1316_ | ~_1522_;
	assign _1524_ = _1523_ | _1319_;
	assign _1525_ = _1310_ & ~_1524_;
	assign _1526_ = (_1326_ ? _1521_ : _1525_);
	assign _1527_ = (_1268_ ? _1525_ : _1353_);
	assign _1528_ = (_1326_ ? _1527_ : _1353_);
	assign _1529_ = (_1328_ ? _1526_ : _1528_);
	assign _1530_ = ~_1413_;
	assign _1531_ = (_1312_ ? _0630_ : _1530_);
	assign _1532_ = _1316_ | ~_1531_;
	assign _1533_ = (_1319_ ? _1331_ : _1532_);
	assign _1534_ = _1310_ & ~_1533_;
	assign _1535_ = (_1326_ ? _1353_ : _1534_);
	assign _1536_ = _1319_ & ~_1331_;
	assign _1537_ = _1356_ & ~_1316_;
	assign _1538_ = _1537_ & ~_1319_;
	assign _1539_ = ~(_1538_ | _1536_);
	assign _1540_ = _1310_ & ~_1539_;
	assign _1541_ = _1319_ & ~_1322_;
	assign _1542_ = ~(_1538_ | _1541_);
	assign _1543_ = _1310_ & ~_1542_;
	assign _1544_ = (_1268_ ? _1540_ : _1543_);
	assign _1545_ = ~(_1407_ | _1313_);
	assign _1546_ = _1316_ | ~_1545_;
	assign _1547_ = _1546_ | _1319_;
	assign _1548_ = _1310_ & ~_1547_;
	assign _1549_ = (_1268_ ? _1543_ : _1548_);
	assign _1550_ = (_1326_ ? _1544_ : _1549_);
	assign _1551_ = (_1328_ ? _1535_ : _1550_);
	assign _1552_ = (_1341_ ? _1529_ : _1551_);
	assign _1553_ = _1316_ | ~_1508_;
	assign _1554_ = ~(_1553_ | _1319_);
	assign _1555_ = ~_1554_;
	assign _1556_ = _1310_ & ~_1555_;
	assign _1557_ = (_1326_ ? _1548_ : _1556_);
	assign _1558_ = (_1319_ ? _1345_ : _1381_);
	assign _1559_ = _1310_ & ~_1558_;
	assign _1560_ = _1559_ & ~_1268_;
	assign _1561_ = (_1326_ ? _1560_ : _1559_);
	assign _1562_ = (_1328_ ? _1557_ : _1561_);
	assign _1563_ = ~(_1500_ | _1312_);
	assign _1564_ = _1563_ | _1316_;
	assign _1565_ = (_1319_ ? _1331_ : _1564_);
	assign _1566_ = _1310_ & ~_1565_;
	assign _1567_ = (_1268_ ? _1353_ : _1371_);
	assign _1568_ = (_1326_ ? _1566_ : _1567_);
	assign _1569_ = (_1268_ ? _1371_ : _1417_);
	assign _1570_ = (_1326_ ? _1569_ : _1417_);
	assign _1571_ = (_1328_ ? _1568_ : _1570_);
	assign _1572_ = (_1341_ ? _1562_ : _1571_);
	assign _1573_ = (_1365_ ? _1552_ : _1572_);
	assign _1574_ = (_1405_ ? _1519_ : _1573_);
	assign _1575_ = _1316_ | ~_1313_;
	assign _1576_ = (_1319_ ? _1345_ : _1575_);
	assign _1577_ = _1310_ & ~_1576_;
	assign _1578_ = (_1326_ ? _1350_ : _1577_);
	assign _1579_ = _1316_ | ~_1406_;
	assign _1580_ = _1579_ | _1319_;
	assign _1581_ = _1310_ & ~_1580_;
	assign _1582_ = (_1268_ ? _1577_ : _1581_);
	assign _1583_ = _1581_ & ~_1520_;
	assign _1584_ = (_1326_ ? _1582_ : _1583_);
	assign _1585_ = (_1328_ ? _1578_ : _1584_);
	assign _1586_ = _1316_ | ~_1487_;
	assign _1587_ = (_1319_ ? _1322_ : _1586_);
	assign _1588_ = _1310_ & ~_1587_;
	assign _1589_ = (_1268_ ? _1588_ : _1371_);
	assign _1590_ = (_1326_ ? _1588_ : _1589_);
	assign _1591_ = _1406_ | _1316_;
	assign _1592_ = (_1319_ ? _1331_ : _1591_);
	assign _1593_ = _1310_ & ~_1592_;
	assign _1594_ = (_1268_ ? _1371_ : _1593_);
	assign _1595_ = (_1326_ ? _1594_ : _1411_);
	assign _1596_ = (_1328_ ? _1590_ : _1595_);
	assign _1597_ = (_1341_ ? _1585_ : _1596_);
	assign _1598_ = (_1326_ ? _1398_ : _1449_);
	assign _1599_ = _1439_ | _1316_;
	assign _1600_ = (_1319_ ? _1331_ : _1599_);
	assign _1601_ = _1310_ & ~_1600_;
	assign _1602_ = (_1268_ ? _1449_ : _1601_);
	assign _1603_ = (_1326_ ? _1602_ : _1601_);
	assign _1604_ = (_1328_ ? _1598_ : _1603_);
	assign _1605_ = _1316_ | ~_1333_;
	assign _1606_ = _1605_ | _1319_;
	assign _1607_ = _1310_ & ~_1606_;
	assign _1608_ = _1545_ | _1316_;
	assign _1609_ = (_1319_ ? _1322_ : _1608_);
	assign _1610_ = _1310_ & ~_1609_;
	assign _1611_ = _1607_ & ~_1268_;
	assign _1612_ = (_1326_ ? _1610_ : _1611_);
	assign _1613_ = (_1328_ ? _1612_ : _1607_);
	assign _1614_ = (_1341_ ? _1604_ : _1613_);
	assign _1615_ = (_1365_ ? _1597_ : _1614_);
	assign _1616_ = _1482_ | _1316_;
	assign _1617_ = (_1319_ ? _1322_ : _1616_);
	assign _1618_ = _1310_ & ~_1617_;
	assign _1619_ = (_1326_ ? _1353_ : _1618_);
	assign _1620_ = (_1328_ ? _1353_ : _1619_);
	assign _1621_ = _1607_ & ~_1520_;
	assign _1622_ = (_1326_ ? _1607_ : _1621_);
	assign _1623_ = _1548_ & ~_1326_;
	assign _1624_ = (_1328_ ? _1622_ : _1623_);
	assign _1625_ = (_1341_ ? _1620_ : _1624_);
	assign _1626_ = (_1319_ ? _1322_ : _1334_);
	assign _1627_ = _1310_ & ~_1626_;
	assign _1628_ = (_1268_ ? _1548_ : _1627_);
	assign _1629_ = (_1268_ ? _1627_ : _1353_);
	assign _1630_ = (_1326_ ? _1628_ : _1629_);
	assign _1631_ = (_1319_ ? _1331_ : _1616_);
	assign _1632_ = (_1319_ ? _1345_ : _1605_);
	assign _1633_ = (_1326_ ? _1631_ : _1632_);
	assign _1634_ = _1310_ & ~_1633_;
	assign _1635_ = (_1328_ ? _1630_ : _1634_);
	assign _1636_ = (_1268_ ? _1577_ : _1627_);
	assign _1637_ = (_1326_ ? _1577_ : _1636_);
	assign _1638_ = (_1326_ ? _1627_ : _1548_);
	assign _1639_ = (_1328_ ? _1637_ : _1638_);
	assign _1640_ = (_1341_ ? _1635_ : _1639_);
	assign _1641_ = (_1365_ ? _1625_ : _1640_);
	assign _1642_ = (_1405_ ? _1615_ : _1641_);
	assign _1643_ = (_1267_ ? _1574_ : _1642_);
	assign _1644_ = (_1469_ ? _1466_ : _1643_);
	assign _1645_ = _1304_ ^ _1303_;
	assign _1646_ = _1644_ & ~_1645_;
	assign _1647_ = \mchip.game2.vga_inst.haddr [8] & ~\mchip.game2.vga_inst.haddr [9];
	assign _1648_ = ~_1647_;
	assign _1649_ = _1270_ & _3178_;
	assign _1650_ = _3185_ & ~_3179_;
	assign _1651_ = ~(_1650_ & _1649_);
	assign _1652_ = _1651_ | _1648_;
	assign _1653_ = ~_0237_;
	assign _1654_ = _1270_ & ~_0771_;
	assign _1655_ = _1654_ & _1651_;
	assign _1656_ = _1647_ & ~_1655_;
	assign _1657_ = _1653_ & ~_1656_;
	assign _1658_ = _1652_ & ~_1657_;
	assign _1659_ = _1272_ & ~_1200_;
	assign _1660_ = _1270_ & ~_1659_;
	assign _1661_ = _1647_ & ~_1660_;
	assign _1662_ = _1661_ | _0237_;
	assign _1663_ = _1658_ & ~_1662_;
	assign _1664_ = _3185_ & ~_0241_;
	assign _1665_ = _1664_ & ~\mchip.game2.vga_inst.haddr [4];
	assign _1666_ = _1665_ ^ _0771_;
	assign _1667_ = ~_1666_;
	assign _1668_ = ~(\mchip.game2.score_inst.score_saved[2] [1] & \mchip.game2.score_inst.score_saved[2] [2]);
	assign _1669_ = ~\mchip.game2.score_inst.score_saved[2] [3];
	assign _1670_ = \mchip.game2.score_inst.score_saved[2] [2] & ~\mchip.game2.score_inst.score_saved[2] [1];
	assign _1671_ = _1670_ & ~_1669_;
	assign _1672_ = _1671_ | ~_1668_;
	assign _1673_ = ~(\mchip.game2.score_inst.score_saved[2] [0] ^ \mchip.game2.score_inst.score_saved[2] [3]);
	assign _1674_ = _1672_ & ~_1673_;
	assign _1675_ = \mchip.game2.score_inst.score_saved[2] [1] & \mchip.game2.score_inst.score_saved[2] [0];
	assign _1676_ = ~(\mchip.game2.score_inst.score_saved[2] [1] ^ \mchip.game2.score_inst.score_saved[2] [2]);
	assign _1677_ = _1675_ & ~_1676_;
	assign _1678_ = _1670_ ^ _1669_;
	assign _1679_ = _1677_ & ~_1678_;
	assign _1680_ = _1673_ ^ _1672_;
	assign _1681_ = _1679_ & ~_1680_;
	assign _1682_ = _1681_ | _1674_;
	assign _1683_ = \mchip.game2.score_inst.score_saved[2] [0] & \mchip.game2.score_inst.score_saved[2] [3];
	assign _1684_ = ~(_1683_ ^ \mchip.game2.score_inst.score_saved[2] [1]);
	assign _1685_ = ~(_1684_ ^ _1682_);
	assign _1686_ = _1685_ & ~_1667_;
	assign _1687_ = _1685_ ^ _1667_;
	assign _1688_ = _1664_ ^ _1199_;
	assign _1689_ = ~(_1680_ ^ _1679_);
	assign _1690_ = _1688_ | ~_1689_;
	assign _1691_ = ~(_1690_ | _1687_);
	assign _1692_ = _1691_ | _1686_;
	assign _1693_ = _1689_ ^ _1688_;
	assign _1694_ = _1693_ | _1687_;
	assign _1695_ = _1232_ & ~_0241_;
	assign _1696_ = _1695_ ^ \mchip.game2.vga_inst.haddr [3];
	assign _1697_ = ~(_1678_ ^ _1677_);
	assign _1698_ = ~(_1697_ & _1696_);
	assign _1699_ = ~(_1697_ ^ _1696_);
	assign _1700_ = _0241_ ^ _1232_;
	assign _1701_ = ~(_1676_ ^ _1675_);
	assign _1702_ = ~(_1701_ & _1700_);
	assign _1703_ = ~(_1702_ | _1699_);
	assign _1704_ = _1698_ & ~_1703_;
	assign _1705_ = _1701_ ^ _1700_;
	assign _1706_ = _1705_ & ~_1699_;
	assign _1707_ = \mchip.game2.score_inst.score_saved[2] [1] ^ \mchip.game2.score_inst.score_saved[2] [0];
	assign _1708_ = ~(_1707_ & _3625_[1]);
	assign _1709_ = \mchip.game2.score_inst.score_saved[2] [0] & ~\mchip.game2.vga_inst.haddr [0];
	assign _1710_ = _1707_ ^ _3625_[1];
	assign _1711_ = _1710_ & _1709_;
	assign _1712_ = _1708_ & ~_1711_;
	assign _1713_ = _1706_ & ~_1712_;
	assign _1714_ = _1704_ & ~_1713_;
	assign _1715_ = ~(_1714_ | _1694_);
	assign _1716_ = _1715_ | _1692_;
	assign _1717_ = ~(\mchip.game2.vga_inst.haddr [4] & \mchip.game2.vga_inst.haddr [5]);
	assign _1718_ = _3178_ & ~_1664_;
	assign _1719_ = _1717_ & ~_1718_;
	assign _1720_ = _1719_ ^ _1256_;
	assign _1721_ = ~(_1683_ & \mchip.game2.score_inst.score_saved[2] [1]);
	assign _1722_ = _1674_ & ~_1684_;
	assign _1723_ = _1721_ & ~_1722_;
	assign _1724_ = _1684_ | _1680_;
	assign _1725_ = _1679_ & ~_1724_;
	assign _1726_ = _1723_ & ~_1725_;
	assign _1727_ = _1726_ ^ \mchip.game2.score_inst.score_saved[2] [2];
	assign _1728_ = _1727_ ^ _1720_;
	assign _1729_ = ~(_1728_ ^ _1716_);
	assign _1730_ = ~(\mchip.game2.score_inst.score_saved[2] [0] ^ \mchip.game2.vga_inst.haddr [0]);
	assign _1731_ = _1270_ & ~_1717_;
	assign _1732_ = ~_1731_;
	assign _1733_ = _1649_ & ~_1664_;
	assign _1734_ = _1732_ & ~_1733_;
	assign _1735_ = _1734_ ^ _1269_;
	assign _1736_ = ~(\mchip.game2.score_inst.score_saved[2] [2] & \mchip.game2.score_inst.score_saved[2] [3]);
	assign _1737_ = _1736_ | _1723_;
	assign _1738_ = _1736_ | _1724_;
	assign _1739_ = _1679_ & ~_1738_;
	assign _1740_ = _1737_ & ~_1739_;
	assign _1741_ = _1735_ & ~_1740_;
	assign _1742_ = \mchip.game2.vga_inst.haddr [6] & ~_1719_;
	assign _1743_ = _1742_ ^ \mchip.game2.vga_inst.haddr [7];
	assign _1744_ = ~_1743_;
	assign _1745_ = \mchip.game2.score_inst.score_saved[2] [2] & ~_1726_;
	assign _1746_ = _1745_ ^ \mchip.game2.score_inst.score_saved[2] [3];
	assign _1747_ = _1746_ & ~_1744_;
	assign _1748_ = _1720_ & ~_1727_;
	assign _1749_ = _1746_ ^ _1744_;
	assign _1750_ = _1748_ & ~_1749_;
	assign _1751_ = _1750_ | _1747_;
	assign _1752_ = _1749_ | _1728_;
	assign _1753_ = _1692_ & ~_1752_;
	assign _1754_ = _1753_ | _1751_;
	assign _1755_ = _1752_ | _1694_;
	assign _1756_ = ~(_1755_ | _1714_);
	assign _1757_ = _1756_ | _1754_;
	assign _1758_ = ~(_1740_ ^ _1735_);
	assign _1759_ = _1758_ & _1757_;
	assign _1760_ = _1759_ | _1741_;
	assign _1761_ = \mchip.game2.vga_inst.haddr [8] & ~_1734_;
	assign _1762_ = _1761_ ^ _1307_;
	assign _1763_ = _1762_ ^ _1760_;
	assign _1764_ = _1763_ | _1323_;
	assign _1765_ = _1764_ | _1730_;
	assign _1766_ = _1710_ ^ _1709_;
	assign _1767_ = _1766_ | _1765_;
	assign _1768_ = ~(_1712_ ^ _1705_);
	assign _1769_ = _1763_ | _1335_;
	assign _1770_ = (_1766_ ? _1764_ : _1769_);
	assign _1771_ = (_1768_ ? _1767_ : _1770_);
	assign _1772_ = _1705_ & ~_1712_;
	assign _1773_ = _1702_ & ~_1772_;
	assign _1774_ = _1773_ ^ _1699_;
	assign _1775_ = ~(_1763_ | _1349_);
	assign _1776_ = ~_1775_;
	assign _1777_ = ~(_1763_ | _1352_);
	assign _1778_ = ~_1777_;
	assign _1779_ = _1763_ | _1358_;
	assign _1780_ = (_1730_ ? _1778_ : _1779_);
	assign _1781_ = (_1730_ ? _1779_ : _1776_);
	assign _1782_ = (_1766_ ? _1780_ : _1781_);
	assign _1783_ = (_1768_ ? _1782_ : _1776_);
	assign _1784_ = (_1774_ ? _1771_ : _1783_);
	assign _1785_ = _1714_ ^ _1693_;
	assign _1786_ = ~(_1763_ | _1370_);
	assign _1787_ = ~_1786_;
	assign _1788_ = _1763_ | _1376_;
	assign _1789_ = (_1730_ ? _1787_ : _1788_);
	assign _1790_ = (_1766_ ? _1787_ : _1789_);
	assign _1791_ = _1788_ | ~_1730_;
	assign _1792_ = _1763_ | _1382_;
	assign _1793_ = (_1766_ ? _1791_ : _1792_);
	assign _1794_ = (_1768_ ? _1790_ : _1793_);
	assign _1795_ = _1763_ | _1388_;
	assign _1796_ = (_1730_ ? _1792_ : _1795_);
	assign _1797_ = (_1730_ ? _1795_ : _1778_);
	assign _1798_ = (_1766_ ? _1796_ : _1797_);
	assign _1799_ = ~(_1763_ | _1397_);
	assign _1800_ = ~_1799_;
	assign _1801_ = (_1768_ ? _1798_ : _1800_);
	assign _1802_ = (_1774_ ? _1794_ : _1801_);
	assign _1803_ = (_1785_ ? _1784_ : _1802_);
	assign _1804_ = ~(_1714_ | _1693_);
	assign _1805_ = _1690_ & ~_1804_;
	assign _1806_ = _1805_ ^ _1687_;
	assign _1807_ = ~(_1763_ | _1410_);
	assign _1808_ = ~_1807_;
	assign _1809_ = ~(_1763_ | _1416_);
	assign _1810_ = ~_1809_;
	assign _1811_ = (_1730_ ? _1808_ : _1810_);
	assign _1812_ = (_1730_ ? _1810_ : _1787_);
	assign _1813_ = (_1766_ ? _1811_ : _1812_);
	assign _1814_ = (_1730_ ? _1787_ : _1778_);
	assign _1815_ = _1763_ | _1424_;
	assign _1816_ = (_1766_ ? _1814_ : _1815_);
	assign _1817_ = (_1768_ ? _1813_ : _1816_);
	assign _1818_ = _1763_ | _1429_;
	assign _1819_ = _1818_ | _1730_;
	assign _1820_ = (_1766_ ? _1819_ : _1818_);
	assign _1821_ = _1763_ | _1433_;
	assign _1822_ = _1763_ | _1437_;
	assign _1823_ = _1763_ | _1441_;
	assign _1824_ = (_1730_ ? _1822_ : _1823_);
	assign _1825_ = (_1766_ ? _1821_ : _1824_);
	assign _1826_ = (_1768_ ? _1820_ : _1825_);
	assign _1827_ = (_1774_ ? _1817_ : _1826_);
	assign _1828_ = ~(_1763_ | _1448_);
	assign _1829_ = ~_1828_;
	assign _1830_ = (_1730_ ? _1823_ : _1829_);
	assign _1831_ = (_1766_ ? _1830_ : _1829_);
	assign _1832_ = _1763_ | _1454_;
	assign _1833_ = (_1766_ ? _1832_ : _1818_);
	assign _1834_ = (_1768_ ? _1831_ : _1833_);
	assign _1835_ = _1818_ | ~_1730_;
	assign _1836_ = (_1766_ ? _1818_ : _1835_);
	assign _1837_ = (_1730_ ? _1792_ : _1829_);
	assign _1838_ = (_1766_ ? _1792_ : _1837_);
	assign _1839_ = (_1768_ ? _1836_ : _1838_);
	assign _1840_ = (_1774_ ? _1834_ : _1839_);
	assign _1841_ = (_1785_ ? _1827_ : _1840_);
	assign _1842_ = (_1806_ ? _1803_ : _1841_);
	assign _1843_ = ~(_1842_ | _1729_);
	assign _1844_ = _1716_ & ~_1728_;
	assign _1845_ = ~(_1844_ | _1748_);
	assign _1846_ = _1845_ ^ _1749_;
	assign _1847_ = (_1766_ ? _1828_ : _1775_);
	assign _1848_ = ~(_1763_ | _1474_);
	assign _1849_ = (_1766_ ? _1775_ : _1848_);
	assign _1850_ = (_1768_ ? _1847_ : _1849_);
	assign _1851_ = ~(_1763_ | _1478_);
	assign _1852_ = (_1730_ ? _1848_ : _1851_);
	assign _1853_ = (_1766_ ? _1852_ : _1851_);
	assign _1854_ = _1484_ & ~_1763_;
	assign _1855_ = ~(_1763_ | _1489_);
	assign _1856_ = _1855_ & ~_1730_;
	assign _1857_ = (_1766_ ? _1854_ : _1856_);
	assign _1858_ = (_1768_ ? _1853_ : _1857_);
	assign _1859_ = (_1774_ ? _1850_ : _1858_);
	assign _1860_ = ~(_1763_ | _1496_);
	assign _1861_ = (_1766_ ? _1855_ : _1860_);
	assign _1862_ = ~(_1763_ | _1503_);
	assign _1863_ = (_1730_ ? _1860_ : _1862_);
	assign _1864_ = (_1766_ ? _1863_ : _1862_);
	assign _1865_ = (_1768_ ? _1861_ : _1864_);
	assign _1866_ = ~(_1763_ | _1510_);
	assign _1867_ = ~(_1763_ | _1513_);
	assign _1868_ = (_1730_ ? _1866_ : _1867_);
	assign _1869_ = (_1766_ ? _1866_ : _1868_);
	assign _1870_ = (_1768_ ? _1862_ : _1869_);
	assign _1871_ = (_1774_ ? _1865_ : _1870_);
	assign _1872_ = (_1785_ ? _1859_ : _1871_);
	assign _1873_ = ~_1730_;
	assign _1874_ = _1867_ & ~_1873_;
	assign _1875_ = ~(_1763_ | _1524_);
	assign _1876_ = (_1766_ ? _1874_ : _1875_);
	assign _1877_ = (_1730_ ? _1875_ : _1777_);
	assign _1878_ = (_1766_ ? _1877_ : _1777_);
	assign _1879_ = (_1768_ ? _1876_ : _1878_);
	assign _1880_ = ~(_1763_ | _1533_);
	assign _1881_ = (_1766_ ? _1777_ : _1880_);
	assign _1882_ = ~_1539_;
	assign _1883_ = _1882_ & ~_1763_;
	assign _1884_ = ~_1542_;
	assign _1885_ = _1884_ & ~_1763_;
	assign _1886_ = (_1730_ ? _1883_ : _1885_);
	assign _1887_ = ~(_1763_ | _1547_);
	assign _1888_ = (_1730_ ? _1885_ : _1887_);
	assign _1889_ = (_1766_ ? _1886_ : _1888_);
	assign _1890_ = (_1768_ ? _1881_ : _1889_);
	assign _1891_ = (_1774_ ? _1879_ : _1890_);
	assign _1892_ = _1554_ & ~_1763_;
	assign _1893_ = (_1766_ ? _1887_ : _1892_);
	assign _1894_ = ~(_1763_ | _1558_);
	assign _1895_ = _1894_ & ~_1730_;
	assign _1896_ = (_1766_ ? _1895_ : _1894_);
	assign _1897_ = (_1768_ ? _1893_ : _1896_);
	assign _1898_ = ~(_1763_ | _1565_);
	assign _1899_ = (_1730_ ? _1777_ : _1786_);
	assign _1900_ = (_1766_ ? _1898_ : _1899_);
	assign _1901_ = (_1730_ ? _1786_ : _1809_);
	assign _1902_ = (_1766_ ? _1901_ : _1809_);
	assign _1903_ = (_1768_ ? _1900_ : _1902_);
	assign _1904_ = (_1774_ ? _1897_ : _1903_);
	assign _1905_ = (_1785_ ? _1891_ : _1904_);
	assign _1906_ = (_1806_ ? _1872_ : _1905_);
	assign _1907_ = ~(_1763_ | _1576_);
	assign _1908_ = (_1766_ ? _1775_ : _1907_);
	assign _1909_ = ~(_1763_ | _1580_);
	assign _1910_ = (_1730_ ? _1907_ : _1909_);
	assign _1911_ = _1909_ & ~_1873_;
	assign _1912_ = (_1766_ ? _1910_ : _1911_);
	assign _1913_ = (_1768_ ? _1908_ : _1912_);
	assign _1914_ = ~(_1763_ | _1587_);
	assign _1915_ = (_1730_ ? _1914_ : _1786_);
	assign _1916_ = (_1766_ ? _1914_ : _1915_);
	assign _1917_ = ~(_1763_ | _1592_);
	assign _1918_ = (_1730_ ? _1786_ : _1917_);
	assign _1919_ = (_1766_ ? _1918_ : _1807_);
	assign _1920_ = (_1768_ ? _1916_ : _1919_);
	assign _1921_ = (_1774_ ? _1913_ : _1920_);
	assign _1922_ = (_1766_ ? _1799_ : _1828_);
	assign _1923_ = ~(_1763_ | _1600_);
	assign _1924_ = (_1730_ ? _1828_ : _1923_);
	assign _1925_ = (_1766_ ? _1924_ : _1923_);
	assign _1926_ = (_1768_ ? _1922_ : _1925_);
	assign _1927_ = ~(_1763_ | _1606_);
	assign _1928_ = ~(_1763_ | _1609_);
	assign _1929_ = _1927_ & ~_1730_;
	assign _1930_ = (_1766_ ? _1928_ : _1929_);
	assign _1931_ = (_1768_ ? _1930_ : _1927_);
	assign _1932_ = (_1774_ ? _1926_ : _1931_);
	assign _1933_ = (_1785_ ? _1921_ : _1932_);
	assign _1934_ = ~_1617_;
	assign _1935_ = _1934_ & ~_1763_;
	assign _1936_ = (_1766_ ? _1777_ : _1935_);
	assign _1937_ = (_1768_ ? _1777_ : _1936_);
	assign _1938_ = _1927_ & ~_1873_;
	assign _1939_ = (_1766_ ? _1927_ : _1938_);
	assign _1940_ = _1887_ & ~_1766_;
	assign _1941_ = (_1768_ ? _1939_ : _1940_);
	assign _1942_ = (_1774_ ? _1937_ : _1941_);
	assign _1943_ = ~(_1763_ | _1626_);
	assign _1944_ = (_1730_ ? _1887_ : _1943_);
	assign _1945_ = (_1730_ ? _1943_ : _1777_);
	assign _1946_ = (_1766_ ? _1944_ : _1945_);
	assign _1947_ = (_1766_ ? _1631_ : _1632_);
	assign _1948_ = ~(_1947_ | _1763_);
	assign _1949_ = (_1768_ ? _1946_ : _1948_);
	assign _1950_ = (_1730_ ? _1907_ : _1943_);
	assign _1951_ = (_1766_ ? _1907_ : _1950_);
	assign _1952_ = (_1766_ ? _1943_ : _1887_);
	assign _1953_ = (_1768_ ? _1951_ : _1952_);
	assign _1954_ = (_1774_ ? _1949_ : _1953_);
	assign _1955_ = (_1785_ ? _1942_ : _1954_);
	assign _1956_ = (_1806_ ? _1933_ : _1955_);
	assign _1957_ = (_1729_ ? _1906_ : _1956_);
	assign _1958_ = (_1846_ ? _1843_ : _1957_);
	assign _1959_ = _1758_ ^ _1757_;
	assign _1960_ = _1958_ & ~_1959_;
	assign _1961_ = \mchip.game2.vga_inst.haddr [0] | ~\mchip.game2.vga_inst.haddr [1];
	assign _1962_ = \mchip.game2.vga_inst.haddr [3] | ~\mchip.game2.vga_inst.haddr [2];
	assign _1963_ = ~(_1962_ | _1961_);
	assign _1964_ = ~(_1963_ & _1731_);
	assign _1965_ = _1964_ | _1648_;
	assign _1966_ = ~(_1962_ | _0241_);
	assign _1967_ = _3186_ & ~_1966_;
	assign _1968_ = _1731_ & ~_1967_;
	assign _1969_ = _1731_ & ~_1968_;
	assign _1970_ = _1647_ & ~_1969_;
	assign _1971_ = _1653_ & ~_1970_;
	assign _1972_ = _1965_ & ~_1971_;
	assign _1973_ = _0241_ | ~_3185_;
	assign _1974_ = _1649_ & ~_1973_;
	assign _1975_ = _1654_ & ~_1974_;
	assign _1976_ = _1647_ & ~_1975_;
	assign _1977_ = _1976_ | _0237_;
	assign _1978_ = _1972_ & ~_1977_;
	assign _1979_ = _3179_ & ~_0242_;
	assign _1980_ = _0248_ & ~_1979_;
	assign _1981_ = \mchip.game2.vga_inst.haddr [4] & ~_1980_;
	assign _1982_ = _1981_ ^ \mchip.game2.vga_inst.haddr [5];
	assign _1983_ = ~_1982_;
	assign _1984_ = \mchip.game2.score_inst.score_saved[1] [2] & \mchip.game2.score_inst.score_saved[1] [3];
	assign _1985_ = ~(\mchip.game2.score_inst.score_saved[1] [0] ^ \mchip.game2.score_inst.score_saved[1] [3]);
	assign _1986_ = _1985_ ^ _1984_;
	assign _1987_ = ~(\mchip.game2.score_inst.score_saved[1] [2] & \mchip.game2.score_inst.score_saved[1] [1]);
	assign _1988_ = ~(\mchip.game2.score_inst.score_saved[1] [2] ^ \mchip.game2.score_inst.score_saved[1] [3]);
	assign _1989_ = _1988_ | _1987_;
	assign _1990_ = _1988_ ^ _1987_;
	assign _1991_ = ~(\mchip.game2.score_inst.score_saved[1] [1] & \mchip.game2.score_inst.score_saved[1] [0]);
	assign _1992_ = ~(\mchip.game2.score_inst.score_saved[1] [2] ^ \mchip.game2.score_inst.score_saved[1] [1]);
	assign _1993_ = _1992_ | _1991_;
	assign _1994_ = _1990_ & ~_1993_;
	assign _1995_ = _1989_ & ~_1994_;
	assign _1996_ = _1995_ | _1986_;
	assign _1997_ = _1984_ & ~_1985_;
	assign _1998_ = ~(\mchip.game2.score_inst.score_saved[1] [0] & \mchip.game2.score_inst.score_saved[1] [3]);
	assign _1999_ = _1998_ ^ \mchip.game2.score_inst.score_saved[1] [1];
	assign _2000_ = _1999_ ^ _1997_;
	assign _2001_ = _2000_ ^ _1996_;
	assign _2002_ = _2001_ & ~_1983_;
	assign _2003_ = _2001_ ^ _1983_;
	assign _2004_ = _1980_ ^ \mchip.game2.vga_inst.haddr [4];
	assign _2005_ = _1995_ ^ _1986_;
	assign _2006_ = _2004_ | ~_2005_;
	assign _2007_ = ~(_2006_ | _2003_);
	assign _2008_ = _2007_ | _2002_;
	assign _2009_ = _2005_ ^ _2004_;
	assign _2010_ = _2009_ | _2003_;
	assign _2011_ = _1238_ ^ _0662_;
	assign _2012_ = ~(_1993_ ^ _1990_);
	assign _2013_ = ~(_2012_ & _2011_);
	assign _2014_ = ~(_2012_ ^ _2011_);
	assign _2015_ = _3179_ ^ _1232_;
	assign _2016_ = _1992_ ^ _1991_;
	assign _2017_ = ~(_2016_ & _2015_);
	assign _2018_ = ~(_2017_ | _2014_);
	assign _2019_ = _2013_ & ~_2018_;
	assign _2020_ = _2016_ ^ _2015_;
	assign _2021_ = _2020_ & ~_2014_;
	assign _2022_ = \mchip.game2.score_inst.score_saved[1] [1] ^ \mchip.game2.score_inst.score_saved[1] [0];
	assign _2023_ = _3625_[1] | ~_2022_;
	assign _2024_ = \mchip.game2.score_inst.score_saved[1] [0] & ~\mchip.game2.vga_inst.haddr [0];
	assign _2025_ = ~(_2022_ ^ _3625_[1]);
	assign _2026_ = _2025_ & _2024_;
	assign _2027_ = _2023_ & ~_2026_;
	assign _2028_ = _2021_ & ~_2027_;
	assign _2029_ = _2019_ & ~_2028_;
	assign _2030_ = ~(_2029_ | _2010_);
	assign _2031_ = _2030_ | _2008_;
	assign _2032_ = ~(_1980_ | _1717_);
	assign _2033_ = _2032_ ^ \mchip.game2.vga_inst.haddr [6];
	assign _2034_ = _1997_ & ~_1999_;
	assign _2035_ = _2000_ | _1986_;
	assign _2036_ = ~(_2035_ | _1995_);
	assign _2037_ = _2036_ | _2034_;
	assign _2038_ = \mchip.game2.score_inst.score_saved[1] [1] & ~_1998_;
	assign _2039_ = ~(_2038_ ^ \mchip.game2.score_inst.score_saved[1] [2]);
	assign _2040_ = _2039_ ^ _2037_;
	assign _2041_ = _2040_ ^ _2033_;
	assign _2042_ = ~(_2041_ ^ _2031_);
	assign _2043_ = ~(\mchip.game2.score_inst.score_saved[1] [0] ^ \mchip.game2.vga_inst.haddr [0]);
	assign _2044_ = ~(_1980_ | _1732_);
	assign _2045_ = _2044_ ^ \mchip.game2.vga_inst.haddr [8];
	assign _2046_ = ~\mchip.game2.score_inst.score_saved[1] [3];
	assign _2047_ = ~(_2038_ & \mchip.game2.score_inst.score_saved[1] [2]);
	assign _2048_ = _2047_ | _2046_;
	assign _2049_ = _2039_ | _2046_;
	assign _2050_ = _2034_ & ~_2049_;
	assign _2051_ = _2048_ & ~_2050_;
	assign _2052_ = _2049_ | _2035_;
	assign _2053_ = ~(_2052_ | _1995_);
	assign _2054_ = _2051_ & ~_2053_;
	assign _2055_ = _2045_ & ~_2054_;
	assign _2056_ = ~(_2032_ & \mchip.game2.vga_inst.haddr [6]);
	assign _2057_ = _2056_ ^ \mchip.game2.vga_inst.haddr [7];
	assign _2058_ = _2037_ & ~_2039_;
	assign _2059_ = _2047_ & ~_2058_;
	assign _2060_ = _2059_ ^ _2046_;
	assign _2061_ = _2060_ & ~_2057_;
	assign _2062_ = _2033_ & ~_2040_;
	assign _2063_ = _2060_ ^ _2057_;
	assign _2064_ = _2062_ & ~_2063_;
	assign _2065_ = _2064_ | _2061_;
	assign _2066_ = _2063_ | _2041_;
	assign _2067_ = _2008_ & ~_2066_;
	assign _2068_ = _2067_ | _2065_;
	assign _2069_ = _2066_ | _2010_;
	assign _2070_ = ~(_2069_ | _2029_);
	assign _2071_ = _2070_ | _2068_;
	assign _2072_ = ~(_2054_ ^ _2045_);
	assign _2073_ = _2072_ & _2071_;
	assign _2074_ = _2073_ | _2055_;
	assign _2075_ = _2044_ & ~_1269_;
	assign _2076_ = _2075_ ^ _1307_;
	assign _2077_ = _2076_ ^ _2074_;
	assign _2078_ = _2077_ | _1323_;
	assign _2079_ = _2078_ | _2043_;
	assign _2080_ = _2025_ ^ _2024_;
	assign _2081_ = _2080_ | _2079_;
	assign _2082_ = ~(_2027_ ^ _2020_);
	assign _2083_ = _2077_ | _1335_;
	assign _2084_ = (_2080_ ? _2078_ : _2083_);
	assign _2085_ = (_2082_ ? _2081_ : _2084_);
	assign _2086_ = _2020_ & ~_2027_;
	assign _2087_ = _2017_ & ~_2086_;
	assign _2088_ = _2087_ ^ _2014_;
	assign _2089_ = _2077_ | _1349_;
	assign _2090_ = _2077_ | _1352_;
	assign _2091_ = _2077_ | _1358_;
	assign _2092_ = (_2043_ ? _2090_ : _2091_);
	assign _2093_ = (_2043_ ? _2091_ : _2089_);
	assign _2094_ = (_2080_ ? _2092_ : _2093_);
	assign _2095_ = (_2082_ ? _2094_ : _2089_);
	assign _2096_ = (_2088_ ? _2085_ : _2095_);
	assign _2097_ = _2029_ ^ _2009_;
	assign _2098_ = _2077_ | _1370_;
	assign _2099_ = _2077_ | _1376_;
	assign _2100_ = (_2043_ ? _2098_ : _2099_);
	assign _2101_ = (_2080_ ? _2098_ : _2100_);
	assign _2102_ = _2099_ | ~_2043_;
	assign _2103_ = _2077_ | _1382_;
	assign _2104_ = (_2080_ ? _2102_ : _2103_);
	assign _2105_ = (_2082_ ? _2101_ : _2104_);
	assign _2106_ = _2077_ | _1388_;
	assign _2107_ = (_2043_ ? _2103_ : _2106_);
	assign _2108_ = (_2043_ ? _2106_ : _2090_);
	assign _2109_ = (_2080_ ? _2107_ : _2108_);
	assign _2110_ = ~(_2077_ | _1397_);
	assign _2111_ = ~_2110_;
	assign _2112_ = (_2082_ ? _2109_ : _2111_);
	assign _2113_ = (_2088_ ? _2105_ : _2112_);
	assign _2114_ = (_2097_ ? _2096_ : _2113_);
	assign _2115_ = ~(_2029_ | _2009_);
	assign _2116_ = _2006_ & ~_2115_;
	assign _2117_ = _2116_ ^ _2003_;
	assign _2118_ = _2077_ | _1410_;
	assign _2119_ = _2077_ | _1416_;
	assign _2120_ = (_2043_ ? _2118_ : _2119_);
	assign _2121_ = (_2043_ ? _2119_ : _2098_);
	assign _2122_ = (_2080_ ? _2120_ : _2121_);
	assign _2123_ = (_2043_ ? _2098_ : _2090_);
	assign _2124_ = _2077_ | _1424_;
	assign _2125_ = (_2080_ ? _2123_ : _2124_);
	assign _2126_ = (_2082_ ? _2122_ : _2125_);
	assign _2127_ = _2077_ | _1429_;
	assign _2128_ = _2127_ | _2043_;
	assign _2129_ = (_2080_ ? _2128_ : _2127_);
	assign _2130_ = _2077_ | _1433_;
	assign _2131_ = _2077_ | _1437_;
	assign _2132_ = _2077_ | _1441_;
	assign _2133_ = (_2043_ ? _2131_ : _2132_);
	assign _2134_ = (_2080_ ? _2130_ : _2133_);
	assign _2135_ = (_2082_ ? _2129_ : _2134_);
	assign _2136_ = (_2088_ ? _2126_ : _2135_);
	assign _2137_ = _2077_ | _1448_;
	assign _2138_ = (_2043_ ? _2132_ : _2137_);
	assign _2139_ = (_2080_ ? _2138_ : _2137_);
	assign _2140_ = _2077_ | _1454_;
	assign _2141_ = (_2080_ ? _2140_ : _2127_);
	assign _2142_ = (_2082_ ? _2139_ : _2141_);
	assign _2143_ = _2127_ | ~_2043_;
	assign _2144_ = (_2080_ ? _2127_ : _2143_);
	assign _2145_ = (_2043_ ? _2103_ : _2137_);
	assign _2146_ = (_2080_ ? _2103_ : _2145_);
	assign _2147_ = (_2082_ ? _2144_ : _2146_);
	assign _2148_ = (_2088_ ? _2142_ : _2147_);
	assign _2149_ = (_2097_ ? _2136_ : _2148_);
	assign _2150_ = (_2117_ ? _2114_ : _2149_);
	assign _2151_ = ~(_2150_ | _2042_);
	assign _2152_ = _2031_ & ~_2041_;
	assign _2153_ = ~(_2152_ | _2062_);
	assign _2154_ = _2153_ ^ _2063_;
	assign _2155_ = ~_2089_;
	assign _2156_ = ~(_2077_ | _1448_);
	assign _2157_ = (_2080_ ? _2156_ : _2155_);
	assign _2158_ = ~(_2077_ | _1474_);
	assign _2159_ = (_2080_ ? _2155_ : _2158_);
	assign _2160_ = (_2082_ ? _2157_ : _2159_);
	assign _2161_ = ~(_2077_ | _1478_);
	assign _2162_ = (_2043_ ? _2158_ : _2161_);
	assign _2163_ = (_2080_ ? _2162_ : _2161_);
	assign _2164_ = _1484_ & ~_2077_;
	assign _2165_ = ~(_2077_ | _1489_);
	assign _2166_ = _2165_ & ~_2043_;
	assign _2167_ = (_2080_ ? _2164_ : _2166_);
	assign _2168_ = (_2082_ ? _2163_ : _2167_);
	assign _2169_ = (_2088_ ? _2160_ : _2168_);
	assign _2170_ = ~(_2077_ | _1496_);
	assign _2171_ = (_2080_ ? _2165_ : _2170_);
	assign _2172_ = ~(_2077_ | _1503_);
	assign _2173_ = (_2043_ ? _2170_ : _2172_);
	assign _2174_ = (_2080_ ? _2173_ : _2172_);
	assign _2175_ = (_2082_ ? _2171_ : _2174_);
	assign _2176_ = ~(_2077_ | _1510_);
	assign _2177_ = ~(_2077_ | _1513_);
	assign _2178_ = (_2043_ ? _2176_ : _2177_);
	assign _2179_ = (_2080_ ? _2176_ : _2178_);
	assign _2180_ = (_2082_ ? _2172_ : _2179_);
	assign _2181_ = (_2088_ ? _2175_ : _2180_);
	assign _2182_ = (_2097_ ? _2169_ : _2181_);
	assign _2183_ = ~_2043_;
	assign _2184_ = _2177_ & ~_2183_;
	assign _2185_ = ~(_2077_ | _1524_);
	assign _2186_ = (_2080_ ? _2184_ : _2185_);
	assign _2187_ = ~(_2077_ | _1352_);
	assign _2188_ = (_2043_ ? _2185_ : _2187_);
	assign _2189_ = (_2080_ ? _2188_ : _2187_);
	assign _2190_ = (_2082_ ? _2186_ : _2189_);
	assign _2191_ = ~(_2077_ | _1533_);
	assign _2192_ = (_2080_ ? _2187_ : _2191_);
	assign _2193_ = _1882_ & ~_2077_;
	assign _2194_ = _1884_ & ~_2077_;
	assign _2195_ = (_2043_ ? _2193_ : _2194_);
	assign _2196_ = ~(_2077_ | _1547_);
	assign _2197_ = (_2043_ ? _2194_ : _2196_);
	assign _2198_ = (_2080_ ? _2195_ : _2197_);
	assign _2199_ = (_2082_ ? _2192_ : _2198_);
	assign _2200_ = (_2088_ ? _2190_ : _2199_);
	assign _2201_ = _1554_ & ~_2077_;
	assign _2202_ = (_2080_ ? _2196_ : _2201_);
	assign _2203_ = ~(_2077_ | _1558_);
	assign _2204_ = _2203_ & ~_2043_;
	assign _2205_ = (_2080_ ? _2204_ : _2203_);
	assign _2206_ = (_2082_ ? _2202_ : _2205_);
	assign _2207_ = ~(_2077_ | _1565_);
	assign _2208_ = ~(_2077_ | _1370_);
	assign _2209_ = (_2043_ ? _2187_ : _2208_);
	assign _2210_ = (_2080_ ? _2207_ : _2209_);
	assign _2211_ = ~(_2077_ | _1416_);
	assign _2212_ = (_2043_ ? _2208_ : _2211_);
	assign _2213_ = (_2080_ ? _2212_ : _2211_);
	assign _2214_ = (_2082_ ? _2210_ : _2213_);
	assign _2215_ = (_2088_ ? _2206_ : _2214_);
	assign _2216_ = (_2097_ ? _2200_ : _2215_);
	assign _2217_ = (_2117_ ? _2182_ : _2216_);
	assign _2218_ = ~(_2077_ | _1576_);
	assign _2219_ = (_2080_ ? _2155_ : _2218_);
	assign _2220_ = ~(_2077_ | _1580_);
	assign _2221_ = (_2043_ ? _2218_ : _2220_);
	assign _2222_ = _2220_ & ~_2183_;
	assign _2223_ = (_2080_ ? _2221_ : _2222_);
	assign _2224_ = (_2082_ ? _2219_ : _2223_);
	assign _2225_ = ~(_2077_ | _1587_);
	assign _2226_ = (_2043_ ? _2225_ : _2208_);
	assign _2227_ = (_2080_ ? _2225_ : _2226_);
	assign _2228_ = ~_2118_;
	assign _2229_ = ~(_2077_ | _1592_);
	assign _2230_ = (_2043_ ? _2208_ : _2229_);
	assign _2231_ = (_2080_ ? _2230_ : _2228_);
	assign _2232_ = (_2082_ ? _2227_ : _2231_);
	assign _2233_ = (_2088_ ? _2224_ : _2232_);
	assign _2234_ = (_2080_ ? _2110_ : _2156_);
	assign _2235_ = ~(_2077_ | _1600_);
	assign _2236_ = (_2043_ ? _2156_ : _2235_);
	assign _2237_ = (_2080_ ? _2236_ : _2235_);
	assign _2238_ = (_2082_ ? _2234_ : _2237_);
	assign _2239_ = _2077_ | _1606_;
	assign _2240_ = ~_2239_;
	assign _2241_ = ~(_2077_ | _1609_);
	assign _2242_ = _2183_ & ~_2239_;
	assign _2243_ = (_2080_ ? _2241_ : _2242_);
	assign _2244_ = (_2082_ ? _2243_ : _2240_);
	assign _2245_ = (_2088_ ? _2238_ : _2244_);
	assign _2246_ = (_2097_ ? _2233_ : _2245_);
	assign _2247_ = _1934_ & ~_2077_;
	assign _2248_ = (_2080_ ? _2187_ : _2247_);
	assign _2249_ = (_2082_ ? _2187_ : _2248_);
	assign _2250_ = _2043_ & ~_2239_;
	assign _2251_ = (_2080_ ? _2240_ : _2250_);
	assign _2252_ = _2196_ & ~_2080_;
	assign _2253_ = (_2082_ ? _2251_ : _2252_);
	assign _2254_ = (_2088_ ? _2249_ : _2253_);
	assign _2255_ = ~(_2077_ | _1626_);
	assign _2256_ = (_2043_ ? _2196_ : _2255_);
	assign _2257_ = (_2043_ ? _2255_ : _2187_);
	assign _2258_ = (_2080_ ? _2256_ : _2257_);
	assign _2259_ = (_2080_ ? _1631_ : _1632_);
	assign _2260_ = ~(_2259_ | _2077_);
	assign _2261_ = (_2082_ ? _2258_ : _2260_);
	assign _2262_ = (_2043_ ? _2218_ : _2255_);
	assign _2263_ = (_2080_ ? _2218_ : _2262_);
	assign _2264_ = (_2080_ ? _2255_ : _2196_);
	assign _2265_ = (_2082_ ? _2263_ : _2264_);
	assign _2266_ = (_2088_ ? _2261_ : _2265_);
	assign _2267_ = (_2097_ ? _2254_ : _2266_);
	assign _2268_ = (_2117_ ? _2246_ : _2267_);
	assign _2269_ = (_2042_ ? _2217_ : _2268_);
	assign _2270_ = (_2154_ ? _2151_ : _2269_);
	assign _2271_ = _2072_ ^ _2071_;
	assign _2272_ = _2270_ & ~_2271_;
	assign _2273_ = \mchip.game2.vga_inst.haddr [9] & ~\mchip.game2.vga_inst.haddr [8];
	assign _2274_ = ~(_2273_ & _3182_);
	assign _2275_ = _0248_ & _0239_;
	assign _2276_ = _2275_ | _2274_;
	assign _2277_ = _2273_ & ~_3182_;
	assign _2278_ = _2277_ | _3181_;
	assign _2279_ = _2276_ & ~_2278_;
	assign _2280_ = ~(_0242_ | _3179_);
	assign _2281_ = \mchip.game2.vga_inst.haddr [3] & ~_2280_;
	assign _2282_ = _1731_ & ~_2281_;
	assign _2283_ = _1731_ & ~_2282_;
	assign _2284_ = _1647_ & ~_2283_;
	assign _2285_ = _2284_ | _0237_;
	assign _2286_ = _2279_ & ~_2285_;
	assign _2287_ = _3227_ & _3174_;
	assign _2288_ = \mchip.game2.vga_inst.haddr [4] | ~\mchip.game2.vga_inst.haddr [3];
	assign _2289_ = _0663_ & ~_2288_;
	assign _2290_ = _1199_ & ~_2289_;
	assign _2291_ = _2287_ & ~_2290_;
	assign _2292_ = _2287_ & ~_2291_;
	assign _2293_ = \mchip.game2.vga_inst.haddr [9] & ~_2292_;
	assign _2294_ = ~(_1961_ | _0248_);
	assign _2295_ = ~(_2294_ & _0257_);
	assign _2296_ = _2273_ & ~_2295_;
	assign _2297_ = _2293_ & ~_2296_;
	assign _2298_ = _3227_ & ~\mchip.game2.vga_inst.haddr [6];
	assign _2299_ = \mchip.game2.vga_inst.haddr [6] | ~\mchip.game2.vga_inst.haddr [5];
	assign _2300_ = _3227_ & ~_2299_;
	assign _2301_ = \mchip.game2.vga_inst.haddr [3] | \mchip.game2.vga_inst.haddr [4];
	assign _2302_ = _0724_ & ~_2301_;
	assign _2303_ = _2300_ & ~_2302_;
	assign _2304_ = _2298_ & ~_2303_;
	assign _2305_ = \mchip.game2.vga_inst.haddr [9] & ~_2304_;
	assign _2306_ = _2297_ & ~_2305_;
	assign _2307_ = _0253_ | ~_0239_;
	assign _2308_ = _1256_ & ~_2307_;
	assign _2309_ = _2308_ ^ \mchip.game2.vga_inst.haddr [7];
	assign _2310_ = \mchip.game2.score_inst.score_saved[0] [0] & \mchip.game2.score_inst.score_saved[0] [3];
	assign _2311_ = ~(_2310_ & \mchip.game2.score_inst.score_saved[0] [1]);
	assign _2312_ = _2310_ ^ \mchip.game2.score_inst.score_saved[0] [1];
	assign _2313_ = ~(\mchip.game2.score_inst.score_saved[0] [1] & \mchip.game2.score_inst.score_saved[0] [2]);
	assign _2314_ = ~\mchip.game2.score_inst.score_saved[0] [3];
	assign _2315_ = \mchip.game2.score_inst.score_saved[0] [2] & ~\mchip.game2.score_inst.score_saved[0] [1];
	assign _2316_ = _2315_ & ~_2314_;
	assign _2317_ = _2316_ | ~_2313_;
	assign _2318_ = \mchip.game2.score_inst.score_saved[0] [0] ^ \mchip.game2.score_inst.score_saved[0] [3];
	assign _2319_ = ~(_2318_ & _2317_);
	assign _2320_ = _2312_ & ~_2319_;
	assign _2321_ = _2311_ & ~_2320_;
	assign _2322_ = _2318_ ^ _2317_;
	assign _2323_ = _2322_ & _2312_;
	assign _2324_ = \mchip.game2.score_inst.score_saved[0] [1] & \mchip.game2.score_inst.score_saved[0] [0];
	assign _2325_ = ~(\mchip.game2.score_inst.score_saved[0] [1] ^ \mchip.game2.score_inst.score_saved[0] [2]);
	assign _2326_ = _2324_ & ~_2325_;
	assign _2327_ = _2315_ ^ _2314_;
	assign _2328_ = _2326_ & ~_2327_;
	assign _2329_ = ~_2328_;
	assign _2330_ = _2323_ & ~_2329_;
	assign _2331_ = _2321_ & ~_2330_;
	assign _2332_ = \mchip.game2.score_inst.score_saved[0] [2] & ~_2331_;
	assign _2333_ = _2332_ ^ \mchip.game2.score_inst.score_saved[0] [3];
	assign _2334_ = _2333_ & _2309_;
	assign _2335_ = _2333_ ^ _2309_;
	assign _2336_ = _2307_ ^ \mchip.game2.vga_inst.haddr [6];
	assign _2337_ = ~(_2331_ ^ \mchip.game2.score_inst.score_saved[0] [2]);
	assign _2338_ = _2336_ | ~_2337_;
	assign _2339_ = _2335_ & ~_2338_;
	assign _2340_ = _2339_ | _2334_;
	assign _2341_ = _2337_ ^ _2336_;
	assign _2342_ = _2335_ & ~_2341_;
	assign _2343_ = _1199_ & ~_0253_;
	assign _2344_ = _2343_ ^ \mchip.game2.vga_inst.haddr [5];
	assign _2345_ = _2322_ & ~_2329_;
	assign _2346_ = _2319_ & ~_2345_;
	assign _2347_ = ~(_2346_ ^ _2312_);
	assign _2348_ = ~(_2347_ & _2344_);
	assign _2349_ = _2347_ ^ _2344_;
	assign _2350_ = _2328_ ^ _2322_;
	assign _2351_ = _3625_[4] | ~_2350_;
	assign _2352_ = _2349_ & ~_2351_;
	assign _2353_ = _2348_ & ~_2352_;
	assign _2354_ = _2342_ & ~_2353_;
	assign _2355_ = _2354_ | _2340_;
	assign _2356_ = _2350_ ^ _3625_[4];
	assign _2357_ = _2356_ | ~_2349_;
	assign _2358_ = _2342_ & ~_2357_;
	assign _2359_ = _0241_ & ~_1232_;
	assign _3625_[3] = _2359_ ^ \mchip.game2.vga_inst.haddr [3];
	assign _2360_ = ~(_2327_ ^ _2326_);
	assign _2361_ = ~(_2360_ & _3625_[3]);
	assign _2362_ = ~(_2360_ ^ _3625_[3]);
	assign _3625_[2] = ~(_2359_ | _1695_);
	assign _2363_ = ~(_2325_ ^ _2324_);
	assign _2364_ = ~(_2363_ & _3625_[2]);
	assign _2365_ = ~(_2364_ | _2362_);
	assign _2366_ = _2361_ & ~_2365_;
	assign _2367_ = _2363_ ^ _3625_[2];
	assign _2368_ = _2367_ & ~_2362_;
	assign _2369_ = \mchip.game2.score_inst.score_saved[0] [1] ^ \mchip.game2.score_inst.score_saved[0] [0];
	assign _2370_ = ~(_2369_ & _3625_[1]);
	assign _2371_ = \mchip.game2.score_inst.score_saved[0] [0] & ~\mchip.game2.vga_inst.haddr [0];
	assign _2372_ = _2369_ ^ _3625_[1];
	assign _2373_ = _2372_ & _2371_;
	assign _2374_ = _2370_ & ~_2373_;
	assign _2375_ = _2368_ & ~_2374_;
	assign _2376_ = _2366_ & ~_2375_;
	assign _2377_ = _2358_ & ~_2376_;
	assign _2378_ = _2377_ | _2355_;
	assign _2379_ = _0253_ & _0257_;
	assign _2380_ = _0257_ & ~_2379_;
	assign _2381_ = _2380_ ^ \mchip.game2.vga_inst.haddr [8];
	assign _2382_ = ~(\mchip.game2.score_inst.score_saved[0] [2] & \mchip.game2.score_inst.score_saved[0] [3]);
	assign _2383_ = _2382_ | _2321_;
	assign _2384_ = _2382_ | ~_2323_;
	assign _2385_ = _2328_ & ~_2384_;
	assign _2386_ = _2383_ & ~_2385_;
	assign _2387_ = ~(_2386_ ^ _2381_);
	assign _2388_ = _2387_ ^ _2378_;
	assign _2389_ = _2381_ & ~_2386_;
	assign _2390_ = _2387_ & _2378_;
	assign _2391_ = _2390_ | _2389_;
	assign _2392_ = _2380_ & ~\mchip.game2.vga_inst.haddr [8];
	assign _2393_ = _2392_ ^ _1307_;
	assign _2394_ = _2393_ ^ _2391_;
	assign _2395_ = _2394_ | _1323_;
	assign _2396_ = ~(\mchip.game2.score_inst.score_saved[0] [0] ^ \mchip.game2.vga_inst.haddr [0]);
	assign _2397_ = _2396_ | _2395_;
	assign _2398_ = _2372_ ^ _2371_;
	assign _2399_ = _2398_ | _2397_;
	assign _2400_ = ~(_2374_ ^ _2367_);
	assign _2401_ = _2394_ | _1335_;
	assign _2402_ = (_2398_ ? _2395_ : _2401_);
	assign _2403_ = (_2400_ ? _2399_ : _2402_);
	assign _2404_ = _2367_ & ~_2374_;
	assign _2405_ = _2364_ & ~_2404_;
	assign _2406_ = _2405_ ^ _2362_;
	assign _2407_ = _2394_ | _1352_;
	assign _2408_ = _2394_ | _1358_;
	assign _2409_ = (_2396_ ? _2407_ : _2408_);
	assign _2410_ = _2394_ | _1349_;
	assign _2411_ = (_2396_ ? _2408_ : _2410_);
	assign _2412_ = (_2398_ ? _2409_ : _2411_);
	assign _2413_ = (_2400_ ? _2412_ : _2410_);
	assign _2414_ = (_2406_ ? _2403_ : _2413_);
	assign _2415_ = _2376_ ^ _2356_;
	assign _2416_ = _2394_ | _1370_;
	assign _2417_ = _2394_ | _1376_;
	assign _2418_ = (_2396_ ? _2416_ : _2417_);
	assign _2419_ = (_2398_ ? _2416_ : _2418_);
	assign _2420_ = _2417_ | ~_2396_;
	assign _2421_ = _2394_ | _1382_;
	assign _2422_ = (_2398_ ? _2420_ : _2421_);
	assign _2423_ = (_2400_ ? _2419_ : _2422_);
	assign _2424_ = _2394_ | _1388_;
	assign _2425_ = (_2396_ ? _2421_ : _2424_);
	assign _2426_ = (_2396_ ? _2424_ : _2407_);
	assign _2427_ = (_2398_ ? _2425_ : _2426_);
	assign _2428_ = _2394_ | _1397_;
	assign _2429_ = (_2400_ ? _2427_ : _2428_);
	assign _2430_ = (_2406_ ? _2423_ : _2429_);
	assign _2431_ = (_2415_ ? _2414_ : _2430_);
	assign _2432_ = ~(_2376_ | _2356_);
	assign _2433_ = _2432_ | ~_2351_;
	assign _2434_ = _2433_ ^ _2349_;
	assign _2435_ = _2394_ | _1410_;
	assign _2436_ = _2394_ | _1416_;
	assign _2437_ = (_2396_ ? _2435_ : _2436_);
	assign _2438_ = (_2396_ ? _2436_ : _2416_);
	assign _2439_ = (_2398_ ? _2437_ : _2438_);
	assign _2440_ = (_2396_ ? _2416_ : _2407_);
	assign _2441_ = _2394_ | _1424_;
	assign _2442_ = (_2398_ ? _2440_ : _2441_);
	assign _2443_ = (_2400_ ? _2439_ : _2442_);
	assign _2444_ = _2394_ | _1429_;
	assign _2445_ = _2444_ | _2396_;
	assign _2446_ = (_2398_ ? _2445_ : _2444_);
	assign _2447_ = _2394_ | _1433_;
	assign _2448_ = _2394_ | _1437_;
	assign _2449_ = _2394_ | _1441_;
	assign _2450_ = (_2396_ ? _2448_ : _2449_);
	assign _2451_ = (_2398_ ? _2447_ : _2450_);
	assign _2452_ = (_2400_ ? _2446_ : _2451_);
	assign _2453_ = (_2406_ ? _2443_ : _2452_);
	assign _2454_ = _2394_ | _1448_;
	assign _2455_ = (_2396_ ? _2449_ : _2454_);
	assign _2456_ = (_2398_ ? _2455_ : _2454_);
	assign _2457_ = _2394_ | _1454_;
	assign _2458_ = (_2398_ ? _2457_ : _2444_);
	assign _2459_ = (_2400_ ? _2456_ : _2458_);
	assign _2460_ = _2444_ | ~_2396_;
	assign _2461_ = (_2398_ ? _2444_ : _2460_);
	assign _2462_ = (_2396_ ? _2421_ : _2454_);
	assign _2463_ = (_2398_ ? _2421_ : _2462_);
	assign _2464_ = (_2400_ ? _2461_ : _2463_);
	assign _2465_ = (_2406_ ? _2459_ : _2464_);
	assign _2466_ = (_2415_ ? _2453_ : _2465_);
	assign _2467_ = (_2434_ ? _2431_ : _2466_);
	assign _2468_ = ~(_2376_ | _2357_);
	assign _2469_ = _2353_ & ~_2468_;
	assign _2470_ = _2469_ ^ _2341_;
	assign _2471_ = _2470_ | _2467_;
	assign _2472_ = ~(_2469_ | _2341_);
	assign _2473_ = _2472_ | ~_2338_;
	assign _2474_ = _2473_ ^ _2335_;
	assign _2475_ = (_2398_ ? _2454_ : _2410_);
	assign _2476_ = _2394_ | _1474_;
	assign _2477_ = (_2398_ ? _2410_ : _2476_);
	assign _2478_ = (_2400_ ? _2475_ : _2477_);
	assign _2479_ = _2394_ | _1478_;
	assign _2480_ = (_2396_ ? _2476_ : _2479_);
	assign _2481_ = (_2398_ ? _2480_ : _2479_);
	assign _2482_ = _2394_ | _1485_;
	assign _2483_ = _2394_ | _1489_;
	assign _2484_ = _2483_ | _2396_;
	assign _2485_ = (_2398_ ? _2482_ : _2484_);
	assign _2486_ = (_2400_ ? _2481_ : _2485_);
	assign _2487_ = (_2406_ ? _2478_ : _2486_);
	assign _2488_ = _2394_ | _1496_;
	assign _2489_ = (_2398_ ? _2483_ : _2488_);
	assign _2490_ = _2394_ | _1503_;
	assign _2491_ = (_2396_ ? _2488_ : _2490_);
	assign _2492_ = (_2398_ ? _2491_ : _2490_);
	assign _2493_ = (_2400_ ? _2489_ : _2492_);
	assign _2494_ = _2394_ | _1510_;
	assign _2495_ = _2394_ | _1513_;
	assign _2496_ = (_2396_ ? _2494_ : _2495_);
	assign _2497_ = (_2398_ ? _2494_ : _2496_);
	assign _2498_ = (_2400_ ? _2490_ : _2497_);
	assign _2499_ = (_2406_ ? _2493_ : _2498_);
	assign _2500_ = (_2415_ ? _2487_ : _2499_);
	assign _2501_ = _2495_ | ~_2396_;
	assign _2502_ = _2394_ | _1524_;
	assign _2503_ = (_2398_ ? _2501_ : _2502_);
	assign _2504_ = (_2396_ ? _2502_ : _2407_);
	assign _2505_ = (_2398_ ? _2504_ : _2407_);
	assign _2506_ = (_2400_ ? _2503_ : _2505_);
	assign _2507_ = _2394_ | _1533_;
	assign _2508_ = (_2398_ ? _2407_ : _2507_);
	assign _2509_ = _2394_ | _1539_;
	assign _2510_ = _2394_ | _1542_;
	assign _2511_ = (_2396_ ? _2509_ : _2510_);
	assign _2512_ = _2394_ | _1547_;
	assign _2513_ = (_2396_ ? _2510_ : _2512_);
	assign _2514_ = (_2398_ ? _2511_ : _2513_);
	assign _2515_ = (_2400_ ? _2508_ : _2514_);
	assign _2516_ = (_2406_ ? _2506_ : _2515_);
	assign _2517_ = _2394_ | _1555_;
	assign _2518_ = (_2398_ ? _2512_ : _2517_);
	assign _2519_ = _2394_ | _1558_;
	assign _2520_ = _2519_ | _2396_;
	assign _2521_ = (_2398_ ? _2520_ : _2519_);
	assign _2522_ = (_2400_ ? _2518_ : _2521_);
	assign _2523_ = _2394_ | _1565_;
	assign _2524_ = (_2396_ ? _2407_ : _2416_);
	assign _2525_ = (_2398_ ? _2523_ : _2524_);
	assign _2526_ = (_2396_ ? _2416_ : _2436_);
	assign _2527_ = (_2398_ ? _2526_ : _2436_);
	assign _2528_ = (_2400_ ? _2525_ : _2527_);
	assign _2529_ = (_2406_ ? _2522_ : _2528_);
	assign _2530_ = (_2415_ ? _2516_ : _2529_);
	assign _2531_ = (_2434_ ? _2500_ : _2530_);
	assign _2532_ = _2394_ | _1576_;
	assign _2533_ = (_2398_ ? _2410_ : _2532_);
	assign _2534_ = _2394_ | _1580_;
	assign _2535_ = (_2396_ ? _2532_ : _2534_);
	assign _2536_ = _2534_ | ~_2396_;
	assign _2537_ = (_2398_ ? _2535_ : _2536_);
	assign _2538_ = (_2400_ ? _2533_ : _2537_);
	assign _2539_ = _2394_ | _1587_;
	assign _2540_ = (_2396_ ? _2539_ : _2416_);
	assign _2541_ = (_2398_ ? _2539_ : _2540_);
	assign _2542_ = _2394_ | _1592_;
	assign _2543_ = (_2396_ ? _2416_ : _2542_);
	assign _2544_ = (_2398_ ? _2543_ : _2435_);
	assign _2545_ = (_2400_ ? _2541_ : _2544_);
	assign _2546_ = (_2406_ ? _2538_ : _2545_);
	assign _2547_ = (_2398_ ? _2428_ : _2454_);
	assign _2548_ = _2394_ | _1600_;
	assign _2549_ = (_2396_ ? _2454_ : _2548_);
	assign _2550_ = (_2398_ ? _2549_ : _2548_);
	assign _2551_ = (_2400_ ? _2547_ : _2550_);
	assign _2552_ = _2394_ | _1609_;
	assign _2553_ = _2394_ | _1606_;
	assign _2554_ = _2553_ | _2396_;
	assign _2555_ = (_2398_ ? _2552_ : _2554_);
	assign _2556_ = (_2400_ ? _2555_ : _2553_);
	assign _2557_ = (_2406_ ? _2551_ : _2556_);
	assign _2558_ = (_2415_ ? _2546_ : _2557_);
	assign _2559_ = _2394_ | _1617_;
	assign _2560_ = (_2398_ ? _2407_ : _2559_);
	assign _2561_ = (_2400_ ? _2407_ : _2560_);
	assign _2562_ = _2553_ | ~_2396_;
	assign _2563_ = (_2398_ ? _2553_ : _2562_);
	assign _2564_ = _2512_ | _2398_;
	assign _2565_ = (_2400_ ? _2563_ : _2564_);
	assign _2566_ = (_2406_ ? _2561_ : _2565_);
	assign _2567_ = _2394_ | _1626_;
	assign _2568_ = (_2396_ ? _2512_ : _2567_);
	assign _2569_ = (_2396_ ? _2567_ : _2407_);
	assign _2570_ = (_2398_ ? _2568_ : _2569_);
	assign _2571_ = _2394_ | _1631_;
	assign _2572_ = _2394_ | _1632_;
	assign _2573_ = (_2398_ ? _2571_ : _2572_);
	assign _2574_ = (_2400_ ? _2570_ : _2573_);
	assign _2575_ = (_2396_ ? _2532_ : _2567_);
	assign _2576_ = (_2398_ ? _2532_ : _2575_);
	assign _2577_ = (_2398_ ? _2567_ : _2512_);
	assign _2578_ = (_2400_ ? _2576_ : _2577_);
	assign _2579_ = (_2406_ ? _2574_ : _2578_);
	assign _2580_ = (_2415_ ? _2566_ : _2579_);
	assign _2581_ = (_2434_ ? _2558_ : _2580_);
	assign _2582_ = (_2470_ ? _2531_ : _2581_);
	assign _2583_ = (_2474_ ? _2471_ : _2582_);
	assign _2584_ = _2583_ | _2388_;
	assign _2585_ = _2306_ & ~_2584_;
	assign _2586_ = (_2286_ ? _2272_ : _2585_);
	assign _2587_ = (_1978_ ? _1960_ : _2586_);
	assign _0093_ = (_1663_ ? _1646_ : _2587_);
	assign _2588_ = ~\mchip.game2.jumping_inst.frame [3];
	assign _2589_ = \mchip.game2.jumping_inst.frame [2] & ~\mchip.game2.jumping_inst.frame [0];
	assign _2590_ = ~_0957_;
	assign _2591_ = (\mchip.game2.jumping_inst.frame [2] ? \mchip.game2.jumping_inst.frame [0] : _2590_);
	assign _2592_ = (\mchip.game2.jumping_inst.frame [3] ? _2591_ : _2589_);
	assign _2593_ = ~_2589_;
	assign _2594_ = (\mchip.game2.jumping_inst.frame [2] ? \mchip.game2.jumping_inst.frame [0] : _0990_);
	assign _2595_ = (\mchip.game2.jumping_inst.frame [3] ? _2594_ : _2593_);
	assign _2596_ = (\mchip.game2.jumping_inst.frame [4] ? _2595_ : _2592_);
	assign _2597_ = \mchip.game2.jumping_inst.frame [2] & ~_0989_;
	assign _2598_ = ~(\mchip.game2.jumping_inst.frame [1] | \mchip.game2.jumping_inst.frame [0]);
	assign _2599_ = ~(_2598_ | _0973_);
	assign _2600_ = (\mchip.game2.jumping_inst.frame [2] ? _2599_ : _0957_);
	assign _2601_ = (\mchip.game2.jumping_inst.frame [3] ? _2600_ : _2597_);
	assign _2602_ = _0962_ & ~_2601_;
	assign _0000_[0] = (\mchip.game2.jumping_inst.frame [5] ? _2602_ : _2596_);
	assign _2603_ = _2598_ | _0957_;
	assign _2604_ = (\mchip.game2.jumping_inst.frame [2] ? _2603_ : \mchip.game2.jumping_inst.frame [0]);
	assign _2605_ = _2603_ | _0976_;
	assign _2606_ = (\mchip.game2.jumping_inst.frame [3] ? _2605_ : _2604_);
	assign _2607_ = (\mchip.game2.jumping_inst.frame [2] ? \mchip.game2.jumping_inst.frame [1] : \mchip.game2.jumping_inst.frame [0]);
	assign _2608_ = (\mchip.game2.jumping_inst.frame [2] ? _2603_ : _0990_);
	assign _2609_ = (\mchip.game2.jumping_inst.frame [3] ? _2608_ : _2607_);
	assign _2610_ = (\mchip.game2.jumping_inst.frame [4] ? _2609_ : _2606_);
	assign _2611_ = \mchip.game2.jumping_inst.frame [2] & ~\mchip.game2.jumping_inst.frame [1];
	assign _2612_ = ~_2611_;
	assign _2613_ = (\mchip.game2.jumping_inst.frame [3] ? _2612_ : _2607_);
	assign _2614_ = (\mchip.game2.jumping_inst.frame [4] ? _0989_ : _2613_);
	assign _0000_[1] = (\mchip.game2.jumping_inst.frame [5] ? _2614_ : _2610_);
	assign _2615_ = (\mchip.game2.jumping_inst.frame [2] ? _0974_ : _0995_);
	assign _2616_ = (\mchip.game2.jumping_inst.frame [2] ? _0989_ : \mchip.game2.jumping_inst.frame [0]);
	assign _2617_ = (\mchip.game2.jumping_inst.frame [3] ? _2616_ : _2615_);
	assign _2618_ = \mchip.game2.jumping_inst.frame [2] | ~\mchip.game2.jumping_inst.frame [1];
	assign _2619_ = (\mchip.game2.jumping_inst.frame [2] ? _2590_ : _0990_);
	assign _2620_ = (\mchip.game2.jumping_inst.frame [3] ? _2619_ : _2618_);
	assign _2621_ = (\mchip.game2.jumping_inst.frame [4] ? _2620_ : _2617_);
	assign _2622_ = ~\mchip.game2.jumping_inst.frame [1];
	assign _2623_ = (\mchip.game2.jumping_inst.frame [2] ? \mchip.game2.jumping_inst.frame [0] : _0995_);
	assign _2624_ = (\mchip.game2.jumping_inst.frame [2] ? _0995_ : \mchip.game2.jumping_inst.frame [0]);
	assign _2625_ = (\mchip.game2.jumping_inst.frame [3] ? _2624_ : _2623_);
	assign _2626_ = (\mchip.game2.jumping_inst.frame [4] ? _2622_ : _2625_);
	assign _0000_[2] = (\mchip.game2.jumping_inst.frame [5] ? _2626_ : _2621_);
	assign _2627_ = (\mchip.game2.jumping_inst.frame [2] ? _0989_ : _0973_);
	assign _2628_ = ~(\mchip.game2.jumping_inst.frame [2] | \mchip.game2.jumping_inst.frame [1]);
	assign _2629_ = _2628_ | _2611_;
	assign _2630_ = (\mchip.game2.jumping_inst.frame [3] ? _2629_ : _2627_);
	assign _2631_ = (\mchip.game2.jumping_inst.frame [3] ? _0989_ : _2622_);
	assign _2632_ = ~(_2631_ & _0976_);
	assign _2633_ = (\mchip.game2.jumping_inst.frame [4] ? _2632_ : _2630_);
	assign _2634_ = (\mchip.game2.jumping_inst.frame [2] ? _0995_ : _2598_);
	assign _2635_ = (\mchip.game2.jumping_inst.frame [2] ? _0989_ : _0995_);
	assign _2636_ = (\mchip.game2.jumping_inst.frame [3] ? _2635_ : _2634_);
	assign _2637_ = (\mchip.game2.jumping_inst.frame [4] ? _2598_ : _2636_);
	assign _0000_[3] = (\mchip.game2.jumping_inst.frame [5] ? _2637_ : _2633_);
	assign _2638_ = (\mchip.game2.jumping_inst.frame [2] ? _2622_ : _0957_);
	assign _2639_ = _2611_ | ~_2618_;
	assign _2640_ = (\mchip.game2.jumping_inst.frame [3] ? _2639_ : _2638_);
	assign _2641_ = ~(_0989_ & _0976_);
	assign _2642_ = \mchip.game2.jumping_inst.frame [3] & ~_2641_;
	assign _2643_ = (\mchip.game2.jumping_inst.frame [4] ? _2642_ : _2640_);
	assign _2644_ = \mchip.game2.jumping_inst.frame [2] & ~_2598_;
	assign _2645_ = ~_2644_;
	assign _2646_ = _2598_ ^ _0976_;
	assign _2647_ = (\mchip.game2.jumping_inst.frame [3] ? _2646_ : _2645_);
	assign _2648_ = _0962_ & ~_2647_;
	assign _0000_[4] = (\mchip.game2.jumping_inst.frame [5] ? _2648_ : _2643_);
	assign _2649_ = \mchip.game2.jumping_inst.frame [2] & \mchip.game2.jumping_inst.frame [1];
	assign _2650_ = _2649_ ^ _2588_;
	assign _2651_ = _2644_ ^ _2588_;
	assign _2652_ = (\mchip.game2.jumping_inst.frame [5] ? _2651_ : _2650_);
	assign _0000_[5] = _0962_ & ~_2652_;
	assign _2653_ = _2649_ & ~_2588_;
	assign _2654_ = _2653_ | \mchip.game2.jumping_inst.frame [4];
	assign _2655_ = _2644_ | \mchip.game2.jumping_inst.frame [3];
	assign _2656_ = _0962_ & ~_2655_;
	assign _0000_[6] = (\mchip.game2.jumping_inst.frame [5] ? _2656_ : _2654_);
	assign _3621_[0] = ~\mchip.game2.no_jump_ctr [0];
	assign _3622_[0] = ~\mchip.game2.start_ctr [0];
	assign _0027_ = ~_0372_;
	assign _2657_ = ~(_3219_ & _3206_);
	assign _2658_ = _2657_ | _3217_;
	assign _2659_ = _3213_ & ~_2658_;
	assign _2660_ = _3206_ & ~_3219_;
	assign _2661_ = ~(_2660_ | _3217_);
	assign _2662_ = _3215_ & ~_2661_;
	assign _2663_ = _3213_ & ~_2662_;
	assign _2664_ = ~(_2663_ | _3188_);
	assign _2665_ = _2664_ | _2659_;
	assign _2666_ = _3217_ | _3191_;
	assign _2667_ = _2666_ | ~_3213_;
	assign _2668_ = ~(_3217_ | _3200_);
	assign _2669_ = _3215_ & ~_2668_;
	assign _2670_ = _3213_ & ~_2669_;
	assign _2671_ = _3197_ & ~_2670_;
	assign _2672_ = _2667_ & ~_2671_;
	assign _0151_ = _2672_ | _2665_;
	assign _2673_ = _2273_ & _1731_;
	assign _2674_ = _2673_ | _3181_;
	assign _2675_ = _3179_ | ~_2273_;
	assign _2676_ = \mchip.game2.vga_inst.haddr [6] | ~\mchip.game2.vga_inst.haddr [7];
	assign _2677_ = _2676_ | _0254_;
	assign _2678_ = _2677_ | _2675_;
	assign _2679_ = _2678_ | _3186_;
	assign _2680_ = _2676_ | _0239_;
	assign _2681_ = _2680_ & ~_1270_;
	assign _2682_ = _2273_ & ~_2681_;
	assign _2683_ = _2682_ | _3181_;
	assign _2684_ = _2679_ & ~_2683_;
	assign _0150_ = _2684_ | _2674_;
	assign _2685_ = _0253_ & ~_1199_;
	assign _3625_[5] = _2685_ ^ \mchip.game2.vga_inst.haddr [5];
	assign _2686_ = _0253_ & ~_1717_;
	assign _3625_[6] = _2686_ ^ \mchip.game2.vga_inst.haddr [6];
	assign _2687_ = _2686_ & ~_1256_;
	assign _3625_[7] = _2687_ ^ \mchip.game2.vga_inst.haddr [7];
	assign _2688_ = _1731_ & _0253_;
	assign _3625_[8] = _2688_ ^ \mchip.game2.vga_inst.haddr [8];
	assign _2689_ = _2688_ & ~_1269_;
	assign _3625_[9] = _2689_ ^ \mchip.game2.vga_inst.haddr [9];
	assign _3624_[1] = \mchip.game2.start_ctr [0] ^ \mchip.game2.start_ctr [1];
	assign _2690_ = \mchip.game2.start_ctr [0] & \mchip.game2.start_ctr [1];
	assign _3624_[2] = _2690_ ^ \mchip.game2.start_ctr [2];
	assign _2691_ = _2690_ & \mchip.game2.start_ctr [2];
	assign _3624_[3] = _2691_ ^ \mchip.game2.start_ctr [3];
	assign _2692_ = ~(\mchip.game2.start_ctr [2] & \mchip.game2.start_ctr [3]);
	assign _2693_ = _2690_ & ~_2692_;
	assign _3624_[4] = _2693_ ^ \mchip.game2.start_ctr [4];
	assign _2694_ = _2693_ & \mchip.game2.start_ctr [4];
	assign _3624_[5] = _2694_ ^ \mchip.game2.start_ctr [5];
	assign _2695_ = ~(\mchip.game2.start_ctr [5] & \mchip.game2.start_ctr [4]);
	assign _2696_ = _2693_ & ~_2695_;
	assign _3624_[6] = _2696_ ^ \mchip.game2.start_ctr [6];
	assign _2697_ = _2696_ & \mchip.game2.start_ctr [6];
	assign _3624_[7] = _2697_ ^ \mchip.game2.start_ctr [7];
	assign _2698_ = ~(\mchip.game2.start_ctr [6] & \mchip.game2.start_ctr [7]);
	assign _2699_ = ~(_2698_ | _2695_);
	assign _2700_ = ~(_2699_ & _2693_);
	assign _3624_[8] = ~(_2700_ ^ \mchip.game2.start_ctr [8]);
	assign _2701_ = \mchip.game2.start_ctr [8] & ~_2700_;
	assign _3624_[9] = _2701_ ^ \mchip.game2.start_ctr [9];
	assign _2702_ = _3258_ & ~_2700_;
	assign _3624_[10] = _2702_ ^ \mchip.game2.start_ctr [10];
	assign _2703_ = _2702_ & \mchip.game2.start_ctr [10];
	assign _3624_[11] = _2703_ ^ \mchip.game2.start_ctr [11];
	assign _2704_ = \mchip.game2.start_ctr [10] & \mchip.game2.start_ctr [11];
	assign _2705_ = ~(_2704_ & _3258_);
	assign _2706_ = ~(_2705_ | _2700_);
	assign _3624_[12] = _2706_ ^ \mchip.game2.start_ctr [12];
	assign _2707_ = _2706_ & \mchip.game2.start_ctr [12];
	assign _3624_[13] = _2707_ ^ \mchip.game2.start_ctr [13];
	assign _2708_ = ~(\mchip.game2.start_ctr [12] & \mchip.game2.start_ctr [13]);
	assign _2709_ = _2706_ & ~_2708_;
	assign _3624_[14] = _2709_ ^ \mchip.game2.start_ctr [14];
	assign _2710_ = _2709_ & \mchip.game2.start_ctr [14];
	assign _3624_[15] = _2710_ ^ \mchip.game2.start_ctr [15];
	assign _2711_ = _2708_ | _3255_;
	assign _2712_ = _2711_ | _2705_;
	assign _2713_ = ~(_2712_ | _2700_);
	assign _3624_[16] = _2713_ ^ \mchip.game2.start_ctr [16];
	assign _2714_ = _2713_ & \mchip.game2.start_ctr [16];
	assign _3624_[17] = _2714_ ^ \mchip.game2.start_ctr [17];
	assign _2715_ = ~(\mchip.game2.start_ctr [17] & \mchip.game2.start_ctr [16]);
	assign _2716_ = _2713_ & ~_2715_;
	assign _3624_[18] = _2716_ ^ \mchip.game2.start_ctr [18];
	assign _2717_ = _2716_ & \mchip.game2.start_ctr [18];
	assign _3624_[19] = _2717_ ^ \mchip.game2.start_ctr [19];
	assign _2718_ = ~(\mchip.game2.start_ctr [18] & \mchip.game2.start_ctr [19]);
	assign _2719_ = _2718_ | _2715_;
	assign _2720_ = _2713_ & ~_2719_;
	assign _3624_[20] = _2720_ ^ \mchip.game2.start_ctr [20];
	assign _2721_ = _2720_ & \mchip.game2.start_ctr [20];
	assign _3624_[21] = _2721_ ^ \mchip.game2.start_ctr [21];
	assign _2722_ = ~(\mchip.game2.start_ctr [20] & \mchip.game2.start_ctr [21]);
	assign _2723_ = _2720_ & ~_2722_;
	assign _3624_[22] = _2723_ ^ \mchip.game2.start_ctr [22];
	assign _2724_ = _2723_ & \mchip.game2.start_ctr [22];
	assign _3624_[23] = _2724_ ^ \mchip.game2.start_ctr [23];
	assign _2725_ = _2722_ | ~_3244_;
	assign _2726_ = _2725_ | _2719_;
	assign _2727_ = _2713_ & ~_2726_;
	assign _3624_[24] = _2727_ ^ \mchip.game2.start_ctr [24];
	assign _2728_ = _2727_ & \mchip.game2.start_ctr [24];
	assign _3624_[25] = _2728_ ^ \mchip.game2.start_ctr [25];
	assign _2729_ = ~(\mchip.game2.start_ctr [24] & \mchip.game2.start_ctr [25]);
	assign _2730_ = _2727_ & ~_2729_;
	assign _3624_[26] = _2730_ ^ \mchip.game2.start_ctr [26];
	assign _2731_ = _2730_ & \mchip.game2.start_ctr [26];
	assign _3624_[27] = _2731_ ^ \mchip.game2.start_ctr [27];
	assign _2732_ = ~(\mchip.game2.start_ctr [26] & \mchip.game2.start_ctr [27]);
	assign _2733_ = _2732_ | _2729_;
	assign _2734_ = _2727_ & ~_2733_;
	assign _3624_[28] = _2734_ ^ \mchip.game2.start_ctr [28];
	assign _2735_ = _2734_ & \mchip.game2.start_ctr [28];
	assign _3624_[29] = _2735_ ^ \mchip.game2.start_ctr [29];
	assign _2736_ = ~(\mchip.game2.start_ctr [29] & \mchip.game2.start_ctr [28]);
	assign _2737_ = _2734_ & ~_2736_;
	assign _3624_[30] = _2737_ ^ \mchip.game2.start_ctr [30];
	assign _2738_ = _2737_ & \mchip.game2.start_ctr [30];
	assign _3624_[31] = _2738_ ^ \mchip.game2.start_ctr [31];
	assign _3623_[1] = \mchip.game2.no_jump_ctr [0] ^ \mchip.game2.no_jump_ctr [1];
	assign _2739_ = \mchip.game2.no_jump_ctr [0] & \mchip.game2.no_jump_ctr [1];
	assign _3623_[2] = _2739_ ^ \mchip.game2.no_jump_ctr [2];
	assign _2740_ = _2739_ & \mchip.game2.no_jump_ctr [2];
	assign _3623_[3] = _2740_ ^ \mchip.game2.no_jump_ctr [3];
	assign _2741_ = ~(\mchip.game2.no_jump_ctr [2] & \mchip.game2.no_jump_ctr [3]);
	assign _2742_ = _2739_ & ~_2741_;
	assign _3623_[4] = _2742_ ^ \mchip.game2.no_jump_ctr [4];
	assign _2743_ = _2742_ & \mchip.game2.no_jump_ctr [4];
	assign _3623_[5] = _2743_ ^ \mchip.game2.no_jump_ctr [5];
	assign _2744_ = ~(\mchip.game2.no_jump_ctr [4] & \mchip.game2.no_jump_ctr [5]);
	assign _2745_ = _2742_ & ~_2744_;
	assign _3623_[6] = _2745_ ^ \mchip.game2.no_jump_ctr [6];
	assign _2746_ = _2745_ & \mchip.game2.no_jump_ctr [6];
	assign _3623_[7] = _2746_ ^ \mchip.game2.no_jump_ctr [7];
	assign _2747_ = ~(\mchip.game2.no_jump_ctr [6] & \mchip.game2.no_jump_ctr [7]);
	assign _2748_ = _2747_ | _2744_;
	assign _2749_ = _2742_ & ~_2748_;
	assign _3623_[8] = _2749_ ^ \mchip.game2.no_jump_ctr [8];
	assign _2750_ = _2749_ & \mchip.game2.no_jump_ctr [8];
	assign _3623_[9] = _2750_ ^ \mchip.game2.no_jump_ctr [9];
	assign _2751_ = ~(\mchip.game2.no_jump_ctr [8] & \mchip.game2.no_jump_ctr [9]);
	assign _2752_ = _2749_ & ~_2751_;
	assign _3623_[10] = _2752_ ^ \mchip.game2.no_jump_ctr [10];
	assign _2753_ = _2752_ & \mchip.game2.no_jump_ctr [10];
	assign _3623_[11] = _2753_ ^ \mchip.game2.no_jump_ctr [11];
	assign _2754_ = ~(\mchip.game2.no_jump_ctr [10] & \mchip.game2.no_jump_ctr [11]);
	assign _2755_ = _2754_ | _2751_;
	assign _2756_ = _2749_ & ~_2755_;
	assign _3623_[12] = _2756_ ^ \mchip.game2.no_jump_ctr [12];
	assign _2757_ = _2756_ & \mchip.game2.no_jump_ctr [12];
	assign _3623_[13] = _2757_ ^ \mchip.game2.no_jump_ctr [13];
	assign _2758_ = ~(\mchip.game2.no_jump_ctr [12] & \mchip.game2.no_jump_ctr [13]);
	assign _2759_ = _2756_ & ~_2758_;
	assign _3623_[14] = _2759_ ^ \mchip.game2.no_jump_ctr [14];
	assign _2760_ = _2759_ & \mchip.game2.no_jump_ctr [14];
	assign _3623_[15] = _2760_ ^ \mchip.game2.no_jump_ctr [15];
	assign _2761_ = ~(\mchip.game2.no_jump_ctr [14] & \mchip.game2.no_jump_ctr [15]);
	assign _2762_ = _2761_ | _2758_;
	assign _2763_ = _2762_ | _2755_;
	assign _2764_ = _2749_ & ~_2763_;
	assign _3623_[16] = _2764_ ^ \mchip.game2.no_jump_ctr [16];
	assign _2765_ = _2764_ & \mchip.game2.no_jump_ctr [16];
	assign _3623_[17] = _2765_ ^ \mchip.game2.no_jump_ctr [17];
	assign _2766_ = ~(\mchip.game2.no_jump_ctr [16] & \mchip.game2.no_jump_ctr [17]);
	assign _2767_ = _2764_ & ~_2766_;
	assign _3623_[18] = _2767_ ^ \mchip.game2.no_jump_ctr [18];
	assign _2768_ = _2767_ & \mchip.game2.no_jump_ctr [18];
	assign _3623_[19] = _2768_ ^ \mchip.game2.no_jump_ctr [19];
	assign _0091_ = \mchip.game2.rng_inst.out [1] ^ \mchip.game2.rng_inst.out [4];
	assign _2769_ = ~_3450_;
	assign _2770_ = _2769_ & ~_3454_;
	assign _2771_ = _3447_ | _3442_;
	assign _2772_ = _2770_ & ~_2771_;
	assign _2773_ = _3470_ | _3436_;
	assign _2774_ = _3441_ | _3435_;
	assign _2775_ = _2774_ | _2773_;
	assign _2776_ = _2772_ & ~_2775_;
	assign _2777_ = _2776_ | _3454_;
	assign _2778_ = ~(_3484_ & _3426_);
	assign _2779_ = _2778_ | _3432_;
	assign _2780_ = _2777_ & ~_2779_;
	assign _2781_ = _3433_ & ~_2780_;
	assign _2782_ = _3450_ | _3447_;
	assign _2783_ = _2782_ | _3455_;
	assign _2784_ = _3437_ | _3435_;
	assign _2785_ = _2784_ | _3443_;
	assign _2786_ = _2785_ | _2783_;
	assign _2787_ = _3432_ | ~_3426_;
	assign _2788_ = _2787_ | _2786_;
	assign _2789_ = _3470_ & ~_2788_;
	assign _2790_ = _3454_ & ~_2778_;
	assign _2791_ = _3426_ & ~_2790_;
	assign _2792_ = _2770_ & ~_2778_;
	assign _2793_ = _3442_ & ~_3447_;
	assign _2794_ = _3441_ & _3435_;
	assign _2795_ = _2793_ & ~_2794_;
	assign _2796_ = _2771_ & ~_2795_;
	assign _2797_ = _2792_ & ~_2796_;
	assign _2798_ = _2791_ & ~_2797_;
	assign _2799_ = _2798_ | _3432_;
	assign _2800_ = _2799_ | _2789_;
	assign _2801_ = _2781_ & ~_2800_;
	assign _2802_ = ~\mchip.game2.cactus_type [0];
	assign _2803_ = _0536_ & _0521_;
	assign _2804_ = _2803_ | ~_0525_;
	assign _2805_ = _2804_ | _0528_;
	assign _2806_ = _2805_ | _2802_;
	assign _2807_ = _2806_ | _3450_;
	assign _2808_ = _2807_ | _3470_;
	assign _2809_ = _2808_ | _3436_;
	assign _2810_ = _2809_ | _3435_;
	assign _2811_ = ~(_0577_ & _0525_);
	assign _2812_ = (_0528_ ? _0562_ : _2811_);
	assign _2813_ = _2812_ | _2802_;
	assign _2814_ = _2813_ | _3450_;
	assign _2815_ = _2814_ | _3470_;
	assign _2816_ = _3470_ & ~_2814_;
	assign _2817_ = _2815_ & ~_2816_;
	assign _2818_ = _0521_ | ~_0555_;
	assign _2819_ = ~(_2818_ | _0525_);
	assign _2820_ = _2819_ & ~_0528_;
	assign _2821_ = (_3470_ ? _0551_ : _2820_);
	assign _2822_ = _2821_ | _2802_;
	assign _2823_ = _2822_ | _3450_;
	assign _2824_ = (_3436_ ? _2817_ : _2823_);
	assign _2825_ = _3198_ | _0516_;
	assign _2826_ = ~(_2825_ | _0521_);
	assign _2827_ = ~(_2826_ & _0525_);
	assign _2828_ = _2827_ | _0528_;
	assign _2829_ = _2828_ | _2802_;
	assign _2830_ = _2829_ | _3450_;
	assign _2831_ = _2830_ | _3470_;
	assign _2832_ = _3470_ & ~_2830_;
	assign _2833_ = _2831_ & ~_2832_;
	assign _2834_ = (_0521_ ? _0541_ : _0518_);
	assign _2835_ = (_0525_ ? _2834_ : _0554_);
	assign _2836_ = (_0528_ ? _2818_ : _2835_);
	assign _2837_ = ~(_0522_ & _0518_);
	assign _2838_ = _0554_ & ~_2837_;
	assign _2839_ = ~(_2838_ & _0528_);
	assign _2840_ = (_3470_ ? _2836_ : _2839_);
	assign _2841_ = _2840_ | _2802_;
	assign _2842_ = _2841_ | _3450_;
	assign _2843_ = (_3436_ ? _2833_ : _2842_);
	assign _2844_ = (_3435_ ? _2824_ : _2843_);
	assign _2845_ = (_3441_ ? _2810_ : _2844_);
	assign _2846_ = _0571_ & ~_0521_;
	assign _2847_ = _2846_ | ~_0525_;
	assign _2848_ = _2847_ & ~_0528_;
	assign _2849_ = _2848_ | _2802_;
	assign _2850_ = _2849_ | _3450_;
	assign _2851_ = _0517_ | _0515_;
	assign _2852_ = ~(_2851_ | _0521_);
	assign _2853_ = ~(_2852_ & _0528_);
	assign _2854_ = _2853_ | _2802_;
	assign _2855_ = _2854_ | _3450_;
	assign _2856_ = (_3470_ ? _2850_ : _2855_);
	assign _2857_ = ~(_0542_ & _0525_);
	assign _2858_ = (_0528_ ? _0549_ : _2857_);
	assign _2859_ = _2858_ | _2802_;
	assign _2860_ = _2859_ | _3450_;
	assign _2861_ = (_3470_ ? _2855_ : _2860_);
	assign _2862_ = (_3436_ ? _2856_ : _2861_);
	assign _2863_ = _0540_ | _2802_;
	assign _2864_ = _2802_ & ~_0540_;
	assign _2865_ = _2863_ & ~_2864_;
	assign _2866_ = _0544_ | _2802_;
	assign _2867_ = _2802_ & ~_0544_;
	assign _2868_ = _2866_ & ~_2867_;
	assign _2869_ = (_3470_ ? _2865_ : _2868_);
	assign _2870_ = _2869_ | _3450_;
	assign _2871_ = (_0521_ ? _0541_ : _0517_);
	assign _2872_ = ~(_2871_ & _0525_);
	assign _2873_ = _2872_ | _0528_;
	assign _2874_ = (\mchip.game2.cactus_type [0] ? _2873_ : _0529_);
	assign _2875_ = (_0528_ ? _0532_ : _2872_);
	assign _2876_ = (\mchip.game2.cactus_type [0] ? _2875_ : _0533_);
	assign _2877_ = (_3470_ ? _2874_ : _2876_);
	assign _2878_ = _2877_ | _3450_;
	assign _2879_ = (_3436_ ? _2870_ : _2878_);
	assign _2880_ = (_3435_ ? _2862_ : _2879_);
	assign _2881_ = (_3470_ ? _0551_ : _0564_);
	assign _2882_ = _2881_ & ~\mchip.game2.cactus_type [0];
	assign _2883_ = _2882_ | _3450_;
	assign _2884_ = (\mchip.game2.cactus_type [0] ? _0564_ : _0551_);
	assign _2885_ = _2884_ | _3450_;
	assign _2886_ = (_0517_ ? _0515_ : _3189_);
	assign _2887_ = _2886_ & _0521_;
	assign _2888_ = ~(_2887_ & _0525_);
	assign _2889_ = _2888_ | _0528_;
	assign _2890_ = (\mchip.game2.cactus_type [0] ? _2889_ : _0559_);
	assign _2891_ = _2890_ | _3450_;
	assign _2892_ = (_3470_ ? _2885_ : _2891_);
	assign _2893_ = (_3436_ ? _2883_ : _2892_);
	assign _2894_ = (_0525_ ? _0572_ : _0570_);
	assign _2895_ = _2894_ | _0528_;
	assign _2896_ = (\mchip.game2.cactus_type [0] ? _2895_ : _0579_);
	assign _2897_ = _2896_ | _3450_;
	assign _2898_ = (_3470_ ? _2891_ : _2897_);
	assign _2899_ = ~(_0521_ & _0518_);
	assign _2900_ = (_0525_ ? _2899_ : _0572_);
	assign _2901_ = _0528_ | ~_2900_;
	assign _2902_ = (\mchip.game2.cactus_type [0] ? _2901_ : _0574_);
	assign _2903_ = _2902_ | _3450_;
	assign _2904_ = _2903_ | _3471_;
	assign _2905_ = (_3436_ ? _2898_ : _2904_);
	assign _2906_ = (_3435_ ? _2893_ : _2905_);
	assign _2907_ = (_3441_ ? _2880_ : _2906_);
	assign _2908_ = (_3442_ ? _2845_ : _2907_);
	assign _2909_ = _2908_ | _3447_;
	assign _0022_ = _2801_ & ~_2909_;
	assign _2910_ = _3432_ ^ \mchip.game2.scroll_inst.pos [10];
	assign _2911_ = ~(_2910_ | _3426_);
	assign _2912_ = _3432_ & ~_0301_;
	assign _2913_ = _2911_ & ~_2912_;
	assign _2914_ = _3434_ & ~_3454_;
	assign _2915_ = _2914_ & ~_3451_;
	assign _2916_ = _3450_ & ~_3447_;
	assign _2917_ = _2916_ & _2914_;
	assign _2918_ = _3442_ | _3441_;
	assign _2919_ = _3438_ & ~_2918_;
	assign _2920_ = _2917_ & ~_2919_;
	assign _2921_ = _2920_ | _2915_;
	assign _2922_ = _2913_ & ~_2921_;
	assign _2923_ = _2921_ ^ _3479_;
	assign _2924_ = _3479_ & ~_2921_;
	assign _2925_ = _2924_ ^ _2910_;
	assign _2926_ = _2911_ & ~_2921_;
	assign _2927_ = _2926_ ^ _2912_;
	assign _2928_ = _2927_ | _2925_;
	assign _2929_ = _2928_ | _2923_;
	assign _2930_ = _2926_ & ~_2912_;
	assign _2931_ = _2930_ | _2922_;
	assign _2932_ = _2931_ | _2929_;
	assign _2933_ = ~_3454_;
	assign _2934_ = _2916_ & ~_2919_;
	assign _2935_ = _3451_ & ~_2934_;
	assign _2936_ = _2933_ & ~_2935_;
	assign _2937_ = _2936_ ^ _3434_;
	assign _2938_ = _2923_ & ~_2937_;
	assign _2939_ = _2928_ | ~_2938_;
	assign _2940_ = ~(_2939_ | _2931_);
	assign _2941_ = _2935_ ^ _2933_;
	assign _2942_ = ~_2941_;
	assign _2943_ = ~(_2919_ ^ _3447_);
	assign _2944_ = _3474_ ^ _3442_;
	assign _2945_ = _2943_ & ~_2944_;
	assign _2946_ = _2919_ & ~_3447_;
	assign _2947_ = _2946_ ^ _2769_;
	assign _2948_ = _2947_ | _2941_;
	assign _2949_ = _2945_ & ~_2948_;
	assign _2950_ = _3441_ ^ _3438_;
	assign _2951_ = _2950_ | _3473_;
	assign _2952_ = _2951_ | _3508_;
	assign _2953_ = _2949_ & ~_2952_;
	assign _2954_ = _2942_ & ~_2953_;
	assign _2955_ = _2940_ & ~_2954_;
	assign _2956_ = _2932_ & ~_2955_;
	assign _2957_ = _2956_ | _2922_;
	assign _2958_ = _2944_ & _2943_;
	assign _2959_ = _2948_ | ~_2958_;
	assign _2960_ = _3473_ | ~_2950_;
	assign _2961_ = _2960_ | _3472_;
	assign _2962_ = ~(_2961_ | _2959_);
	assign _2963_ = ~(_2962_ & _2940_);
	assign _2964_ = ~(_2963_ | _2922_);
	assign _2965_ = _2938_ & ~_2942_;
	assign _2966_ = _2923_ & ~_2965_;
	assign _2967_ = _2938_ & ~_2948_;
	assign _2968_ = _2950_ & _3473_;
	assign _2969_ = _2968_ | ~_2958_;
	assign _2970_ = _2969_ & ~_2945_;
	assign _2971_ = _2967_ & ~_2970_;
	assign _2972_ = _2966_ & ~_2971_;
	assign _2973_ = _2931_ | _2928_;
	assign _2974_ = _2973_ | _2922_;
	assign _2975_ = _2974_ | _2972_;
	assign _2976_ = _2975_ | _2922_;
	assign _2977_ = _2976_ | _2964_;
	assign _2978_ = _2957_ & ~_2977_;
	assign _2979_ = ~(\mchip.game2.scroll_inst.pos [4] ^ \mchip.game2.vga_inst.haddr [4]);
	assign _2980_ = _2979_ & ~_3400_;
	assign _2981_ = _2979_ ^ _3400_;
	assign _2982_ = ~(\mchip.game2.scroll_inst.pos [3] ^ \mchip.game2.vga_inst.haddr [3]);
	assign _2983_ = _3410_ | ~_2982_;
	assign _2984_ = _2982_ ^ _3410_;
	assign _2985_ = ~(\mchip.game2.scroll_inst.pos [2] ^ \mchip.game2.vga_inst.haddr [2]);
	assign _2986_ = _3406_ | ~_2985_;
	assign _2987_ = ~(_2986_ | _2984_);
	assign _2988_ = _2983_ & ~_2987_;
	assign _2989_ = ~(\mchip.game2.scroll_inst.pos [1] ^ \mchip.game2.vga_inst.haddr [1]);
	assign _2990_ = _2989_ & _3405_;
	assign _2991_ = ~(_2985_ ^ _3406_);
	assign _2992_ = _2984_ | ~_2991_;
	assign _2993_ = _2990_ & ~_2992_;
	assign _2994_ = _2988_ & ~_2993_;
	assign _2995_ = ~(_2994_ | _2981_);
	assign _2996_ = _2995_ | _2980_;
	assign _2997_ = ~(\mchip.game2.scroll_inst.pos [5] ^ \mchip.game2.vga_inst.haddr [5]);
	assign _2998_ = ~(_2997_ ^ _3415_);
	assign _2999_ = _2998_ ^ _2996_;
	assign _3000_ = _2989_ ^ _3405_;
	assign _3001_ = ~\mchip.game2.cactus_type [2];
	assign _3002_ = _2805_ | _3001_;
	assign _3003_ = _2997_ & ~_3415_;
	assign _3004_ = _2998_ & _2980_;
	assign _3005_ = _3004_ | _3003_;
	assign _3006_ = _2981_ | ~_2998_;
	assign _3007_ = ~(_3006_ | _2994_);
	assign _3008_ = _3007_ | _3005_;
	assign _3009_ = _3393_ ^ _3389_;
	assign _3010_ = _3009_ ^ _3008_;
	assign _3011_ = _3010_ | _3002_;
	assign _3012_ = _3011_ | _3470_;
	assign _3013_ = _3012_ | _3000_;
	assign _3014_ = _2991_ ^ _2990_;
	assign _3015_ = _3014_ | _3013_;
	assign _3016_ = _2991_ & _2990_;
	assign _3017_ = _2986_ & ~_3016_;
	assign _3018_ = _3017_ ^ _2984_;
	assign _3019_ = _2812_ | _3001_;
	assign _3020_ = _3019_ | _3010_;
	assign _3021_ = _3020_ | _3470_;
	assign _3022_ = _3470_ & ~_3020_;
	assign _3023_ = _3021_ & ~_3022_;
	assign _3024_ = _2821_ | _3001_;
	assign _3025_ = _3024_ | _3010_;
	assign _3026_ = (_3000_ ? _3023_ : _3025_);
	assign _3027_ = _2828_ | _3001_;
	assign _3028_ = _3027_ | _3010_;
	assign _3029_ = _3028_ | _3470_;
	assign _3030_ = _3470_ & ~_3028_;
	assign _3031_ = _3029_ & ~_3030_;
	assign _3032_ = _2840_ | _3001_;
	assign _3033_ = _3032_ | _3010_;
	assign _3034_ = (_3000_ ? _3031_ : _3033_);
	assign _3035_ = (_3014_ ? _3026_ : _3034_);
	assign _3036_ = (_3018_ ? _3015_ : _3035_);
	assign _3037_ = _2994_ ^ _2981_;
	assign _3038_ = _2848_ | _3001_;
	assign _3039_ = _3038_ | _3010_;
	assign _3040_ = _2853_ | _3001_;
	assign _3041_ = _3040_ | _3010_;
	assign _3042_ = (_3470_ ? _3039_ : _3041_);
	assign _3043_ = _2858_ | _3001_;
	assign _3044_ = _3043_ | _3010_;
	assign _3045_ = (_3470_ ? _3041_ : _3044_);
	assign _3046_ = (_3000_ ? _3042_ : _3045_);
	assign _3047_ = (_0525_ ? _0532_ : _0577_);
	assign _3048_ = ~(_3047_ & _0568_);
	assign _3049_ = (\mchip.game2.cactus_type [2] ? _0540_ : _3048_);
	assign _3050_ = ~(_0577_ | _0525_);
	assign _3051_ = _3050_ | _0528_;
	assign _3052_ = (\mchip.game2.cactus_type [2] ? _0544_ : _3051_);
	assign _3053_ = (_3470_ ? _3049_ : _3052_);
	assign _3054_ = _3053_ | _3010_;
	assign _3055_ = ~(_0569_ & _0525_);
	assign _3056_ = _3055_ | _0528_;
	assign _3057_ = (\mchip.game2.cactus_type [2] ? _2873_ : _3056_);
	assign _3058_ = _3057_ | _3010_;
	assign _3059_ = _0517_ & _0497_;
	assign _3060_ = ~(_3059_ & _0521_);
	assign _3061_ = _3060_ | _0525_;
	assign _3062_ = (_0528_ ? _3061_ : _3055_);
	assign _3063_ = (\mchip.game2.cactus_type [2] ? _2875_ : _3062_);
	assign _3064_ = _3063_ | _3010_;
	assign _3065_ = (_3470_ ? _3058_ : _3064_);
	assign _3066_ = (_3000_ ? _3054_ : _3065_);
	assign _3067_ = (_3014_ ? _3046_ : _3066_);
	assign _3068_ = ~(_2803_ | _0525_);
	assign _3069_ = (_0528_ ? _3068_ : _0550_);
	assign _3070_ = ~_3068_;
	assign _3071_ = (_0528_ ? _3070_ : _0563_);
	assign _3072_ = ~_3071_;
	assign _3073_ = (_3470_ ? _3069_ : _3072_);
	assign _3074_ = _3001_ & ~_3073_;
	assign _3075_ = (\mchip.game2.cactus_type [2] ? _0564_ : _3071_);
	assign _3076_ = (_0528_ ? _0553_ : _0558_);
	assign _3077_ = (\mchip.game2.cactus_type [2] ? _2889_ : _3076_);
	assign _3078_ = (_3470_ ? _3075_ : _3077_);
	assign _3079_ = (_3000_ ? _3074_ : _3078_);
	assign _3080_ = _3079_ | _3010_;
	assign _3081_ = (\mchip.game2.cactus_type [2] ? _2889_ : _0559_);
	assign _3082_ = (_0525_ ? _0531_ : _0570_);
	assign _3083_ = _3082_ | _0528_;
	assign _3084_ = (\mchip.game2.cactus_type [2] ? _2895_ : _3083_);
	assign _3085_ = (_3470_ ? _3081_ : _3084_);
	assign _3086_ = _3085_ | _3010_;
	assign _3087_ = (\mchip.game2.cactus_type [2] ? _2901_ : _2895_);
	assign _3088_ = _3087_ | _3010_;
	assign _3089_ = _3088_ | ~_3470_;
	assign _3090_ = (_3000_ ? _3086_ : _3089_);
	assign _3091_ = (_3014_ ? _3080_ : _3090_);
	assign _3092_ = (_3018_ ? _3067_ : _3091_);
	assign _3093_ = (_3037_ ? _3036_ : _3092_);
	assign _3094_ = _3093_ | _2999_;
	assign _0021_ = _2978_ & ~_3094_;
	assign _3095_ = \mchip.game2.scroll_inst.tick_time [0] | ~_3171_;
	assign _3096_ = io_in[8] & io_in[11];
	assign _3097_ = ~(_3096_ ^ \mchip.game2.scroll_inst.tick_time [1]);
	assign _3628_[1] = _3097_ ^ _3095_;
	assign _3098_ = \mchip.game2.scroll_inst.tick_time [1] & ~_3096_;
	assign _3099_ = _3097_ & _3095_;
	assign _3100_ = _3099_ | _3098_;
	assign _3101_ = io_in[11] & ~io_in[9];
	assign _3102_ = _3101_ ^ \mchip.game2.scroll_inst.tick_time [2];
	assign _3628_[2] = _3102_ ^ _3100_;
	assign _3103_ = _3101_ & \mchip.game2.scroll_inst.tick_time [2];
	assign _3104_ = _3102_ & _3100_;
	assign _3105_ = _3104_ | _3103_;
	assign _3106_ = io_in[10] & io_in[11];
	assign _3107_ = ~(_3106_ ^ \mchip.game2.scroll_inst.tick_time [3]);
	assign _3628_[3] = _3107_ ^ _3105_;
	assign _3108_ = ~(_3107_ & _3102_);
	assign _3109_ = _3100_ & ~_3108_;
	assign _3110_ = \mchip.game2.scroll_inst.tick_time [3] & ~_3106_;
	assign _3111_ = _3107_ & _3103_;
	assign _3112_ = _3111_ | _3110_;
	assign _3113_ = ~(_3112_ | _3109_);
	assign _3628_[4] = _3113_ ^ \mchip.game2.scroll_inst.tick_time [4];
	assign _3114_ = _3113_ & ~\mchip.game2.scroll_inst.tick_time [4];
	assign _3628_[5] = _3114_ ^ \mchip.game2.scroll_inst.tick_time [5];
	assign _3115_ = \mchip.game2.scroll_inst.tick_time [4] | \mchip.game2.scroll_inst.tick_time [5];
	assign _3116_ = _3113_ & ~_3115_;
	assign _3628_[6] = _3116_ ^ \mchip.game2.scroll_inst.tick_time [6];
	assign _3117_ = _3116_ & ~\mchip.game2.scroll_inst.tick_time [6];
	assign _3628_[7] = _3117_ ^ \mchip.game2.scroll_inst.tick_time [7];
	assign _3118_ = ~\mchip.game2.scroll_inst.tick_time [8];
	assign _3119_ = \mchip.game2.scroll_inst.tick_time [6] | \mchip.game2.scroll_inst.tick_time [7];
	assign _3120_ = ~(_3119_ | _3115_);
	assign _3121_ = _3120_ & ~_3113_;
	assign _3122_ = _3119_ | _3115_;
	assign _3123_ = _3122_ | _3121_;
	assign _3628_[8] = _3123_ ^ _3118_;
	assign _3124_ = _3118_ & ~_3123_;
	assign _3628_[9] = _3124_ ^ \mchip.game2.scroll_inst.tick_time [9];
	assign _3125_ = \mchip.game2.scroll_inst.tick_time [8] | \mchip.game2.scroll_inst.tick_time [9];
	assign _3126_ = ~(_3125_ | _3123_);
	assign _3628_[10] = _3126_ ^ \mchip.game2.scroll_inst.tick_time [10];
	assign _3127_ = _3126_ & ~\mchip.game2.scroll_inst.tick_time [10];
	assign _3628_[11] = _3127_ ^ \mchip.game2.scroll_inst.tick_time [11];
	assign _3128_ = \mchip.game2.scroll_inst.tick_time [10] | \mchip.game2.scroll_inst.tick_time [11];
	assign _3129_ = _3128_ | _3125_;
	assign _3130_ = _3123_ & ~_3129_;
	assign _3131_ = ~(_3129_ | _3130_);
	assign _3628_[12] = _3131_ ^ \mchip.game2.scroll_inst.tick_time [12];
	assign _3132_ = _3131_ & ~\mchip.game2.scroll_inst.tick_time [12];
	assign _3628_[13] = _3132_ ^ \mchip.game2.scroll_inst.tick_time [13];
	assign _3133_ = ~(\mchip.game2.scroll_inst.tick_time [12] | \mchip.game2.scroll_inst.tick_time [13]);
	assign _3134_ = _3133_ & _3131_;
	assign _3628_[14] = _3134_ ^ \mchip.game2.scroll_inst.tick_time [14];
	assign _3135_ = _3134_ & ~\mchip.game2.scroll_inst.tick_time [14];
	assign _3628_[15] = _3135_ ^ \mchip.game2.scroll_inst.tick_time [15];
	assign _3136_ = \mchip.game2.scroll_inst.tick_time [14] | \mchip.game2.scroll_inst.tick_time [15];
	assign _3137_ = _3133_ & ~_3136_;
	assign _3138_ = _3136_ | ~_3133_;
	assign _3139_ = _3129_ & ~_3138_;
	assign _3140_ = _3137_ & ~_3139_;
	assign _3141_ = _3138_ | _3129_;
	assign _3142_ = _3123_ & ~_3141_;
	assign _3143_ = _3140_ & ~_3142_;
	assign _3628_[16] = _3143_ ^ \mchip.game2.scroll_inst.tick_time [16];
	assign _3144_ = _3143_ & ~\mchip.game2.scroll_inst.tick_time [16];
	assign _3628_[17] = _3144_ ^ \mchip.game2.scroll_inst.tick_time [17];
	assign _3145_ = io_in[3] & io_in[11];
	assign _3146_ = _3145_ & \mchip.game2.scroll_inst.pos [0];
	assign _3147_ = io_in[11] & ~io_in[4];
	assign _3148_ = _3147_ ^ \mchip.game2.scroll_inst.pos [1];
	assign _3627_[1] = ~(_3148_ ^ _3146_);
	assign _3149_ = _3146_ & ~_3148_;
	assign _3150_ = \mchip.game2.scroll_inst.pos [1] & ~_3147_;
	assign _3151_ = _3150_ | _3149_;
	assign _3152_ = io_in[5] & io_in[11];
	assign _3153_ = _3152_ ^ \mchip.game2.scroll_inst.pos [2];
	assign _3627_[2] = _3153_ ^ _3151_;
	assign _3154_ = _3152_ & \mchip.game2.scroll_inst.pos [2];
	assign _3155_ = _3153_ & _3151_;
	assign _3156_ = _3155_ | _3154_;
	assign _3157_ = io_in[6] & io_in[11];
	assign _3158_ = _3157_ ^ \mchip.game2.scroll_inst.pos [3];
	assign _3627_[3] = _3158_ ^ _3156_;
	assign _3159_ = ~(_3157_ & \mchip.game2.scroll_inst.pos [3]);
	assign _3160_ = _3158_ & _3154_;
	assign _3161_ = _3159_ & ~_3160_;
	assign _3162_ = ~(_3158_ & _3153_);
	assign _3163_ = _3151_ & ~_3162_;
	assign _3164_ = _3161_ & ~_3163_;
	assign _3627_[4] = ~(_3164_ ^ \mchip.game2.scroll_inst.pos [4]);
	assign _3165_ = \mchip.game2.scroll_inst.pos [4] & ~_3164_;
	assign _3627_[5] = _3165_ ^ \mchip.game2.scroll_inst.pos [5];
	assign _3166_ = ~(_3164_ | _0327_);
	assign _3627_[6] = _3166_ ^ \mchip.game2.scroll_inst.pos [6];
	assign _3167_ = _3166_ & \mchip.game2.scroll_inst.pos [6];
	assign _3627_[7] = _3167_ ^ \mchip.game2.scroll_inst.pos [7];
	assign _3168_ = _0328_ & ~_3164_;
	assign _3627_[8] = _3168_ ^ \mchip.game2.scroll_inst.pos [8];
	assign _3169_ = _3168_ & \mchip.game2.scroll_inst.pos [8];
	assign _3627_[9] = _3169_ ^ \mchip.game2.scroll_inst.pos [9];
	assign _3170_ = _3168_ & ~_0378_;
	assign _3627_[10] = _3170_ ^ \mchip.game2.scroll_inst.pos [10];
	assign _3626_[0] = _3145_ ^ \mchip.game2.scroll_inst.pos [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.hsync  <= 1'h1;
		else
			\mchip.game2.vga_inst.hsync  <= _0150_;
	always @(posedge io_in[12])
		if (_0016_)
			\mchip.game2.rendering_inst.layers [4] <= 1'h0;
		else
			\mchip.game2.rendering_inst.layers [4] <= _0021_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.game2.rendering_inst.layers [1] <= 1'h0;
		else
			\mchip.game2.rendering_inst.layers [1] <= _0022_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.game_over  <= 1'h1;
		else if (_0001_)
			\mchip.game2.game_over  <= _0027_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.cactus_type [2] <= 1'h0;
		else if (_0024_)
			\mchip.game2.cactus_type [2] <= \mchip.game2.rng_inst.out [4];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [0] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [0] <= _3622_[0];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [1] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [1] <= _3624_[1];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [2] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [2] <= _3624_[2];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [3] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [3] <= _3624_[3];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [4] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [4] <= _3624_[4];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [5] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [5] <= _3624_[5];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [6] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [6] <= _3624_[6];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [7] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [7] <= _3624_[7];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [8] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [8] <= _3624_[8];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [9] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [9] <= _3624_[9];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [10] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [10] <= _3624_[10];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [11] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [11] <= _3624_[11];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [12] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [12] <= _3624_[12];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [13] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [13] <= _3624_[13];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [14] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [14] <= _3624_[14];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [15] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [15] <= _3624_[15];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [16] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [16] <= _3624_[16];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [17] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [17] <= _3624_[17];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [18] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [18] <= _3624_[18];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [19] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [19] <= _3624_[19];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [20] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [20] <= _3624_[20];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [21] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [21] <= _3624_[21];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [22] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [22] <= _3624_[22];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [23] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [23] <= _3624_[23];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [24] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [24] <= _3624_[24];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [25] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [25] <= _3624_[25];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [26] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [26] <= _3624_[26];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [27] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [27] <= _3624_[27];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [28] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [28] <= _3624_[28];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [29] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [29] <= _3624_[29];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [30] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [30] <= _3624_[30];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.start_ctr [31] <= 1'h0;
		else if (_0162_)
			\mchip.game2.start_ctr [31] <= _3624_[31];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.cactus_select_last [0] <= 1'h0;
		else
			\mchip.game2.cactus_select_last [0] <= \mchip.game2.rendering_inst.cactus_select [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.cactus_select_last [1] <= 1'h0;
		else
			\mchip.game2.cactus_select_last [1] <= \mchip.game2.rendering_inst.cactus_select [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.cactus_select_last [2] <= 1'h0;
		else
			\mchip.game2.cactus_select_last [2] <= \mchip.game2.rendering_inst.cactus_select [2];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.in_air  <= 1'h0;
		else if (_0163_)
			\mchip.game2.jumping_inst.in_air  <= _0054_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.frame [0] <= 1'h0;
		else if (_0010_)
			\mchip.game2.jumping_inst.frame [0] <= _0055_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.frame [1] <= 1'h0;
		else if (_0010_)
			\mchip.game2.jumping_inst.frame [1] <= _0056_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.frame [2] <= 1'h0;
		else if (_0010_)
			\mchip.game2.jumping_inst.frame [2] <= _0057_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.frame [3] <= 1'h0;
		else if (_0010_)
			\mchip.game2.jumping_inst.frame [3] <= _0058_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.frame [4] <= 1'h0;
		else if (_0010_)
			\mchip.game2.jumping_inst.frame [4] <= _0059_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.frame [5] <= 1'h0;
		else if (_0010_)
			\mchip.game2.jumping_inst.frame [5] <= _0060_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.frame [6] <= 1'h0;
		else if (_0010_)
			\mchip.game2.jumping_inst.frame [6] <= _0061_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.frame [7] <= 1'h0;
		else if (_0010_)
			\mchip.game2.jumping_inst.frame [7] <= _0062_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.frame [8] <= 1'h0;
		else if (_0010_)
			\mchip.game2.jumping_inst.frame [8] <= _0063_;
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [0] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [0] <= _3621_[0];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [1] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [1] <= _3623_[1];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [2] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [2] <= _3623_[2];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [3] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [3] <= _3623_[3];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [4] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [4] <= _3623_[4];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [5] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [5] <= _3623_[5];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [6] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [6] <= _3623_[6];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [7] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [7] <= _3623_[7];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [8] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [8] <= _3623_[8];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [9] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [9] <= _3623_[9];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [10] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [10] <= _3623_[10];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [11] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [11] <= _3623_[11];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [12] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [12] <= _3623_[12];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [13] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [13] <= _3623_[13];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [14] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [14] <= _3623_[14];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [15] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [15] <= _3623_[15];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [16] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [16] <= _3623_[16];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [17] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [17] <= _3623_[17];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [18] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [18] <= _3623_[18];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.game2.no_jump_ctr [19] <= 1'h0;
		else
			\mchip.game2.no_jump_ctr [19] <= _3623_[19];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [0] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [0] <= _0064_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [1] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [1] <= _0075_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [2] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [2] <= _0080_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [3] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [3] <= _0081_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [4] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [4] <= _0082_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [5] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [5] <= _0083_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [6] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [6] <= _0084_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [7] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [7] <= _0085_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [8] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [8] <= _0086_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [9] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [9] <= _0087_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [10] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [10] <= _0065_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [11] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [11] <= _0066_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [12] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [12] <= _0067_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [13] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [13] <= _0068_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [14] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [14] <= _0069_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [15] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [15] <= _0070_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [16] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [16] <= _0071_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [17] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [17] <= _0072_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [18] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [18] <= _0073_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [19] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [19] <= _0074_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [20] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [20] <= _0076_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [21] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [21] <= _0077_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [22] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [22] <= _0078_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.jumping_inst.ctr [23] <= 1'h0;
		else if (_0011_)
			\mchip.game2.jumping_inst.ctr [23] <= _0079_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [0] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [0] <= _0029_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [1] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [1] <= _0040_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [2] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [2] <= _0046_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [3] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [3] <= _0047_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [4] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [4] <= _0048_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [5] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [5] <= _0049_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [6] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [6] <= _0050_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [7] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [7] <= _0051_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [8] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [8] <= _0052_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [9] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [9] <= _0053_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [10] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [10] <= _0030_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [11] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [11] <= _0031_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [12] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [12] <= _0032_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [13] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [13] <= _0033_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [14] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [14] <= _0034_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [15] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [15] <= _0035_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [16] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [16] <= _0036_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [17] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [17] <= _0037_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [18] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [18] <= _0038_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [19] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [19] <= _0039_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [20] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [20] <= _0041_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [21] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [21] <= _0042_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [22] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [22] <= _0043_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [23] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [23] <= _0044_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.ctr [24] <= 1'h0;
		else if (_0163_)
			\mchip.game2.dinosprite_inst.ctr [24] <= _0045_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.dinosprite_inst.sprite  <= 1'h0;
		else if (_0012_)
			\mchip.game2.dinosprite_inst.sprite  <= _0028_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [0] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [0] <= _3628_[0];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [1] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [1] <= _3628_[1];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [2] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [2] <= _3628_[2];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [3] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [3] <= _3628_[3];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [4] <= 1'h1;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [4] <= _3628_[4];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [5] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [5] <= _3628_[5];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [6] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [6] <= _3628_[6];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [7] <= 1'h1;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [7] <= _3628_[7];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [8] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [8] <= _3628_[8];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [9] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [9] <= _3628_[9];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [10] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [10] <= _3628_[10];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [11] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [11] <= _3628_[11];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [12] <= 1'h1;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [12] <= _3628_[12];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [13] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [13] <= _3628_[13];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [14] <= 1'h1;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [14] <= _3628_[14];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [15] <= 1'h1;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [15] <= _3628_[15];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [16] <= 1'h1;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [16] <= _3628_[16];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.tick_time [17] <= 1'h1;
		else if (_0002_)
			\mchip.game2.scroll_inst.tick_time [17] <= _3628_[17];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [0] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [0] <= _3626_[0];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [1] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [1] <= _3627_[1];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [2] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [2] <= _3627_[2];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [3] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [3] <= _3627_[3];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [4] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [4] <= _3627_[4];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [5] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [5] <= _3627_[5];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [6] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [6] <= _3627_[6];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [7] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [7] <= _3627_[7];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [8] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [8] <= _3627_[8];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [9] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [9] <= _3627_[9];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.pos [10] <= 1'h0;
		else if (_0002_)
			\mchip.game2.scroll_inst.pos [10] <= _3627_[10];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [0] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [0] <= _0132_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [1] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [1] <= _0141_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [2] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [2] <= _0142_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [3] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [3] <= _0143_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [4] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [4] <= _0144_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [5] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [5] <= _0145_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [6] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [6] <= _0146_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [7] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [7] <= _0147_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [8] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [8] <= _0148_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [9] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [9] <= _0149_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [10] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [10] <= _0133_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [11] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [11] <= _0134_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [12] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [12] <= _0135_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [13] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [13] <= _0136_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [14] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [14] <= _0137_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [15] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [15] <= _0138_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [16] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [16] <= _0139_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.scroll_inst.ctr [17] <= 1'h0;
		else if (_0163_)
			\mchip.game2.scroll_inst.ctr [17] <= _0140_;
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [0] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [0] <= _3620_[0];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [1] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [1] <= _3625_[1];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [2] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [2] <= _3625_[2];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [3] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [3] <= _3625_[3];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [4] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [4] <= _3625_[4];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [5] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [5] <= _3625_[5];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [6] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [6] <= _3625_[6];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [7] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [7] <= _3625_[7];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [8] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [8] <= _3625_[8];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.game2.vga_inst.haddr [9] <= 1'h0;
		else
			\mchip.game2.vga_inst.haddr [9] <= _3625_[9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vsync  <= 1'h1;
		else if (_0023_)
			\mchip.game2.vga_inst.vsync  <= _0151_;
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[3] [0] <= \mchip.game2.score_inst.score[3] [0];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[3] [1] <= \mchip.game2.score_inst.score[3] [1];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[3] [2] <= \mchip.game2.score_inst.score[3] [2];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[3] [3] <= \mchip.game2.score_inst.score[3] [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [0] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [0] <= _0152_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [1] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [1] <= _0153_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [2] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [2] <= _0154_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [3] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [3] <= _0155_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [4] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [4] <= _0156_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [5] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [5] <= _0157_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [6] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [6] <= _0158_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [7] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [7] <= _0159_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [8] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [8] <= _0160_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.vga_inst.vaddr [9] <= 1'h0;
		else if (_0023_)
			\mchip.game2.vga_inst.vaddr [9] <= _0161_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.rng_inst.out [0] <= 1'h1;
		else if (io_in[0])
			\mchip.game2.rng_inst.out [0] <= _0091_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.rng_inst.out [1] <= 1'h0;
		else if (io_in[0])
			\mchip.game2.rng_inst.out [1] <= \mchip.game2.rng_inst.out [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.rng_inst.out [2] <= 1'h0;
		else if (io_in[0])
			\mchip.game2.rng_inst.out [2] <= \mchip.game2.rng_inst.out [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.rng_inst.out [3] <= 1'h0;
		else if (io_in[0])
			\mchip.game2.rng_inst.out [3] <= \mchip.game2.rng_inst.out [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.rng_inst.out [4] <= 1'h0;
		else if (io_in[0])
			\mchip.game2.rng_inst.out [4] <= \mchip.game2.rng_inst.out [3];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[3] [0] <= 1'h0;
		else if (_0003_)
			\mchip.game2.score_inst.score[3] [0] <= _0094_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[3] [1] <= 1'h0;
		else if (_0003_)
			\mchip.game2.score_inst.score[3] [1] <= _0095_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[3] [2] <= 1'h0;
		else if (_0003_)
			\mchip.game2.score_inst.score[3] [2] <= _0096_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[3] [3] <= 1'h0;
		else if (_0003_)
			\mchip.game2.score_inst.score[3] [3] <= _0097_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[2] [0] <= 1'h0;
		else if (_0004_)
			\mchip.game2.score_inst.score[2] [0] <= _0098_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[2] [1] <= 1'h0;
		else if (_0004_)
			\mchip.game2.score_inst.score[2] [1] <= _0099_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[2] [2] <= 1'h0;
		else if (_0004_)
			\mchip.game2.score_inst.score[2] [2] <= _0100_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[2] [3] <= 1'h0;
		else if (_0004_)
			\mchip.game2.score_inst.score[2] [3] <= _0101_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[1] [0] <= 1'h0;
		else if (_0005_)
			\mchip.game2.score_inst.score[1] [0] <= _0102_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[1] [1] <= 1'h0;
		else if (_0005_)
			\mchip.game2.score_inst.score[1] [1] <= _0103_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[1] [2] <= 1'h0;
		else if (_0005_)
			\mchip.game2.score_inst.score[1] [2] <= _0104_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[1] [3] <= 1'h0;
		else if (_0005_)
			\mchip.game2.score_inst.score[1] [3] <= _0105_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[0] [0] <= 1'h0;
		else if (_0006_)
			\mchip.game2.score_inst.score[0] [0] <= _0106_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[0] [1] <= 1'h0;
		else if (_0006_)
			\mchip.game2.score_inst.score[0] [1] <= _0107_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[0] [2] <= 1'h0;
		else if (_0006_)
			\mchip.game2.score_inst.score[0] [2] <= _0108_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.score[0] [3] <= 1'h0;
		else if (_0006_)
			\mchip.game2.score_inst.score[0] [3] <= _0109_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [0] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [0] <= _0110_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [1] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [1] <= _0121_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [2] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [2] <= _0124_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [3] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [3] <= _0125_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [4] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [4] <= _0126_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [5] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [5] <= _0127_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [6] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [6] <= _0128_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [7] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [7] <= _0129_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [8] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [8] <= _0130_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [9] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [9] <= _0131_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [10] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [10] <= _0111_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [11] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [11] <= _0112_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [12] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [12] <= _0113_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [13] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [13] <= _0114_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [14] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [14] <= _0115_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [15] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [15] <= _0116_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [16] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [16] <= _0117_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [17] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [17] <= _0118_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [18] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [18] <= _0119_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [19] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [19] <= _0120_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [20] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [20] <= _0122_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.game2.score_inst.ctr [21] <= 1'h0;
		else if (_0163_)
			\mchip.game2.score_inst.ctr [21] <= _0123_;
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[2] [0] <= \mchip.game2.score_inst.score[2] [0];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[2] [1] <= \mchip.game2.score_inst.score[2] [1];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[2] [2] <= \mchip.game2.score_inst.score[2] [2];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[2] [3] <= \mchip.game2.score_inst.score[2] [3];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[1] [0] <= \mchip.game2.score_inst.score[1] [0];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[1] [1] <= \mchip.game2.score_inst.score[1] [1];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[1] [2] <= \mchip.game2.score_inst.score[1] [2];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[1] [3] <= \mchip.game2.score_inst.score[1] [3];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[0] [0] <= \mchip.game2.score_inst.score[0] [0];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[0] [1] <= \mchip.game2.score_inst.score[0] [1];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[0] [2] <= \mchip.game2.score_inst.score[0] [2];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.score_saved[0] [3] <= \mchip.game2.score_inst.score[0] [3];
	always @(posedge io_in[12])
		if (!_0092_)
			\mchip.game2.score_inst.pixel  <= 1'h0;
		else
			\mchip.game2.score_inst.pixel  <= _0093_;
	always @(posedge io_in[12])
		if (_0014_)
			\mchip.game2.rendering_inst.layers [3] <= 1'h0;
		else
			\mchip.game2.rendering_inst.layers [3] <= _3631_;
	always @(posedge io_in[12])
		if (_0017_)
			\mchip.game2.rendering_inst.layers [2] <= 1'h0;
		else
			\mchip.game2.rendering_inst.layers [2] <= _3630_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.rendering_inst.cactus_select [1] <= 1'h0;
		else if (_0008_)
			\mchip.game2.rendering_inst.cactus_select [1] <= _0089_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.rendering_inst.cactus_select [2] <= 1'h0;
		else if (_0007_)
			\mchip.game2.rendering_inst.cactus_select [2] <= _0090_;
	always @(posedge io_in[12])
		if (!_0020_)
			\mchip.game2.jumping_inst.jump_pos [0] <= _0000_[0];
	always @(posedge io_in[12])
		if (!_0020_)
			\mchip.game2.jumping_inst.jump_pos [1] <= _0000_[1];
	always @(posedge io_in[12])
		if (!_0020_)
			\mchip.game2.jumping_inst.jump_pos [2] <= _0000_[2];
	always @(posedge io_in[12])
		if (!_0020_)
			\mchip.game2.jumping_inst.jump_pos [3] <= _0000_[3];
	always @(posedge io_in[12])
		if (!_0020_)
			\mchip.game2.jumping_inst.jump_pos [4] <= _0000_[4];
	always @(posedge io_in[12])
		if (!_0020_)
			\mchip.game2.jumping_inst.jump_pos [5] <= _0000_[5];
	always @(posedge io_in[12])
		if (!_0020_)
			\mchip.game2.jumping_inst.jump_pos [6] <= _0000_[6];
	always @(posedge io_in[12])
		if (_0018_)
			\mchip.game2.rendering_inst.layers [0] <= 1'h0;
		else
			\mchip.game2.rendering_inst.layers [0] <= _3629_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.rendering_inst.cactus_select [0] <= 1'h0;
		else if (_0009_)
			\mchip.game2.rendering_inst.cactus_select [0] <= _0088_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.cactus_type [1] <= 1'h0;
		else if (_0025_)
			\mchip.game2.cactus_type [1] <= \mchip.game2.rng_inst.out [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.game2.cactus_type [0] <= 1'h0;
		else if (_0026_)
			\mchip.game2.cactus_type [0] <= \mchip.game2.rng_inst.out [2];
	assign _3620_[9:1] = 9'h000;
	assign _3621_[19:1] = 19'h00000;
	assign _3622_[31:1] = 31'h00000000;
	assign _3623_[0] = _3621_[0];
	assign _3624_[0] = _3622_[0];
	assign _3625_[0] = _3620_[0];
	assign _3626_[10:1] = {\mchip.game2.scroll_inst.pos [10:4], 3'h0};
	assign _3627_[0] = _3626_[0];
	assign io_out = {8'h00, \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.vga_inst.vsync , \mchip.game2.vga_inst.hsync };
	assign \mchip.clock  = io_in[12];
	assign \mchip.game2.cactus_select  = \mchip.game2.rendering_inst.cactus_select ;
	assign \mchip.game2.clk  = io_in[12];
	assign \mchip.game2.dbg_score  = {\mchip.game2.score_inst.score[3] , \mchip.game2.score_inst.score[2] , \mchip.game2.score_inst.score[1] , \mchip.game2.score_inst.score[0] };
	assign \mchip.game2.dbg_scrolladdr  = \mchip.game2.scroll_inst.pos ;
	assign \mchip.game2.dbg_speed  = {6'h00, \mchip.game2.scroll_inst.tick_time };
	assign \mchip.game2.debug_in  = io_in[2];
	assign \mchip.game2.dinosprite_inst.clk  = io_in[12];
	assign \mchip.game2.dinosprite_inst.sys_rst  = io_in[13];
	assign \mchip.game2.dinosprite_num  = \mchip.game2.dinosprite_inst.sprite ;
	assign \mchip.game2.haddr  = \mchip.game2.vga_inst.haddr ;
	assign \mchip.game2.halt_in  = io_in[1];
	assign \mchip.game2.jump_in  = io_in[0];
	assign \mchip.game2.jump_pos  = \mchip.game2.jumping_inst.jump_pos ;
	assign \mchip.game2.jumping_inst.clk  = io_in[12];
	assign \mchip.game2.jumping_inst.jump  = io_in[0];
	assign \mchip.game2.jumping_inst.speed  = 24'h03d090;
	assign \mchip.game2.jumping_inst.sys_rst  = io_in[13];
	assign \mchip.game2.random  = \mchip.game2.rng_inst.out ;
	assign \mchip.game2.rendering_inst.cactus_type  = \mchip.game2.cactus_type ;
	assign \mchip.game2.rendering_inst.clk  = io_in[12];
	assign \mchip.game2.rendering_inst.dinosprite_num  = \mchip.game2.dinosprite_inst.sprite ;
	assign \mchip.game2.rendering_inst.game_over  = \mchip.game2.game_over ;
	assign \mchip.game2.rendering_inst.haddr  = \mchip.game2.vga_inst.haddr ;
	assign \mchip.game2.rendering_inst.jump_pos  = \mchip.game2.jumping_inst.jump_pos ;
	assign \mchip.game2.rendering_inst.pixel  = \mchip.game2.dbg_pixel ;
	assign \mchip.game2.rendering_inst.score_pixel  = \mchip.game2.score_inst.pixel ;
	assign \mchip.game2.rendering_inst.scrolladdr  = \mchip.game2.scroll_inst.pos ;
	assign \mchip.game2.rendering_inst.sys_rst  = io_in[13];
	assign \mchip.game2.rendering_inst.vaddr  = \mchip.game2.vga_inst.vaddr ;
	assign \mchip.game2.rng_inst.clk  = io_in[12];
	assign \mchip.game2.rng_inst.entropy_in  = io_in[0];
	assign \mchip.game2.rng_inst.sys_rst  = io_in[13];
	assign \mchip.game2.score_inst.clk  = io_in[12];
	assign \mchip.game2.score_inst.haddr  = \mchip.game2.vga_inst.haddr ;
	assign \mchip.game2.score_inst.score_out  = {\mchip.game2.score_inst.score[3] , \mchip.game2.score_inst.score[2] , \mchip.game2.score_inst.score[1] , \mchip.game2.score_inst.score[0] };
	assign \mchip.game2.score_inst.sys_rst  = io_in[13];
	assign \mchip.game2.score_inst.vaddr  = \mchip.game2.vga_inst.vaddr ;
	assign \mchip.game2.score_out  = {\mchip.game2.score_inst.score[3] , \mchip.game2.score_inst.score[2] , \mchip.game2.score_inst.score[1] , \mchip.game2.score_inst.score[0] };
	assign \mchip.game2.score_pixel  = \mchip.game2.score_inst.pixel ;
	assign \mchip.game2.scroll_inst.clk  = io_in[12];
	assign \mchip.game2.scroll_inst.move_amt  = 8'h00;
	assign \mchip.game2.scroll_inst.speed  = {6'h00, \mchip.game2.scroll_inst.tick_time };
	assign \mchip.game2.scroll_inst.speed_change  = 8'h00;
	assign \mchip.game2.scroll_inst.sys_rst  = io_in[13];
	assign \mchip.game2.scrolladdr  = \mchip.game2.scroll_inst.pos ;
	assign \mchip.game2.speed  = {6'h00, \mchip.game2.scroll_inst.tick_time };
	assign \mchip.game2.sys_rst  = io_in[13];
	assign \mchip.game2.vaddr  = \mchip.game2.vga_inst.vaddr ;
	assign \mchip.game2.vga_blue  = {\mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel };
	assign \mchip.game2.vga_green  = {\mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel };
	assign \mchip.game2.vga_hsync  = \mchip.game2.vga_inst.hsync ;
	assign \mchip.game2.vga_inst.clk  = io_in[12];
	assign \mchip.game2.vga_inst.sys_rst  = io_in[13];
	assign \mchip.game2.vga_pixel  = \mchip.game2.dbg_pixel ;
	assign \mchip.game2.vga_red  = {\mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel };
	assign \mchip.game2.vga_vsync  = \mchip.game2.vga_inst.vsync ;
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {6'h00, \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.dbg_pixel , \mchip.game2.vga_inst.vsync , \mchip.game2.vga_inst.hsync };
	assign \mchip.reset  = io_in[13];
endmodule
module d10_jjalacce_connect4 (
	io_in,
	io_out
);
	wire _00000_;
	wire _00001_;
	wire _00002_;
	wire _00003_;
	wire _00004_;
	wire _00005_;
	wire _00006_;
	wire _00007_;
	wire _00008_;
	wire _00009_;
	wire _00010_;
	wire _00011_;
	wire _00012_;
	wire _00013_;
	wire _00014_;
	wire _00015_;
	wire _00016_;
	wire _00017_;
	wire _00018_;
	wire _00019_;
	wire _00020_;
	wire _00021_;
	wire _00022_;
	wire _00023_;
	wire _00024_;
	wire _00025_;
	wire _00026_;
	wire _00027_;
	wire _00028_;
	wire _00029_;
	wire _00030_;
	wire _00031_;
	wire _00032_;
	wire _00033_;
	wire _00034_;
	wire _00035_;
	wire _00036_;
	wire _00037_;
	wire _00038_;
	wire _00039_;
	wire _00040_;
	wire _00041_;
	wire _00042_;
	wire _00043_;
	wire _00044_;
	wire _00045_;
	wire _00046_;
	wire _00047_;
	wire _00048_;
	wire _00049_;
	wire _00050_;
	wire _00051_;
	wire _00052_;
	wire _00053_;
	wire _00054_;
	wire _00055_;
	wire _00056_;
	wire _00057_;
	wire _00058_;
	wire _00059_;
	wire _00060_;
	wire _00061_;
	wire _00062_;
	wire _00063_;
	wire _00064_;
	wire _00065_;
	wire _00066_;
	wire _00067_;
	wire _00068_;
	wire _00069_;
	wire _00070_;
	wire _00071_;
	wire _00072_;
	wire _00073_;
	wire _00074_;
	wire _00075_;
	wire _00076_;
	wire _00077_;
	wire _00078_;
	wire _00079_;
	wire _00080_;
	wire _00081_;
	wire _00082_;
	wire _00083_;
	wire _00084_;
	wire _00085_;
	wire _00086_;
	wire _00087_;
	wire _00088_;
	wire _00089_;
	wire _00090_;
	wire _00091_;
	wire _00092_;
	wire _00093_;
	wire _00094_;
	wire _00095_;
	wire _00096_;
	wire _00097_;
	wire _00098_;
	wire _00099_;
	wire _00100_;
	wire _00101_;
	wire _00102_;
	wire _00103_;
	wire _00104_;
	wire _00105_;
	wire _00106_;
	wire _00107_;
	wire _00108_;
	wire _00109_;
	wire _00110_;
	wire _00111_;
	wire _00112_;
	wire _00113_;
	wire _00114_;
	wire _00115_;
	wire _00116_;
	wire _00117_;
	wire _00118_;
	wire _00119_;
	wire _00120_;
	wire _00121_;
	wire _00122_;
	wire _00123_;
	wire _00124_;
	wire _00125_;
	wire _00126_;
	wire _00127_;
	wire _00128_;
	wire _00129_;
	wire _00130_;
	wire _00131_;
	wire _00132_;
	wire _00133_;
	wire _00134_;
	wire _00135_;
	wire _00136_;
	wire _00137_;
	wire _00138_;
	wire _00139_;
	wire _00140_;
	wire _00141_;
	wire _00142_;
	wire _00143_;
	wire _00144_;
	wire _00145_;
	wire _00146_;
	wire _00147_;
	wire _00148_;
	wire _00149_;
	wire _00150_;
	wire _00151_;
	wire _00152_;
	wire _00153_;
	wire _00154_;
	wire _00155_;
	wire _00156_;
	wire _00157_;
	wire _00158_;
	wire _00159_;
	wire _00160_;
	wire _00161_;
	wire _00162_;
	wire _00163_;
	wire _00164_;
	wire _00165_;
	wire _00166_;
	wire _00167_;
	wire _00168_;
	wire _00169_;
	wire _00170_;
	wire _00171_;
	wire _00172_;
	wire _00173_;
	wire _00174_;
	wire _00175_;
	wire _00176_;
	wire _00177_;
	wire _00178_;
	wire _00179_;
	wire _00180_;
	wire _00181_;
	wire _00182_;
	wire _00183_;
	wire _00184_;
	wire _00185_;
	wire _00186_;
	wire _00187_;
	wire _00188_;
	wire _00189_;
	wire _00190_;
	wire _00191_;
	wire _00192_;
	wire _00193_;
	wire _00194_;
	wire _00195_;
	wire _00196_;
	wire _00197_;
	wire _00198_;
	wire _00199_;
	wire _00200_;
	wire _00201_;
	wire _00202_;
	wire _00203_;
	wire _00204_;
	wire _00205_;
	wire _00206_;
	wire _00207_;
	wire _00208_;
	wire _00209_;
	wire _00210_;
	wire _00211_;
	wire _00212_;
	wire _00213_;
	wire _00214_;
	wire _00215_;
	wire _00216_;
	wire _00217_;
	wire _00218_;
	wire _00219_;
	wire _00220_;
	wire _00221_;
	wire _00222_;
	wire _00223_;
	wire _00224_;
	wire _00225_;
	wire _00226_;
	wire _00227_;
	wire _00228_;
	wire _00229_;
	wire _00230_;
	wire _00231_;
	wire _00232_;
	wire _00233_;
	wire _00234_;
	wire _00235_;
	wire _00236_;
	wire _00237_;
	wire _00238_;
	wire _00239_;
	wire _00240_;
	wire _00241_;
	wire _00242_;
	wire _00243_;
	wire _00244_;
	wire _00245_;
	wire _00246_;
	wire _00247_;
	wire _00248_;
	wire _00249_;
	wire _00250_;
	wire _00251_;
	wire _00252_;
	wire _00253_;
	wire _00254_;
	wire _00255_;
	wire _00256_;
	wire _00257_;
	wire _00258_;
	wire _00259_;
	wire _00260_;
	wire _00261_;
	wire _00262_;
	wire _00263_;
	wire _00264_;
	wire _00265_;
	wire _00266_;
	wire _00267_;
	wire _00268_;
	wire _00269_;
	wire _00270_;
	wire _00271_;
	wire _00272_;
	wire _00273_;
	wire _00274_;
	wire _00275_;
	wire _00276_;
	wire _00277_;
	wire _00278_;
	wire _00279_;
	wire _00280_;
	wire _00281_;
	wire _00282_;
	wire _00283_;
	wire _00284_;
	wire _00285_;
	wire _00286_;
	wire _00287_;
	wire _00288_;
	wire _00289_;
	wire _00290_;
	wire _00291_;
	wire _00292_;
	wire _00293_;
	wire _00294_;
	wire _00295_;
	wire _00296_;
	wire _00297_;
	wire _00298_;
	wire _00299_;
	wire _00300_;
	wire _00301_;
	wire _00302_;
	wire _00303_;
	wire _00304_;
	wire _00305_;
	wire _00306_;
	wire _00307_;
	wire _00308_;
	wire _00309_;
	wire _00310_;
	wire _00311_;
	wire _00312_;
	wire _00313_;
	wire _00314_;
	wire _00315_;
	wire _00316_;
	wire _00317_;
	wire _00318_;
	wire _00319_;
	wire _00320_;
	wire _00321_;
	wire _00322_;
	wire _00323_;
	wire _00324_;
	wire _00325_;
	wire _00326_;
	wire _00327_;
	wire _00328_;
	wire _00329_;
	wire _00330_;
	wire _00331_;
	wire _00332_;
	wire _00333_;
	wire _00334_;
	wire _00335_;
	wire _00336_;
	wire _00337_;
	wire _00338_;
	wire _00339_;
	wire _00340_;
	wire _00341_;
	wire _00342_;
	wire _00343_;
	wire _00344_;
	wire _00345_;
	wire _00346_;
	wire _00347_;
	wire _00348_;
	wire _00349_;
	wire _00350_;
	wire _00351_;
	wire _00352_;
	wire _00353_;
	wire _00354_;
	wire _00355_;
	wire _00356_;
	wire _00357_;
	wire _00358_;
	wire _00359_;
	wire _00360_;
	wire _00361_;
	wire _00362_;
	wire _00363_;
	wire _00364_;
	wire _00365_;
	wire _00366_;
	wire _00367_;
	wire _00368_;
	wire _00369_;
	wire _00370_;
	wire _00371_;
	wire _00372_;
	wire _00373_;
	wire _00374_;
	wire _00375_;
	wire _00376_;
	wire _00377_;
	wire _00378_;
	wire _00379_;
	wire _00380_;
	wire _00381_;
	wire _00382_;
	wire _00383_;
	wire _00384_;
	wire _00385_;
	wire _00386_;
	wire _00387_;
	wire _00388_;
	wire _00389_;
	wire _00390_;
	wire _00391_;
	wire _00392_;
	wire _00393_;
	wire _00394_;
	wire _00395_;
	wire _00396_;
	wire _00397_;
	wire _00398_;
	wire _00399_;
	wire _00400_;
	wire _00401_;
	wire _00402_;
	wire _00403_;
	wire _00404_;
	wire _00405_;
	wire _00406_;
	wire _00407_;
	wire _00408_;
	wire _00409_;
	wire _00410_;
	wire _00411_;
	wire _00412_;
	wire _00413_;
	wire _00414_;
	wire _00415_;
	wire _00416_;
	wire _00417_;
	wire _00418_;
	wire _00419_;
	wire _00420_;
	wire _00421_;
	wire _00422_;
	wire _00423_;
	wire _00424_;
	wire _00425_;
	wire _00426_;
	wire _00427_;
	wire _00428_;
	wire _00429_;
	wire _00430_;
	wire _00431_;
	wire _00432_;
	wire _00433_;
	wire _00434_;
	wire _00435_;
	wire _00436_;
	wire _00437_;
	wire _00438_;
	wire _00439_;
	wire _00440_;
	wire _00441_;
	wire _00442_;
	wire _00443_;
	wire _00444_;
	wire _00445_;
	wire _00446_;
	wire _00447_;
	wire _00448_;
	wire _00449_;
	wire _00450_;
	wire _00451_;
	wire _00452_;
	wire _00453_;
	wire _00454_;
	wire _00455_;
	wire _00456_;
	wire _00457_;
	wire _00458_;
	wire _00459_;
	wire _00460_;
	wire _00461_;
	wire _00462_;
	wire _00463_;
	wire _00464_;
	wire _00465_;
	wire _00466_;
	wire _00467_;
	wire _00468_;
	wire _00469_;
	wire _00470_;
	wire _00471_;
	wire _00472_;
	wire _00473_;
	wire _00474_;
	wire _00475_;
	wire _00476_;
	wire _00477_;
	wire _00478_;
	wire _00479_;
	wire _00480_;
	wire _00481_;
	wire _00482_;
	wire _00483_;
	wire _00484_;
	wire _00485_;
	wire _00486_;
	wire _00487_;
	wire _00488_;
	wire _00489_;
	wire _00490_;
	wire _00491_;
	wire _00492_;
	wire _00493_;
	wire _00494_;
	wire _00495_;
	wire _00496_;
	wire _00497_;
	wire _00498_;
	wire _00499_;
	wire _00500_;
	wire _00501_;
	wire _00502_;
	wire _00503_;
	wire _00504_;
	wire _00505_;
	wire _00506_;
	wire _00507_;
	wire _00508_;
	wire _00509_;
	wire _00510_;
	wire _00511_;
	wire _00512_;
	wire _00513_;
	wire _00514_;
	wire _00515_;
	wire _00516_;
	wire _00517_;
	wire _00518_;
	wire _00519_;
	wire _00520_;
	wire _00521_;
	wire _00522_;
	wire _00523_;
	wire _00524_;
	wire _00525_;
	wire _00526_;
	wire _00527_;
	wire _00528_;
	wire _00529_;
	wire _00530_;
	wire _00531_;
	wire _00532_;
	wire _00533_;
	wire _00534_;
	wire _00535_;
	wire _00536_;
	wire _00537_;
	wire _00538_;
	wire _00539_;
	wire _00540_;
	wire _00541_;
	wire _00542_;
	wire _00543_;
	wire _00544_;
	wire _00545_;
	wire _00546_;
	wire _00547_;
	wire _00548_;
	wire _00549_;
	wire _00550_;
	wire _00551_;
	wire _00552_;
	wire _00553_;
	wire _00554_;
	wire _00555_;
	wire _00556_;
	wire _00557_;
	wire _00558_;
	wire _00559_;
	wire _00560_;
	wire _00561_;
	wire _00562_;
	wire _00563_;
	wire _00564_;
	wire _00565_;
	wire _00566_;
	wire _00567_;
	wire _00568_;
	wire _00569_;
	wire _00570_;
	wire _00571_;
	wire _00572_;
	wire _00573_;
	wire _00574_;
	wire _00575_;
	wire _00576_;
	wire _00577_;
	wire _00578_;
	wire _00579_;
	wire _00580_;
	wire _00581_;
	wire _00582_;
	wire _00583_;
	wire _00584_;
	wire _00585_;
	wire _00586_;
	wire _00587_;
	wire _00588_;
	wire _00589_;
	wire _00590_;
	wire _00591_;
	wire _00592_;
	wire _00593_;
	wire _00594_;
	wire _00595_;
	wire _00596_;
	wire _00597_;
	wire _00598_;
	wire _00599_;
	wire _00600_;
	wire _00601_;
	wire _00602_;
	wire _00603_;
	wire _00604_;
	wire _00605_;
	wire _00606_;
	wire _00607_;
	wire _00608_;
	wire _00609_;
	wire _00610_;
	wire _00611_;
	wire _00612_;
	wire _00613_;
	wire _00614_;
	wire _00615_;
	wire _00616_;
	wire _00617_;
	wire _00618_;
	wire _00619_;
	wire _00620_;
	wire _00621_;
	wire _00622_;
	wire _00623_;
	wire _00624_;
	wire _00625_;
	wire _00626_;
	wire _00627_;
	wire _00628_;
	wire _00629_;
	wire _00630_;
	wire _00631_;
	wire _00632_;
	wire _00633_;
	wire _00634_;
	wire _00635_;
	wire _00636_;
	wire _00637_;
	wire _00638_;
	wire _00639_;
	wire _00640_;
	wire _00641_;
	wire _00642_;
	wire _00643_;
	wire _00644_;
	wire _00645_;
	wire _00646_;
	wire _00647_;
	wire _00648_;
	wire _00649_;
	wire _00650_;
	wire _00651_;
	wire _00652_;
	wire _00653_;
	wire _00654_;
	wire _00655_;
	wire _00656_;
	wire _00657_;
	wire _00658_;
	wire _00659_;
	wire _00660_;
	wire _00661_;
	wire _00662_;
	wire _00663_;
	wire _00664_;
	wire _00665_;
	wire _00666_;
	wire _00667_;
	wire _00668_;
	wire _00669_;
	wire _00670_;
	wire _00671_;
	wire _00672_;
	wire _00673_;
	wire _00674_;
	wire _00675_;
	wire _00676_;
	wire _00677_;
	wire _00678_;
	wire _00679_;
	wire _00680_;
	wire _00681_;
	wire _00682_;
	wire _00683_;
	wire _00684_;
	wire _00685_;
	wire _00686_;
	wire _00687_;
	wire _00688_;
	wire _00689_;
	wire _00690_;
	wire _00691_;
	wire _00692_;
	wire _00693_;
	wire _00694_;
	wire _00695_;
	wire _00696_;
	wire _00697_;
	wire _00698_;
	wire _00699_;
	wire _00700_;
	wire _00701_;
	wire _00702_;
	wire _00703_;
	wire _00704_;
	wire _00705_;
	wire _00706_;
	wire _00707_;
	wire _00708_;
	wire _00709_;
	wire _00710_;
	wire _00711_;
	wire _00712_;
	wire _00713_;
	wire _00714_;
	wire _00715_;
	wire _00716_;
	wire _00717_;
	wire _00718_;
	wire _00719_;
	wire _00720_;
	wire _00721_;
	wire _00722_;
	wire _00723_;
	wire _00724_;
	wire _00725_;
	wire _00726_;
	wire _00727_;
	wire _00728_;
	wire _00729_;
	wire _00730_;
	wire _00731_;
	wire _00732_;
	wire _00733_;
	wire _00734_;
	wire _00735_;
	wire _00736_;
	wire _00737_;
	wire _00738_;
	wire _00739_;
	wire _00740_;
	wire _00741_;
	wire _00742_;
	wire _00743_;
	wire _00744_;
	wire _00745_;
	wire _00746_;
	wire _00747_;
	wire _00748_;
	wire _00749_;
	wire _00750_;
	wire _00751_;
	wire _00752_;
	wire _00753_;
	wire _00754_;
	wire _00755_;
	wire _00756_;
	wire _00757_;
	wire _00758_;
	wire _00759_;
	wire _00760_;
	wire _00761_;
	wire _00762_;
	wire _00763_;
	wire _00764_;
	wire _00765_;
	wire _00766_;
	wire _00767_;
	wire _00768_;
	wire _00769_;
	wire _00770_;
	wire _00771_;
	wire _00772_;
	wire _00773_;
	wire _00774_;
	wire _00775_;
	wire _00776_;
	wire _00777_;
	wire _00778_;
	wire _00779_;
	wire _00780_;
	wire _00781_;
	wire _00782_;
	wire _00783_;
	wire _00784_;
	wire _00785_;
	wire _00786_;
	wire _00787_;
	wire _00788_;
	wire _00789_;
	wire _00790_;
	wire _00791_;
	wire _00792_;
	wire _00793_;
	wire _00794_;
	wire _00795_;
	wire _00796_;
	wire _00797_;
	wire _00798_;
	wire _00799_;
	wire _00800_;
	wire _00801_;
	wire _00802_;
	wire _00803_;
	wire _00804_;
	wire _00805_;
	wire _00806_;
	wire _00807_;
	wire _00808_;
	wire _00809_;
	wire _00810_;
	wire _00811_;
	wire _00812_;
	wire _00813_;
	wire _00814_;
	wire _00815_;
	wire _00816_;
	wire _00817_;
	wire _00818_;
	wire _00819_;
	wire _00820_;
	wire _00821_;
	wire _00822_;
	wire _00823_;
	wire _00824_;
	wire _00825_;
	wire _00826_;
	wire _00827_;
	wire _00828_;
	wire _00829_;
	wire _00830_;
	wire _00831_;
	wire _00832_;
	wire _00833_;
	wire _00834_;
	wire _00835_;
	wire _00836_;
	wire _00837_;
	wire _00838_;
	wire _00839_;
	wire _00840_;
	wire _00841_;
	wire _00842_;
	wire _00843_;
	wire _00844_;
	wire _00845_;
	wire _00846_;
	wire _00847_;
	wire _00848_;
	wire _00849_;
	wire _00850_;
	wire _00851_;
	wire _00852_;
	wire _00853_;
	wire _00854_;
	wire _00855_;
	wire _00856_;
	wire _00857_;
	wire _00858_;
	wire _00859_;
	wire _00860_;
	wire _00861_;
	wire _00862_;
	wire _00863_;
	wire _00864_;
	wire _00865_;
	wire _00866_;
	wire _00867_;
	wire _00868_;
	wire _00869_;
	wire _00870_;
	wire _00871_;
	wire _00872_;
	wire _00873_;
	wire _00874_;
	wire _00875_;
	wire _00876_;
	wire _00877_;
	wire _00878_;
	wire _00879_;
	wire _00880_;
	wire _00881_;
	wire _00882_;
	wire _00883_;
	wire _00884_;
	wire _00885_;
	wire _00886_;
	wire _00887_;
	wire _00888_;
	wire _00889_;
	wire _00890_;
	wire _00891_;
	wire _00892_;
	wire _00893_;
	wire _00894_;
	wire _00895_;
	wire _00896_;
	wire _00897_;
	wire _00898_;
	wire _00899_;
	wire _00900_;
	wire _00901_;
	wire _00902_;
	wire _00903_;
	wire _00904_;
	wire _00905_;
	wire _00906_;
	wire _00907_;
	wire _00908_;
	wire _00909_;
	wire _00910_;
	wire _00911_;
	wire _00912_;
	wire _00913_;
	wire _00914_;
	wire _00915_;
	wire _00916_;
	wire _00917_;
	wire _00918_;
	wire _00919_;
	wire _00920_;
	wire _00921_;
	wire _00922_;
	wire _00923_;
	wire _00924_;
	wire _00925_;
	wire _00926_;
	wire _00927_;
	wire _00928_;
	wire _00929_;
	wire _00930_;
	wire _00931_;
	wire _00932_;
	wire _00933_;
	wire _00934_;
	wire _00935_;
	wire _00936_;
	wire _00937_;
	wire _00938_;
	wire _00939_;
	wire _00940_;
	wire _00941_;
	wire _00942_;
	wire _00943_;
	wire _00944_;
	wire _00945_;
	wire _00946_;
	wire _00947_;
	wire _00948_;
	wire _00949_;
	wire _00950_;
	wire _00951_;
	wire _00952_;
	wire _00953_;
	wire _00954_;
	wire _00955_;
	wire _00956_;
	wire _00957_;
	wire _00958_;
	wire _00959_;
	wire _00960_;
	wire _00961_;
	wire _00962_;
	wire _00963_;
	wire _00964_;
	wire _00965_;
	wire _00966_;
	wire _00967_;
	wire _00968_;
	wire _00969_;
	wire _00970_;
	wire _00971_;
	wire _00972_;
	wire _00973_;
	wire _00974_;
	wire _00975_;
	wire _00976_;
	wire _00977_;
	wire _00978_;
	wire _00979_;
	wire _00980_;
	wire _00981_;
	wire _00982_;
	wire _00983_;
	wire _00984_;
	wire _00985_;
	wire _00986_;
	wire _00987_;
	wire _00988_;
	wire _00989_;
	wire _00990_;
	wire _00991_;
	wire _00992_;
	wire _00993_;
	wire _00994_;
	wire _00995_;
	wire _00996_;
	wire _00997_;
	wire _00998_;
	wire _00999_;
	wire _01000_;
	wire _01001_;
	wire _01002_;
	wire _01003_;
	wire _01004_;
	wire _01005_;
	wire _01006_;
	wire _01007_;
	wire _01008_;
	wire _01009_;
	wire _01010_;
	wire _01011_;
	wire _01012_;
	wire _01013_;
	wire _01014_;
	wire _01015_;
	wire _01016_;
	wire _01017_;
	wire _01018_;
	wire _01019_;
	wire _01020_;
	wire _01021_;
	wire _01022_;
	wire _01023_;
	wire _01024_;
	wire _01025_;
	wire _01026_;
	wire _01027_;
	wire _01028_;
	wire _01029_;
	wire _01030_;
	wire _01031_;
	wire _01032_;
	wire _01033_;
	wire _01034_;
	wire _01035_;
	wire _01036_;
	wire _01037_;
	wire _01038_;
	wire _01039_;
	wire _01040_;
	wire _01041_;
	wire _01042_;
	wire _01043_;
	wire _01044_;
	wire _01045_;
	wire _01046_;
	wire _01047_;
	wire _01048_;
	wire _01049_;
	wire _01050_;
	wire _01051_;
	wire _01052_;
	wire _01053_;
	wire _01054_;
	wire _01055_;
	wire _01056_;
	wire _01057_;
	wire _01058_;
	wire _01059_;
	wire _01060_;
	wire _01061_;
	wire _01062_;
	wire _01063_;
	wire _01064_;
	wire _01065_;
	wire _01066_;
	wire _01067_;
	wire _01068_;
	wire _01069_;
	wire _01070_;
	wire _01071_;
	wire _01072_;
	wire _01073_;
	wire _01074_;
	wire _01075_;
	wire _01076_;
	wire _01077_;
	wire _01078_;
	wire _01079_;
	wire _01080_;
	wire _01081_;
	wire _01082_;
	wire _01083_;
	wire _01084_;
	wire _01085_;
	wire _01086_;
	wire _01087_;
	wire _01088_;
	wire _01089_;
	wire _01090_;
	wire _01091_;
	wire _01092_;
	wire _01093_;
	wire _01094_;
	wire _01095_;
	wire _01096_;
	wire _01097_;
	wire _01098_;
	wire _01099_;
	wire _01100_;
	wire _01101_;
	wire _01102_;
	wire _01103_;
	wire _01104_;
	wire _01105_;
	wire _01106_;
	wire _01107_;
	wire _01108_;
	wire _01109_;
	wire _01110_;
	wire _01111_;
	wire _01112_;
	wire _01113_;
	wire _01114_;
	wire _01115_;
	wire _01116_;
	wire _01117_;
	wire _01118_;
	wire _01119_;
	wire _01120_;
	wire _01121_;
	wire _01122_;
	wire _01123_;
	wire _01124_;
	wire _01125_;
	wire _01126_;
	wire _01127_;
	wire _01128_;
	wire _01129_;
	wire _01130_;
	wire _01131_;
	wire _01132_;
	wire _01133_;
	wire _01134_;
	wire _01135_;
	wire _01136_;
	wire _01137_;
	wire _01138_;
	wire _01139_;
	wire _01140_;
	wire _01141_;
	wire _01142_;
	wire _01143_;
	wire _01144_;
	wire _01145_;
	wire _01146_;
	wire _01147_;
	wire _01148_;
	wire _01149_;
	wire _01150_;
	wire _01151_;
	wire _01152_;
	wire _01153_;
	wire _01154_;
	wire _01155_;
	wire _01156_;
	wire _01157_;
	wire _01158_;
	wire _01159_;
	wire _01160_;
	wire _01161_;
	wire _01162_;
	wire _01163_;
	wire _01164_;
	wire _01165_;
	wire _01166_;
	wire _01167_;
	wire _01168_;
	wire _01169_;
	wire _01170_;
	wire _01171_;
	wire _01172_;
	wire _01173_;
	wire _01174_;
	wire _01175_;
	wire _01176_;
	wire _01177_;
	wire _01178_;
	wire _01179_;
	wire _01180_;
	wire _01181_;
	wire _01182_;
	wire _01183_;
	wire _01184_;
	wire _01185_;
	wire _01186_;
	wire _01187_;
	wire _01188_;
	wire _01189_;
	wire _01190_;
	wire _01191_;
	wire _01192_;
	wire _01193_;
	wire _01194_;
	wire _01195_;
	wire _01196_;
	wire _01197_;
	wire _01198_;
	wire _01199_;
	wire _01200_;
	wire _01201_;
	wire _01202_;
	wire _01203_;
	wire _01204_;
	wire _01205_;
	wire _01206_;
	wire _01207_;
	wire _01208_;
	wire _01209_;
	wire _01210_;
	wire _01211_;
	wire _01212_;
	wire _01213_;
	wire _01214_;
	wire _01215_;
	wire _01216_;
	wire _01217_;
	wire _01218_;
	wire _01219_;
	wire _01220_;
	wire _01221_;
	wire _01222_;
	wire _01223_;
	wire _01224_;
	wire _01225_;
	wire _01226_;
	wire _01227_;
	wire _01228_;
	wire _01229_;
	wire _01230_;
	wire _01231_;
	wire _01232_;
	wire _01233_;
	wire _01234_;
	wire _01235_;
	wire _01236_;
	wire _01237_;
	wire _01238_;
	wire _01239_;
	wire _01240_;
	wire _01241_;
	wire _01242_;
	wire _01243_;
	wire _01244_;
	wire _01245_;
	wire _01246_;
	wire _01247_;
	wire _01248_;
	wire _01249_;
	wire _01250_;
	wire _01251_;
	wire _01252_;
	wire _01253_;
	wire _01254_;
	wire _01255_;
	wire _01256_;
	wire _01257_;
	wire _01258_;
	wire _01259_;
	wire _01260_;
	wire _01261_;
	wire _01262_;
	wire _01263_;
	wire _01264_;
	wire _01265_;
	wire _01266_;
	wire _01267_;
	wire _01268_;
	wire _01269_;
	wire _01270_;
	wire _01271_;
	wire _01272_;
	wire _01273_;
	wire _01274_;
	wire _01275_;
	wire _01276_;
	wire _01277_;
	wire _01278_;
	wire _01279_;
	wire _01280_;
	wire _01281_;
	wire _01282_;
	wire _01283_;
	wire _01284_;
	wire _01285_;
	wire _01286_;
	wire _01287_;
	wire _01288_;
	wire _01289_;
	wire _01290_;
	wire _01291_;
	wire _01292_;
	wire _01293_;
	wire _01294_;
	wire _01295_;
	wire _01296_;
	wire _01297_;
	wire _01298_;
	wire _01299_;
	wire _01300_;
	wire _01301_;
	wire _01302_;
	wire _01303_;
	wire _01304_;
	wire _01305_;
	wire _01306_;
	wire _01307_;
	wire _01308_;
	wire _01309_;
	wire _01310_;
	wire _01311_;
	wire _01312_;
	wire _01313_;
	wire _01314_;
	wire _01315_;
	wire _01316_;
	wire _01317_;
	wire _01318_;
	wire _01319_;
	wire _01320_;
	wire _01321_;
	wire _01322_;
	wire _01323_;
	wire _01324_;
	wire _01325_;
	wire _01326_;
	wire _01327_;
	wire _01328_;
	wire _01329_;
	wire _01330_;
	wire _01331_;
	wire _01332_;
	wire _01333_;
	wire _01334_;
	wire _01335_;
	wire _01336_;
	wire _01337_;
	wire _01338_;
	wire _01339_;
	wire _01340_;
	wire _01341_;
	wire _01342_;
	wire _01343_;
	wire _01344_;
	wire _01345_;
	wire _01346_;
	wire _01347_;
	wire _01348_;
	wire _01349_;
	wire _01350_;
	wire _01351_;
	wire _01352_;
	wire _01353_;
	wire _01354_;
	wire _01355_;
	wire _01356_;
	wire _01357_;
	wire _01358_;
	wire _01359_;
	wire _01360_;
	wire _01361_;
	wire _01362_;
	wire _01363_;
	wire _01364_;
	wire _01365_;
	wire _01366_;
	wire _01367_;
	wire _01368_;
	wire _01369_;
	wire _01370_;
	wire _01371_;
	wire _01372_;
	wire _01373_;
	wire _01374_;
	wire _01375_;
	wire _01376_;
	wire _01377_;
	wire _01378_;
	wire _01379_;
	wire _01380_;
	wire _01381_;
	wire _01382_;
	wire _01383_;
	wire _01384_;
	wire _01385_;
	wire _01386_;
	wire _01387_;
	wire _01388_;
	wire _01389_;
	wire _01390_;
	wire _01391_;
	wire _01392_;
	wire _01393_;
	wire _01394_;
	wire _01395_;
	wire _01396_;
	wire _01397_;
	wire _01398_;
	wire _01399_;
	wire _01400_;
	wire _01401_;
	wire _01402_;
	wire _01403_;
	wire _01404_;
	wire _01405_;
	wire _01406_;
	wire _01407_;
	wire _01408_;
	wire _01409_;
	wire _01410_;
	wire _01411_;
	wire _01412_;
	wire _01413_;
	wire _01414_;
	wire _01415_;
	wire _01416_;
	wire _01417_;
	wire _01418_;
	wire _01419_;
	wire _01420_;
	wire _01421_;
	wire _01422_;
	wire _01423_;
	wire _01424_;
	wire _01425_;
	wire _01426_;
	wire _01427_;
	wire _01428_;
	wire _01429_;
	wire _01430_;
	wire _01431_;
	wire _01432_;
	wire _01433_;
	wire _01434_;
	wire _01435_;
	wire _01436_;
	wire _01437_;
	wire _01438_;
	wire _01439_;
	wire _01440_;
	wire _01441_;
	wire _01442_;
	wire _01443_;
	wire _01444_;
	wire _01445_;
	wire _01446_;
	wire _01447_;
	wire _01448_;
	wire _01449_;
	wire _01450_;
	wire _01451_;
	wire _01452_;
	wire _01453_;
	wire _01454_;
	wire _01455_;
	wire _01456_;
	wire _01457_;
	wire _01458_;
	wire _01459_;
	wire _01460_;
	wire _01461_;
	wire _01462_;
	wire _01463_;
	wire _01464_;
	wire _01465_;
	wire _01466_;
	wire _01467_;
	wire _01468_;
	wire _01469_;
	wire _01470_;
	wire _01471_;
	wire _01472_;
	wire _01473_;
	wire _01474_;
	wire _01475_;
	wire _01476_;
	wire _01477_;
	wire _01478_;
	wire _01479_;
	wire _01480_;
	wire _01481_;
	wire _01482_;
	wire _01483_;
	wire _01484_;
	wire _01485_;
	wire _01486_;
	wire _01487_;
	wire _01488_;
	wire _01489_;
	wire _01490_;
	wire _01491_;
	wire _01492_;
	wire _01493_;
	wire _01494_;
	wire _01495_;
	wire _01496_;
	wire _01497_;
	wire _01498_;
	wire _01499_;
	wire _01500_;
	wire _01501_;
	wire _01502_;
	wire _01503_;
	wire _01504_;
	wire _01505_;
	wire _01506_;
	wire _01507_;
	wire _01508_;
	wire _01509_;
	wire _01510_;
	wire _01511_;
	wire _01512_;
	wire _01513_;
	wire _01514_;
	wire _01515_;
	wire _01516_;
	wire _01517_;
	wire _01518_;
	wire _01519_;
	wire _01520_;
	wire _01521_;
	wire _01522_;
	wire _01523_;
	wire _01524_;
	wire _01525_;
	wire _01526_;
	wire _01527_;
	wire _01528_;
	wire _01529_;
	wire _01530_;
	wire _01531_;
	wire _01532_;
	wire _01533_;
	wire _01534_;
	wire _01535_;
	wire _01536_;
	wire _01537_;
	wire _01538_;
	wire _01539_;
	wire _01540_;
	wire _01541_;
	wire _01542_;
	wire _01543_;
	wire _01544_;
	wire _01545_;
	wire _01546_;
	wire _01547_;
	wire _01548_;
	wire _01549_;
	wire _01550_;
	wire _01551_;
	wire _01552_;
	wire _01553_;
	wire _01554_;
	wire _01555_;
	wire _01556_;
	wire _01557_;
	wire _01558_;
	wire _01559_;
	wire _01560_;
	wire _01561_;
	wire _01562_;
	wire _01563_;
	wire _01564_;
	wire _01565_;
	wire _01566_;
	wire _01567_;
	wire _01568_;
	wire _01569_;
	wire _01570_;
	wire _01571_;
	wire _01572_;
	wire _01573_;
	wire _01574_;
	wire _01575_;
	wire _01576_;
	wire _01577_;
	wire _01578_;
	wire _01579_;
	wire _01580_;
	wire _01581_;
	wire _01582_;
	wire _01583_;
	wire _01584_;
	wire _01585_;
	wire _01586_;
	wire _01587_;
	wire _01588_;
	wire _01589_;
	wire _01590_;
	wire _01591_;
	wire _01592_;
	wire _01593_;
	wire _01594_;
	wire _01595_;
	wire _01596_;
	wire _01597_;
	wire _01598_;
	wire _01599_;
	wire _01600_;
	wire _01601_;
	wire _01602_;
	wire _01603_;
	wire _01604_;
	wire _01605_;
	wire _01606_;
	wire _01607_;
	wire _01608_;
	wire _01609_;
	wire _01610_;
	wire _01611_;
	wire _01612_;
	wire _01613_;
	wire _01614_;
	wire _01615_;
	wire _01616_;
	wire _01617_;
	wire _01618_;
	wire _01619_;
	wire _01620_;
	wire _01621_;
	wire _01622_;
	wire _01623_;
	wire _01624_;
	wire _01625_;
	wire _01626_;
	wire _01627_;
	wire _01628_;
	wire _01629_;
	wire _01630_;
	wire _01631_;
	wire _01632_;
	wire _01633_;
	wire _01634_;
	wire _01635_;
	wire _01636_;
	wire _01637_;
	wire _01638_;
	wire _01639_;
	wire _01640_;
	wire _01641_;
	wire _01642_;
	wire _01643_;
	wire _01644_;
	wire _01645_;
	wire _01646_;
	wire _01647_;
	wire _01648_;
	wire _01649_;
	wire _01650_;
	wire _01651_;
	wire _01652_;
	wire _01653_;
	wire _01654_;
	wire _01655_;
	wire _01656_;
	wire _01657_;
	wire _01658_;
	wire _01659_;
	wire _01660_;
	wire _01661_;
	wire _01662_;
	wire _01663_;
	wire _01664_;
	wire _01665_;
	wire _01666_;
	wire _01667_;
	wire _01668_;
	wire _01669_;
	wire _01670_;
	wire _01671_;
	wire _01672_;
	wire _01673_;
	wire _01674_;
	wire _01675_;
	wire _01676_;
	wire _01677_;
	wire _01678_;
	wire _01679_;
	wire _01680_;
	wire _01681_;
	wire _01682_;
	wire _01683_;
	wire _01684_;
	wire _01685_;
	wire _01686_;
	wire _01687_;
	wire _01688_;
	wire _01689_;
	wire _01690_;
	wire _01691_;
	wire _01692_;
	wire _01693_;
	wire _01694_;
	wire _01695_;
	wire _01696_;
	wire _01697_;
	wire _01698_;
	wire _01699_;
	wire _01700_;
	wire _01701_;
	wire _01702_;
	wire _01703_;
	wire _01704_;
	wire _01705_;
	wire _01706_;
	wire _01707_;
	wire _01708_;
	wire _01709_;
	wire _01710_;
	wire _01711_;
	wire _01712_;
	wire _01713_;
	wire _01714_;
	wire _01715_;
	wire _01716_;
	wire _01717_;
	wire _01718_;
	wire _01719_;
	wire _01720_;
	wire _01721_;
	wire _01722_;
	wire _01723_;
	wire _01724_;
	wire _01725_;
	wire _01726_;
	wire _01727_;
	wire _01728_;
	wire _01729_;
	wire _01730_;
	wire _01731_;
	wire _01732_;
	wire _01733_;
	wire _01734_;
	wire _01735_;
	wire _01736_;
	wire _01737_;
	wire _01738_;
	wire _01739_;
	wire _01740_;
	wire _01741_;
	wire _01742_;
	wire _01743_;
	wire _01744_;
	wire _01745_;
	wire _01746_;
	wire _01747_;
	wire _01748_;
	wire _01749_;
	wire _01750_;
	wire _01751_;
	wire _01752_;
	wire _01753_;
	wire _01754_;
	wire _01755_;
	wire _01756_;
	wire _01757_;
	wire _01758_;
	wire _01759_;
	wire _01760_;
	wire _01761_;
	wire _01762_;
	wire _01763_;
	wire _01764_;
	wire _01765_;
	wire _01766_;
	wire _01767_;
	wire _01768_;
	wire _01769_;
	wire _01770_;
	wire _01771_;
	wire _01772_;
	wire _01773_;
	wire _01774_;
	wire _01775_;
	wire _01776_;
	wire _01777_;
	wire _01778_;
	wire _01779_;
	wire _01780_;
	wire _01781_;
	wire _01782_;
	wire _01783_;
	wire _01784_;
	wire _01785_;
	wire _01786_;
	wire _01787_;
	wire _01788_;
	wire _01789_;
	wire _01790_;
	wire _01791_;
	wire _01792_;
	wire _01793_;
	wire _01794_;
	wire _01795_;
	wire _01796_;
	wire _01797_;
	wire _01798_;
	wire _01799_;
	wire _01800_;
	wire _01801_;
	wire _01802_;
	wire _01803_;
	wire _01804_;
	wire _01805_;
	wire _01806_;
	wire _01807_;
	wire _01808_;
	wire _01809_;
	wire _01810_;
	wire _01811_;
	wire _01812_;
	wire _01813_;
	wire _01814_;
	wire _01815_;
	wire _01816_;
	wire _01817_;
	wire _01818_;
	wire _01819_;
	wire _01820_;
	wire _01821_;
	wire _01822_;
	wire _01823_;
	wire _01824_;
	wire _01825_;
	wire _01826_;
	wire _01827_;
	wire _01828_;
	wire _01829_;
	wire _01830_;
	wire _01831_;
	wire _01832_;
	wire _01833_;
	wire _01834_;
	wire _01835_;
	wire _01836_;
	wire _01837_;
	wire _01838_;
	wire _01839_;
	wire _01840_;
	wire _01841_;
	wire _01842_;
	wire _01843_;
	wire _01844_;
	wire _01845_;
	wire _01846_;
	wire _01847_;
	wire _01848_;
	wire _01849_;
	wire _01850_;
	wire _01851_;
	wire _01852_;
	wire _01853_;
	wire _01854_;
	wire _01855_;
	wire _01856_;
	wire _01857_;
	wire _01858_;
	wire _01859_;
	wire _01860_;
	wire _01861_;
	wire _01862_;
	wire _01863_;
	wire _01864_;
	wire _01865_;
	wire _01866_;
	wire _01867_;
	wire _01868_;
	wire _01869_;
	wire _01870_;
	wire _01871_;
	wire _01872_;
	wire _01873_;
	wire _01874_;
	wire _01875_;
	wire _01876_;
	wire _01877_;
	wire _01878_;
	wire _01879_;
	wire _01880_;
	wire _01881_;
	wire _01882_;
	wire _01883_;
	wire _01884_;
	wire _01885_;
	wire _01886_;
	wire _01887_;
	wire _01888_;
	wire _01889_;
	wire _01890_;
	wire _01891_;
	wire _01892_;
	wire _01893_;
	wire _01894_;
	wire _01895_;
	wire _01896_;
	wire _01897_;
	wire _01898_;
	wire _01899_;
	wire _01900_;
	wire _01901_;
	wire _01902_;
	wire _01903_;
	wire _01904_;
	wire _01905_;
	wire _01906_;
	wire _01907_;
	wire _01908_;
	wire _01909_;
	wire _01910_;
	wire _01911_;
	wire _01912_;
	wire _01913_;
	wire _01914_;
	wire _01915_;
	wire _01916_;
	wire _01917_;
	wire _01918_;
	wire _01919_;
	wire _01920_;
	wire _01921_;
	wire _01922_;
	wire _01923_;
	wire _01924_;
	wire _01925_;
	wire _01926_;
	wire _01927_;
	wire _01928_;
	wire _01929_;
	wire _01930_;
	wire _01931_;
	wire _01932_;
	wire _01933_;
	wire _01934_;
	wire _01935_;
	wire _01936_;
	wire _01937_;
	wire _01938_;
	wire _01939_;
	wire _01940_;
	wire _01941_;
	wire _01942_;
	wire _01943_;
	wire _01944_;
	wire _01945_;
	wire _01946_;
	wire _01947_;
	wire _01948_;
	wire _01949_;
	wire _01950_;
	wire _01951_;
	wire _01952_;
	wire _01953_;
	wire _01954_;
	wire _01955_;
	wire _01956_;
	wire _01957_;
	wire _01958_;
	wire _01959_;
	wire _01960_;
	wire _01961_;
	wire _01962_;
	wire _01963_;
	wire _01964_;
	wire _01965_;
	wire _01966_;
	wire _01967_;
	wire _01968_;
	wire _01969_;
	wire _01970_;
	wire _01971_;
	wire _01972_;
	wire _01973_;
	wire _01974_;
	wire _01975_;
	wire _01976_;
	wire _01977_;
	wire _01978_;
	wire _01979_;
	wire _01980_;
	wire _01981_;
	wire _01982_;
	wire _01983_;
	wire _01984_;
	wire _01985_;
	wire _01986_;
	wire _01987_;
	wire _01988_;
	wire _01989_;
	wire _01990_;
	wire _01991_;
	wire _01992_;
	wire _01993_;
	wire _01994_;
	wire _01995_;
	wire _01996_;
	wire _01997_;
	wire _01998_;
	wire _01999_;
	wire _02000_;
	wire _02001_;
	wire _02002_;
	wire _02003_;
	wire _02004_;
	wire _02005_;
	wire _02006_;
	wire _02007_;
	wire _02008_;
	wire _02009_;
	wire _02010_;
	wire _02011_;
	wire _02012_;
	wire _02013_;
	wire _02014_;
	wire _02015_;
	wire _02016_;
	wire _02017_;
	wire _02018_;
	wire _02019_;
	wire _02020_;
	wire _02021_;
	wire _02022_;
	wire _02023_;
	wire _02024_;
	wire _02025_;
	wire _02026_;
	wire _02027_;
	wire _02028_;
	wire _02029_;
	wire _02030_;
	wire _02031_;
	wire _02032_;
	wire _02033_;
	wire _02034_;
	wire _02035_;
	wire _02036_;
	wire _02037_;
	wire _02038_;
	wire _02039_;
	wire _02040_;
	wire _02041_;
	wire _02042_;
	wire _02043_;
	wire _02044_;
	wire _02045_;
	wire _02046_;
	wire _02047_;
	wire _02048_;
	wire _02049_;
	wire _02050_;
	wire _02051_;
	wire _02052_;
	wire _02053_;
	wire _02054_;
	wire _02055_;
	wire _02056_;
	wire _02057_;
	wire _02058_;
	wire _02059_;
	wire _02060_;
	wire _02061_;
	wire _02062_;
	wire _02063_;
	wire _02064_;
	wire _02065_;
	wire _02066_;
	wire _02067_;
	wire _02068_;
	wire _02069_;
	wire _02070_;
	wire _02071_;
	wire _02072_;
	wire _02073_;
	wire _02074_;
	wire _02075_;
	wire _02076_;
	wire _02077_;
	wire _02078_;
	wire _02079_;
	wire _02080_;
	wire _02081_;
	wire _02082_;
	wire _02083_;
	wire _02084_;
	wire _02085_;
	wire _02086_;
	wire _02087_;
	wire _02088_;
	wire _02089_;
	wire _02090_;
	wire _02091_;
	wire _02092_;
	wire _02093_;
	wire _02094_;
	wire _02095_;
	wire _02096_;
	wire _02097_;
	wire _02098_;
	wire _02099_;
	wire _02100_;
	wire _02101_;
	wire _02102_;
	wire _02103_;
	wire _02104_;
	wire _02105_;
	wire _02106_;
	wire _02107_;
	wire _02108_;
	wire _02109_;
	wire _02110_;
	wire _02111_;
	wire _02112_;
	wire _02113_;
	wire _02114_;
	wire _02115_;
	wire _02116_;
	wire _02117_;
	wire _02118_;
	wire _02119_;
	wire _02120_;
	wire _02121_;
	wire _02122_;
	wire _02123_;
	wire _02124_;
	wire _02125_;
	wire _02126_;
	wire _02127_;
	wire _02128_;
	wire _02129_;
	wire _02130_;
	wire _02131_;
	wire _02132_;
	wire _02133_;
	wire _02134_;
	wire _02135_;
	wire _02136_;
	wire _02137_;
	wire _02138_;
	wire _02139_;
	wire _02140_;
	wire _02141_;
	wire _02142_;
	wire _02143_;
	wire _02144_;
	wire _02145_;
	wire _02146_;
	wire _02147_;
	wire _02148_;
	wire _02149_;
	wire _02150_;
	wire _02151_;
	wire _02152_;
	wire _02153_;
	wire _02154_;
	wire _02155_;
	wire _02156_;
	wire _02157_;
	wire _02158_;
	wire _02159_;
	wire _02160_;
	wire _02161_;
	wire _02162_;
	wire _02163_;
	wire _02164_;
	wire _02165_;
	wire _02166_;
	wire _02167_;
	wire _02168_;
	wire _02169_;
	wire _02170_;
	wire _02171_;
	wire _02172_;
	wire _02173_;
	wire _02174_;
	wire _02175_;
	wire _02176_;
	wire _02177_;
	wire _02178_;
	wire _02179_;
	wire _02180_;
	wire _02181_;
	wire _02182_;
	wire _02183_;
	wire _02184_;
	wire _02185_;
	wire _02186_;
	wire _02187_;
	wire _02188_;
	wire _02189_;
	wire _02190_;
	wire _02191_;
	wire _02192_;
	wire _02193_;
	wire _02194_;
	wire _02195_;
	wire _02196_;
	wire _02197_;
	wire _02198_;
	wire _02199_;
	wire _02200_;
	wire _02201_;
	wire _02202_;
	wire _02203_;
	wire _02204_;
	wire _02205_;
	wire _02206_;
	wire _02207_;
	wire _02208_;
	wire _02209_;
	wire _02210_;
	wire _02211_;
	wire _02212_;
	wire _02213_;
	wire _02214_;
	wire _02215_;
	wire _02216_;
	wire _02217_;
	wire _02218_;
	wire _02219_;
	wire _02220_;
	wire _02221_;
	wire _02222_;
	wire _02223_;
	wire _02224_;
	wire _02225_;
	wire _02226_;
	wire _02227_;
	wire _02228_;
	wire _02229_;
	wire _02230_;
	wire _02231_;
	wire _02232_;
	wire _02233_;
	wire _02234_;
	wire _02235_;
	wire _02236_;
	wire _02237_;
	wire _02238_;
	wire _02239_;
	wire _02240_;
	wire _02241_;
	wire _02242_;
	wire _02243_;
	wire _02244_;
	wire _02245_;
	wire _02246_;
	wire _02247_;
	wire _02248_;
	wire _02249_;
	wire _02250_;
	wire _02251_;
	wire _02252_;
	wire _02253_;
	wire _02254_;
	wire _02255_;
	wire _02256_;
	wire _02257_;
	wire _02258_;
	wire _02259_;
	wire _02260_;
	wire _02261_;
	wire _02262_;
	wire _02263_;
	wire _02264_;
	wire _02265_;
	wire _02266_;
	wire _02267_;
	wire _02268_;
	wire _02269_;
	wire _02270_;
	wire _02271_;
	wire _02272_;
	wire _02273_;
	wire _02274_;
	wire _02275_;
	wire _02276_;
	wire _02277_;
	wire _02278_;
	wire _02279_;
	wire _02280_;
	wire _02281_;
	wire _02282_;
	wire _02283_;
	wire _02284_;
	wire _02285_;
	wire _02286_;
	wire _02287_;
	wire _02288_;
	wire _02289_;
	wire _02290_;
	wire _02291_;
	wire _02292_;
	wire _02293_;
	wire _02294_;
	wire _02295_;
	wire _02296_;
	wire _02297_;
	wire _02298_;
	wire _02299_;
	wire _02300_;
	wire _02301_;
	wire _02302_;
	wire _02303_;
	wire _02304_;
	wire _02305_;
	wire _02306_;
	wire _02307_;
	wire _02308_;
	wire _02309_;
	wire _02310_;
	wire _02311_;
	wire _02312_;
	wire _02313_;
	wire _02314_;
	wire _02315_;
	wire _02316_;
	wire _02317_;
	wire _02318_;
	wire _02319_;
	wire _02320_;
	wire _02321_;
	wire _02322_;
	wire _02323_;
	wire _02324_;
	wire _02325_;
	wire _02326_;
	wire _02327_;
	wire _02328_;
	wire _02329_;
	wire _02330_;
	wire _02331_;
	wire _02332_;
	wire _02333_;
	wire _02334_;
	wire _02335_;
	wire _02336_;
	wire _02337_;
	wire _02338_;
	wire _02339_;
	wire _02340_;
	wire _02341_;
	wire _02342_;
	wire _02343_;
	wire _02344_;
	wire _02345_;
	wire _02346_;
	wire _02347_;
	wire _02348_;
	wire _02349_;
	wire _02350_;
	wire _02351_;
	wire _02352_;
	wire _02353_;
	wire _02354_;
	wire _02355_;
	wire _02356_;
	wire _02357_;
	wire _02358_;
	wire _02359_;
	wire _02360_;
	wire _02361_;
	wire _02362_;
	wire _02363_;
	wire _02364_;
	wire _02365_;
	wire _02366_;
	wire _02367_;
	wire _02368_;
	wire _02369_;
	wire _02370_;
	wire _02371_;
	wire _02372_;
	wire _02373_;
	wire _02374_;
	wire _02375_;
	wire _02376_;
	wire _02377_;
	wire _02378_;
	wire _02379_;
	wire _02380_;
	wire _02381_;
	wire _02382_;
	wire _02383_;
	wire _02384_;
	wire _02385_;
	wire _02386_;
	wire _02387_;
	wire _02388_;
	wire _02389_;
	wire _02390_;
	wire _02391_;
	wire _02392_;
	wire _02393_;
	wire _02394_;
	wire _02395_;
	wire _02396_;
	wire _02397_;
	wire _02398_;
	wire _02399_;
	wire _02400_;
	wire _02401_;
	wire _02402_;
	wire _02403_;
	wire _02404_;
	wire _02405_;
	wire _02406_;
	wire _02407_;
	wire _02408_;
	wire _02409_;
	wire _02410_;
	wire _02411_;
	wire _02412_;
	wire _02413_;
	wire _02414_;
	wire _02415_;
	wire _02416_;
	wire _02417_;
	wire _02418_;
	wire _02419_;
	wire _02420_;
	wire _02421_;
	wire _02422_;
	wire _02423_;
	wire _02424_;
	wire _02425_;
	wire _02426_;
	wire _02427_;
	wire _02428_;
	wire _02429_;
	wire _02430_;
	wire _02431_;
	wire _02432_;
	wire _02433_;
	wire _02434_;
	wire _02435_;
	wire _02436_;
	wire _02437_;
	wire _02438_;
	wire _02439_;
	wire _02440_;
	wire _02441_;
	wire _02442_;
	wire _02443_;
	wire _02444_;
	wire _02445_;
	wire _02446_;
	wire _02447_;
	wire _02448_;
	wire _02449_;
	wire _02450_;
	wire _02451_;
	wire _02452_;
	wire _02453_;
	wire _02454_;
	wire _02455_;
	wire _02456_;
	wire _02457_;
	wire _02458_;
	wire _02459_;
	wire _02460_;
	wire _02461_;
	wire _02462_;
	wire _02463_;
	wire _02464_;
	wire _02465_;
	wire _02466_;
	wire _02467_;
	wire _02468_;
	wire _02469_;
	wire _02470_;
	wire _02471_;
	wire _02472_;
	wire _02473_;
	wire _02474_;
	wire _02475_;
	wire _02476_;
	wire _02477_;
	wire _02478_;
	wire _02479_;
	wire _02480_;
	wire _02481_;
	wire _02482_;
	wire _02483_;
	wire _02484_;
	wire _02485_;
	wire _02486_;
	wire _02487_;
	wire _02488_;
	wire _02489_;
	wire _02490_;
	wire _02491_;
	wire _02492_;
	wire _02493_;
	wire _02494_;
	wire _02495_;
	wire _02496_;
	wire _02497_;
	wire _02498_;
	wire _02499_;
	wire _02500_;
	wire _02501_;
	wire _02502_;
	wire _02503_;
	wire _02504_;
	wire _02505_;
	wire _02506_;
	wire _02507_;
	wire _02508_;
	wire _02509_;
	wire _02510_;
	wire _02511_;
	wire _02512_;
	wire _02513_;
	wire _02514_;
	wire _02515_;
	wire _02516_;
	wire _02517_;
	wire _02518_;
	wire _02519_;
	wire _02520_;
	wire _02521_;
	wire _02522_;
	wire _02523_;
	wire _02524_;
	wire _02525_;
	wire _02526_;
	wire _02527_;
	wire _02528_;
	wire _02529_;
	wire _02530_;
	wire _02531_;
	wire _02532_;
	wire _02533_;
	wire _02534_;
	wire _02535_;
	wire _02536_;
	wire _02537_;
	wire _02538_;
	wire _02539_;
	wire _02540_;
	wire _02541_;
	wire _02542_;
	wire _02543_;
	wire _02544_;
	wire _02545_;
	wire _02546_;
	wire _02547_;
	wire _02548_;
	wire _02549_;
	wire _02550_;
	wire _02551_;
	wire _02552_;
	wire _02553_;
	wire _02554_;
	wire _02555_;
	wire _02556_;
	wire _02557_;
	wire _02558_;
	wire _02559_;
	wire _02560_;
	wire _02561_;
	wire _02562_;
	wire _02563_;
	wire _02564_;
	wire _02565_;
	wire _02566_;
	wire _02567_;
	wire _02568_;
	wire _02569_;
	wire _02570_;
	wire _02571_;
	wire _02572_;
	wire _02573_;
	wire _02574_;
	wire _02575_;
	wire _02576_;
	wire _02577_;
	wire _02578_;
	wire _02579_;
	wire _02580_;
	wire _02581_;
	wire _02582_;
	wire _02583_;
	wire _02584_;
	wire _02585_;
	wire _02586_;
	wire _02587_;
	wire _02588_;
	wire _02589_;
	wire _02590_;
	wire _02591_;
	wire _02592_;
	wire _02593_;
	wire _02594_;
	wire _02595_;
	wire _02596_;
	wire _02597_;
	wire _02598_;
	wire _02599_;
	wire _02600_;
	wire _02601_;
	wire _02602_;
	wire _02603_;
	wire _02604_;
	wire _02605_;
	wire _02606_;
	wire _02607_;
	wire _02608_;
	wire _02609_;
	wire _02610_;
	wire _02611_;
	wire _02612_;
	wire _02613_;
	wire _02614_;
	wire _02615_;
	wire _02616_;
	wire _02617_;
	wire _02618_;
	wire _02619_;
	wire _02620_;
	wire _02621_;
	wire _02622_;
	wire _02623_;
	wire _02624_;
	wire _02625_;
	wire _02626_;
	wire _02627_;
	wire _02628_;
	wire _02629_;
	wire _02630_;
	wire _02631_;
	wire _02632_;
	wire _02633_;
	wire _02634_;
	wire _02635_;
	wire _02636_;
	wire _02637_;
	wire _02638_;
	wire _02639_;
	wire _02640_;
	wire _02641_;
	wire _02642_;
	wire _02643_;
	wire _02644_;
	wire _02645_;
	wire _02646_;
	wire _02647_;
	wire _02648_;
	wire _02649_;
	wire _02650_;
	wire _02651_;
	wire _02652_;
	wire _02653_;
	wire _02654_;
	wire _02655_;
	wire _02656_;
	wire _02657_;
	wire _02658_;
	wire _02659_;
	wire _02660_;
	wire _02661_;
	wire _02662_;
	wire _02663_;
	wire _02664_;
	wire _02665_;
	wire _02666_;
	wire _02667_;
	wire _02668_;
	wire _02669_;
	wire _02670_;
	wire _02671_;
	wire _02672_;
	wire _02673_;
	wire _02674_;
	wire _02675_;
	wire _02676_;
	wire _02677_;
	wire _02678_;
	wire _02679_;
	wire _02680_;
	wire _02681_;
	wire _02682_;
	wire _02683_;
	wire _02684_;
	wire _02685_;
	wire _02686_;
	wire _02687_;
	wire _02688_;
	wire _02689_;
	wire _02690_;
	wire _02691_;
	wire _02692_;
	wire _02693_;
	wire _02694_;
	wire _02695_;
	wire _02696_;
	wire _02697_;
	wire _02698_;
	wire _02699_;
	wire _02700_;
	wire _02701_;
	wire _02702_;
	wire _02703_;
	wire _02704_;
	wire _02705_;
	wire _02706_;
	wire _02707_;
	wire _02708_;
	wire _02709_;
	wire _02710_;
	wire _02711_;
	wire _02712_;
	wire _02713_;
	wire _02714_;
	wire _02715_;
	wire _02716_;
	wire _02717_;
	wire _02718_;
	wire _02719_;
	wire _02720_;
	wire _02721_;
	wire _02722_;
	wire _02723_;
	wire _02724_;
	wire _02725_;
	wire _02726_;
	wire _02727_;
	wire _02728_;
	wire _02729_;
	wire _02730_;
	wire _02731_;
	wire _02732_;
	wire _02733_;
	wire _02734_;
	wire _02735_;
	wire _02736_;
	wire _02737_;
	wire _02738_;
	wire _02739_;
	wire _02740_;
	wire _02741_;
	wire _02742_;
	wire _02743_;
	wire _02744_;
	wire _02745_;
	wire _02746_;
	wire _02747_;
	wire _02748_;
	wire _02749_;
	wire _02750_;
	wire _02751_;
	wire _02752_;
	wire _02753_;
	wire _02754_;
	wire _02755_;
	wire _02756_;
	wire _02757_;
	wire _02758_;
	wire _02759_;
	wire _02760_;
	wire _02761_;
	wire _02762_;
	wire _02763_;
	wire _02764_;
	wire _02765_;
	wire _02766_;
	wire _02767_;
	wire _02768_;
	wire _02769_;
	wire _02770_;
	wire _02771_;
	wire _02772_;
	wire _02773_;
	wire _02774_;
	wire _02775_;
	wire _02776_;
	wire _02777_;
	wire _02778_;
	wire _02779_;
	wire _02780_;
	wire _02781_;
	wire _02782_;
	wire _02783_;
	wire _02784_;
	wire _02785_;
	wire _02786_;
	wire _02787_;
	wire _02788_;
	wire _02789_;
	wire _02790_;
	wire _02791_;
	wire _02792_;
	wire _02793_;
	wire _02794_;
	wire _02795_;
	wire _02796_;
	wire _02797_;
	wire _02798_;
	wire _02799_;
	wire _02800_;
	wire _02801_;
	wire _02802_;
	wire _02803_;
	wire _02804_;
	wire _02805_;
	wire _02806_;
	wire _02807_;
	wire _02808_;
	wire _02809_;
	wire _02810_;
	wire _02811_;
	wire _02812_;
	wire _02813_;
	wire _02814_;
	wire _02815_;
	wire _02816_;
	wire _02817_;
	wire _02818_;
	wire _02819_;
	wire _02820_;
	wire _02821_;
	wire _02822_;
	wire _02823_;
	wire _02824_;
	wire _02825_;
	wire _02826_;
	wire _02827_;
	wire _02828_;
	wire _02829_;
	wire _02830_;
	wire _02831_;
	wire _02832_;
	wire _02833_;
	wire _02834_;
	wire _02835_;
	wire _02836_;
	wire _02837_;
	wire _02838_;
	wire _02839_;
	wire _02840_;
	wire _02841_;
	wire _02842_;
	wire _02843_;
	wire _02844_;
	wire _02845_;
	wire _02846_;
	wire _02847_;
	wire _02848_;
	wire _02849_;
	wire _02850_;
	wire _02851_;
	wire _02852_;
	wire _02853_;
	wire _02854_;
	wire _02855_;
	wire _02856_;
	wire _02857_;
	wire _02858_;
	wire _02859_;
	wire _02860_;
	wire _02861_;
	wire _02862_;
	wire _02863_;
	wire _02864_;
	wire _02865_;
	wire _02866_;
	wire _02867_;
	wire _02868_;
	wire _02869_;
	wire _02870_;
	wire _02871_;
	wire _02872_;
	wire _02873_;
	wire _02874_;
	wire _02875_;
	wire _02876_;
	wire _02877_;
	wire _02878_;
	wire _02879_;
	wire _02880_;
	wire _02881_;
	wire _02882_;
	wire _02883_;
	wire _02884_;
	wire _02885_;
	wire _02886_;
	wire _02887_;
	wire _02888_;
	wire _02889_;
	wire _02890_;
	wire _02891_;
	wire _02892_;
	wire _02893_;
	wire _02894_;
	wire _02895_;
	wire _02896_;
	wire _02897_;
	wire _02898_;
	wire _02899_;
	wire _02900_;
	wire _02901_;
	wire _02902_;
	wire _02903_;
	wire _02904_;
	wire _02905_;
	wire _02906_;
	wire _02907_;
	wire _02908_;
	wire _02909_;
	wire _02910_;
	wire _02911_;
	wire _02912_;
	wire _02913_;
	wire _02914_;
	wire _02915_;
	wire _02916_;
	wire _02917_;
	wire _02918_;
	wire _02919_;
	wire _02920_;
	wire _02921_;
	wire _02922_;
	wire _02923_;
	wire _02924_;
	wire _02925_;
	wire _02926_;
	wire _02927_;
	wire _02928_;
	wire _02929_;
	wire _02930_;
	wire _02931_;
	wire _02932_;
	wire _02933_;
	wire _02934_;
	wire _02935_;
	wire _02936_;
	wire _02937_;
	wire _02938_;
	wire _02939_;
	wire _02940_;
	wire _02941_;
	wire _02942_;
	wire _02943_;
	wire _02944_;
	wire _02945_;
	wire _02946_;
	wire _02947_;
	wire _02948_;
	wire _02949_;
	wire _02950_;
	wire _02951_;
	wire _02952_;
	wire _02953_;
	wire _02954_;
	wire _02955_;
	wire _02956_;
	wire _02957_;
	wire _02958_;
	wire _02959_;
	wire _02960_;
	wire _02961_;
	wire _02962_;
	wire _02963_;
	wire _02964_;
	wire _02965_;
	wire _02966_;
	wire _02967_;
	wire _02968_;
	wire _02969_;
	wire _02970_;
	wire _02971_;
	wire _02972_;
	wire _02973_;
	wire _02974_;
	wire _02975_;
	wire _02976_;
	wire _02977_;
	wire _02978_;
	wire _02979_;
	wire _02980_;
	wire _02981_;
	wire _02982_;
	wire _02983_;
	wire _02984_;
	wire _02985_;
	wire _02986_;
	wire _02987_;
	wire _02988_;
	wire _02989_;
	wire _02990_;
	wire _02991_;
	wire _02992_;
	wire _02993_;
	wire _02994_;
	wire _02995_;
	wire _02996_;
	wire _02997_;
	wire _02998_;
	wire _02999_;
	wire _03000_;
	wire _03001_;
	wire _03002_;
	wire _03003_;
	wire _03004_;
	wire _03005_;
	wire _03006_;
	wire _03007_;
	wire _03008_;
	wire _03009_;
	wire _03010_;
	wire _03011_;
	wire _03012_;
	wire _03013_;
	wire _03014_;
	wire _03015_;
	wire _03016_;
	wire _03017_;
	wire _03018_;
	wire _03019_;
	wire _03020_;
	wire _03021_;
	wire _03022_;
	wire _03023_;
	wire _03024_;
	wire _03025_;
	wire _03026_;
	wire _03027_;
	wire _03028_;
	wire _03029_;
	wire _03030_;
	wire _03031_;
	wire _03032_;
	wire _03033_;
	wire _03034_;
	wire _03035_;
	wire _03036_;
	wire _03037_;
	wire _03038_;
	wire _03039_;
	wire _03040_;
	wire _03041_;
	wire _03042_;
	wire _03043_;
	wire _03044_;
	wire _03045_;
	wire _03046_;
	wire _03047_;
	wire _03048_;
	wire _03049_;
	wire _03050_;
	wire _03051_;
	wire _03052_;
	wire _03053_;
	wire _03054_;
	wire _03055_;
	wire _03056_;
	wire _03057_;
	wire _03058_;
	wire _03059_;
	wire _03060_;
	wire _03061_;
	wire _03062_;
	wire _03063_;
	wire _03064_;
	wire _03065_;
	wire _03066_;
	wire _03067_;
	wire _03068_;
	wire _03069_;
	wire _03070_;
	wire _03071_;
	wire _03072_;
	wire _03073_;
	wire _03074_;
	wire _03075_;
	wire _03076_;
	wire _03077_;
	wire _03078_;
	wire _03079_;
	wire _03080_;
	wire _03081_;
	wire _03082_;
	wire _03083_;
	wire _03084_;
	wire _03085_;
	wire _03086_;
	wire _03087_;
	wire _03088_;
	wire _03089_;
	wire _03090_;
	wire _03091_;
	wire _03092_;
	wire _03093_;
	wire _03094_;
	wire _03095_;
	wire _03096_;
	wire _03097_;
	wire _03098_;
	wire _03099_;
	wire _03100_;
	wire _03101_;
	wire _03102_;
	wire _03103_;
	wire _03104_;
	wire _03105_;
	wire _03106_;
	wire _03107_;
	wire _03108_;
	wire _03109_;
	wire _03110_;
	wire _03111_;
	wire _03112_;
	wire _03113_;
	wire _03114_;
	wire _03115_;
	wire _03116_;
	wire _03117_;
	wire _03118_;
	wire _03119_;
	wire _03120_;
	wire _03121_;
	wire _03122_;
	wire _03123_;
	wire _03124_;
	wire _03125_;
	wire _03126_;
	wire _03127_;
	wire _03128_;
	wire _03129_;
	wire _03130_;
	wire _03131_;
	wire _03132_;
	wire _03133_;
	wire _03134_;
	wire _03135_;
	wire _03136_;
	wire _03137_;
	wire _03138_;
	wire _03139_;
	wire _03140_;
	wire _03141_;
	wire _03142_;
	wire _03143_;
	wire _03144_;
	wire _03145_;
	wire _03146_;
	wire _03147_;
	wire _03148_;
	wire _03149_;
	wire _03150_;
	wire _03151_;
	wire _03152_;
	wire _03153_;
	wire _03154_;
	wire _03155_;
	wire _03156_;
	wire _03157_;
	wire _03158_;
	wire _03159_;
	wire _03160_;
	wire _03161_;
	wire _03162_;
	wire _03163_;
	wire _03164_;
	wire _03165_;
	wire _03166_;
	wire _03167_;
	wire _03168_;
	wire _03169_;
	wire _03170_;
	wire _03171_;
	wire _03172_;
	wire _03173_;
	wire _03174_;
	wire _03175_;
	wire _03176_;
	wire _03177_;
	wire _03178_;
	wire _03179_;
	wire _03180_;
	wire _03181_;
	wire _03182_;
	wire _03183_;
	wire _03184_;
	wire _03185_;
	wire _03186_;
	wire _03187_;
	wire _03188_;
	wire _03189_;
	wire _03190_;
	wire _03191_;
	wire _03192_;
	wire _03193_;
	wire _03194_;
	wire _03195_;
	wire _03196_;
	wire _03197_;
	wire _03198_;
	wire _03199_;
	wire _03200_;
	wire _03201_;
	wire _03202_;
	wire _03203_;
	wire _03204_;
	wire _03205_;
	wire _03206_;
	wire _03207_;
	wire _03208_;
	wire _03209_;
	wire _03210_;
	wire _03211_;
	wire _03212_;
	wire _03213_;
	wire _03214_;
	wire _03215_;
	wire _03216_;
	wire _03217_;
	wire _03218_;
	wire _03219_;
	wire _03220_;
	wire _03221_;
	wire _03222_;
	wire _03223_;
	wire _03224_;
	wire _03225_;
	wire _03226_;
	wire _03227_;
	wire _03228_;
	wire _03229_;
	wire _03230_;
	wire _03231_;
	wire _03232_;
	wire _03233_;
	wire _03234_;
	wire _03235_;
	wire _03236_;
	wire _03237_;
	wire _03238_;
	wire _03239_;
	wire _03240_;
	wire _03241_;
	wire _03242_;
	wire _03243_;
	wire _03244_;
	wire _03245_;
	wire _03246_;
	wire _03247_;
	wire _03248_;
	wire _03249_;
	wire _03250_;
	wire _03251_;
	wire _03252_;
	wire _03253_;
	wire _03254_;
	wire _03255_;
	wire _03256_;
	wire _03257_;
	wire _03258_;
	wire _03259_;
	wire _03260_;
	wire _03261_;
	wire _03262_;
	wire _03263_;
	wire _03264_;
	wire _03265_;
	wire _03266_;
	wire _03267_;
	wire _03268_;
	wire _03269_;
	wire _03270_;
	wire _03271_;
	wire _03272_;
	wire _03273_;
	wire _03274_;
	wire _03275_;
	wire _03276_;
	wire _03277_;
	wire _03278_;
	wire _03279_;
	wire _03280_;
	wire _03281_;
	wire _03282_;
	wire _03283_;
	wire _03284_;
	wire _03285_;
	wire _03286_;
	wire _03287_;
	wire _03288_;
	wire _03289_;
	wire _03290_;
	wire _03291_;
	wire _03292_;
	wire _03293_;
	wire _03294_;
	wire _03295_;
	wire _03296_;
	wire _03297_;
	wire _03298_;
	wire _03299_;
	wire _03300_;
	wire _03301_;
	wire _03302_;
	wire _03303_;
	wire _03304_;
	wire _03305_;
	wire _03306_;
	wire _03307_;
	wire _03308_;
	wire _03309_;
	wire _03310_;
	wire _03311_;
	wire _03312_;
	wire _03313_;
	wire _03314_;
	wire _03315_;
	wire _03316_;
	wire _03317_;
	wire _03318_;
	wire _03319_;
	wire _03320_;
	wire _03321_;
	wire _03322_;
	wire _03323_;
	wire _03324_;
	wire _03325_;
	wire _03326_;
	wire _03327_;
	wire _03328_;
	wire _03329_;
	wire _03330_;
	wire _03331_;
	wire _03332_;
	wire _03333_;
	wire _03334_;
	wire _03335_;
	wire _03336_;
	wire _03337_;
	wire _03338_;
	wire _03339_;
	wire _03340_;
	wire _03341_;
	wire _03342_;
	wire _03343_;
	wire _03344_;
	wire _03345_;
	wire _03346_;
	wire _03347_;
	wire _03348_;
	wire _03349_;
	wire _03350_;
	wire _03351_;
	wire _03352_;
	wire _03353_;
	wire _03354_;
	wire _03355_;
	wire _03356_;
	wire _03357_;
	wire _03358_;
	wire _03359_;
	wire _03360_;
	wire _03361_;
	wire _03362_;
	wire _03363_;
	wire _03364_;
	wire _03365_;
	wire _03366_;
	wire _03367_;
	wire _03368_;
	wire _03369_;
	wire _03370_;
	wire _03371_;
	wire _03372_;
	wire _03373_;
	wire _03374_;
	wire _03375_;
	wire _03376_;
	wire _03377_;
	wire _03378_;
	wire _03379_;
	wire _03380_;
	wire _03381_;
	wire _03382_;
	wire _03383_;
	wire _03384_;
	wire _03385_;
	wire _03386_;
	wire _03387_;
	wire _03388_;
	wire _03389_;
	wire _03390_;
	wire _03391_;
	wire _03392_;
	wire _03393_;
	wire _03394_;
	wire _03395_;
	wire _03396_;
	wire _03397_;
	wire _03398_;
	wire _03399_;
	wire _03400_;
	wire _03401_;
	wire _03402_;
	wire _03403_;
	wire _03404_;
	wire _03405_;
	wire _03406_;
	wire _03407_;
	wire _03408_;
	wire _03409_;
	wire _03410_;
	wire _03411_;
	wire _03412_;
	wire _03413_;
	wire _03414_;
	wire _03415_;
	wire _03416_;
	wire _03417_;
	wire _03418_;
	wire _03419_;
	wire _03420_;
	wire _03421_;
	wire _03422_;
	wire _03423_;
	wire _03424_;
	wire _03425_;
	wire _03426_;
	wire _03427_;
	wire _03428_;
	wire _03429_;
	wire _03430_;
	wire _03431_;
	wire _03432_;
	wire _03433_;
	wire _03434_;
	wire _03435_;
	wire _03436_;
	wire _03437_;
	wire _03438_;
	wire _03439_;
	wire _03440_;
	wire _03441_;
	wire _03442_;
	wire _03443_;
	wire _03444_;
	wire _03445_;
	wire _03446_;
	wire _03447_;
	wire _03448_;
	wire _03449_;
	wire _03450_;
	wire _03451_;
	wire _03452_;
	wire _03453_;
	wire _03454_;
	wire _03455_;
	wire _03456_;
	wire _03457_;
	wire _03458_;
	wire _03459_;
	wire _03460_;
	wire _03461_;
	wire _03462_;
	wire _03463_;
	wire _03464_;
	wire _03465_;
	wire _03466_;
	wire _03467_;
	wire _03468_;
	wire _03469_;
	wire _03470_;
	wire _03471_;
	wire _03472_;
	wire _03473_;
	wire _03474_;
	wire _03475_;
	wire _03476_;
	wire _03477_;
	wire _03478_;
	wire _03479_;
	wire _03480_;
	wire _03481_;
	wire _03482_;
	wire _03483_;
	wire _03484_;
	wire _03485_;
	wire _03486_;
	wire _03487_;
	wire _03488_;
	wire _03489_;
	wire _03490_;
	wire _03491_;
	wire _03492_;
	wire _03493_;
	wire _03494_;
	wire _03495_;
	wire _03496_;
	wire _03497_;
	wire _03498_;
	wire _03499_;
	wire _03500_;
	wire _03501_;
	wire _03502_;
	wire _03503_;
	wire _03504_;
	wire _03505_;
	wire _03506_;
	wire _03507_;
	wire _03508_;
	wire _03509_;
	wire _03510_;
	wire _03511_;
	wire _03512_;
	wire _03513_;
	wire _03514_;
	wire _03515_;
	wire _03516_;
	wire _03517_;
	wire _03518_;
	wire _03519_;
	wire _03520_;
	wire _03521_;
	wire _03522_;
	wire _03523_;
	wire _03524_;
	wire _03525_;
	wire _03526_;
	wire _03527_;
	wire _03528_;
	wire _03529_;
	wire _03530_;
	wire _03531_;
	wire _03532_;
	wire _03533_;
	wire _03534_;
	wire _03535_;
	wire _03536_;
	wire _03537_;
	wire _03538_;
	wire _03539_;
	wire _03540_;
	wire _03541_;
	wire _03542_;
	wire _03543_;
	wire _03544_;
	wire _03545_;
	wire _03546_;
	wire _03547_;
	wire _03548_;
	wire _03549_;
	wire _03550_;
	wire _03551_;
	wire _03552_;
	wire _03553_;
	wire _03554_;
	wire _03555_;
	wire _03556_;
	wire _03557_;
	wire _03558_;
	wire _03559_;
	wire _03560_;
	wire _03561_;
	wire _03562_;
	wire _03563_;
	wire _03564_;
	wire _03565_;
	wire _03566_;
	wire _03567_;
	wire _03568_;
	wire _03569_;
	wire _03570_;
	wire _03571_;
	wire _03572_;
	wire _03573_;
	wire _03574_;
	wire _03575_;
	wire _03576_;
	wire _03577_;
	wire _03578_;
	wire _03579_;
	wire _03580_;
	wire _03581_;
	wire _03582_;
	wire _03583_;
	wire _03584_;
	wire _03585_;
	wire _03586_;
	wire _03587_;
	wire _03588_;
	wire _03589_;
	wire _03590_;
	wire _03591_;
	wire _03592_;
	wire _03593_;
	wire _03594_;
	wire _03595_;
	wire _03596_;
	wire _03597_;
	wire _03598_;
	wire _03599_;
	wire _03600_;
	wire _03601_;
	wire _03602_;
	wire _03603_;
	wire _03604_;
	wire _03605_;
	wire _03606_;
	wire _03607_;
	wire _03608_;
	wire _03609_;
	wire _03610_;
	wire _03611_;
	wire _03612_;
	wire _03613_;
	wire _03614_;
	wire _03615_;
	wire _03616_;
	wire _03617_;
	wire _03618_;
	wire _03619_;
	wire _03620_;
	wire _03621_;
	wire _03622_;
	wire _03623_;
	wire _03624_;
	wire _03625_;
	wire _03626_;
	wire _03627_;
	wire _03628_;
	wire _03629_;
	wire _03630_;
	wire _03631_;
	wire _03632_;
	wire _03633_;
	wire _03634_;
	wire _03635_;
	wire _03636_;
	wire _03637_;
	wire _03638_;
	wire _03639_;
	wire _03640_;
	wire _03641_;
	wire _03642_;
	wire _03643_;
	wire _03644_;
	wire _03645_;
	wire _03646_;
	wire _03647_;
	wire _03648_;
	wire _03649_;
	wire _03650_;
	wire _03651_;
	wire _03652_;
	wire _03653_;
	wire _03654_;
	wire _03655_;
	wire _03656_;
	wire _03657_;
	wire _03658_;
	wire _03659_;
	wire _03660_;
	wire _03661_;
	wire _03662_;
	wire _03663_;
	wire _03664_;
	wire _03665_;
	wire _03666_;
	wire _03667_;
	wire _03668_;
	wire _03669_;
	wire _03670_;
	wire _03671_;
	wire _03672_;
	wire _03673_;
	wire _03674_;
	wire _03675_;
	wire _03676_;
	wire _03677_;
	wire _03678_;
	wire _03679_;
	wire _03680_;
	wire _03681_;
	wire _03682_;
	wire _03683_;
	wire _03684_;
	wire _03685_;
	wire _03686_;
	wire _03687_;
	wire _03688_;
	wire _03689_;
	wire _03690_;
	wire _03691_;
	wire _03692_;
	wire _03693_;
	wire _03694_;
	wire _03695_;
	wire _03696_;
	wire _03697_;
	wire _03698_;
	wire _03699_;
	wire _03700_;
	wire _03701_;
	wire _03702_;
	wire _03703_;
	wire _03704_;
	wire _03705_;
	wire _03706_;
	wire _03707_;
	wire _03708_;
	wire _03709_;
	wire _03710_;
	wire _03711_;
	wire _03712_;
	wire _03713_;
	wire _03714_;
	wire _03715_;
	wire _03716_;
	wire _03717_;
	wire _03718_;
	wire _03719_;
	wire _03720_;
	wire _03721_;
	wire _03722_;
	wire _03723_;
	wire _03724_;
	wire _03725_;
	wire _03726_;
	wire _03727_;
	wire _03728_;
	wire _03729_;
	wire _03730_;
	wire _03731_;
	wire _03732_;
	wire _03733_;
	wire _03734_;
	wire _03735_;
	wire _03736_;
	wire _03737_;
	wire _03738_;
	wire _03739_;
	wire _03740_;
	wire _03741_;
	wire _03742_;
	wire _03743_;
	wire _03744_;
	wire _03745_;
	wire _03746_;
	wire _03747_;
	wire _03748_;
	wire _03749_;
	wire _03750_;
	wire _03751_;
	wire _03752_;
	wire _03753_;
	wire _03754_;
	wire _03755_;
	wire _03756_;
	wire _03757_;
	wire _03758_;
	wire _03759_;
	wire _03760_;
	wire _03761_;
	wire _03762_;
	wire _03763_;
	wire _03764_;
	wire _03765_;
	wire _03766_;
	wire _03767_;
	wire _03768_;
	wire _03769_;
	wire _03770_;
	wire _03771_;
	wire _03772_;
	wire _03773_;
	wire _03774_;
	wire _03775_;
	wire _03776_;
	wire _03777_;
	wire _03778_;
	wire _03779_;
	wire _03780_;
	wire _03781_;
	wire _03782_;
	wire _03783_;
	wire _03784_;
	wire _03785_;
	wire _03786_;
	wire _03787_;
	wire _03788_;
	wire _03789_;
	wire _03790_;
	wire _03791_;
	wire _03792_;
	wire _03793_;
	wire _03794_;
	wire _03795_;
	wire _03796_;
	wire _03797_;
	wire _03798_;
	wire _03799_;
	wire _03800_;
	wire _03801_;
	wire _03802_;
	wire _03803_;
	wire _03804_;
	wire _03805_;
	wire _03806_;
	wire _03807_;
	wire _03808_;
	wire _03809_;
	wire _03810_;
	wire _03811_;
	wire _03812_;
	wire _03813_;
	wire _03814_;
	wire _03815_;
	wire _03816_;
	wire _03817_;
	wire _03818_;
	wire _03819_;
	wire _03820_;
	wire _03821_;
	wire _03822_;
	wire _03823_;
	wire _03824_;
	wire _03825_;
	wire _03826_;
	wire _03827_;
	wire _03828_;
	wire _03829_;
	wire _03830_;
	wire _03831_;
	wire _03832_;
	wire _03833_;
	wire _03834_;
	wire _03835_;
	wire _03836_;
	wire _03837_;
	wire _03838_;
	wire _03839_;
	wire _03840_;
	wire _03841_;
	wire _03842_;
	wire _03843_;
	wire _03844_;
	wire _03845_;
	wire _03846_;
	wire _03847_;
	wire _03848_;
	wire _03849_;
	wire _03850_;
	wire _03851_;
	wire _03852_;
	wire _03853_;
	wire _03854_;
	wire _03855_;
	wire _03856_;
	wire _03857_;
	wire _03858_;
	wire _03859_;
	wire _03860_;
	wire _03861_;
	wire _03862_;
	wire _03863_;
	wire _03864_;
	wire _03865_;
	wire _03866_;
	wire _03867_;
	wire _03868_;
	wire _03869_;
	wire _03870_;
	wire _03871_;
	wire _03872_;
	wire _03873_;
	wire _03874_;
	wire _03875_;
	wire _03876_;
	wire _03877_;
	wire _03878_;
	wire _03879_;
	wire _03880_;
	wire _03881_;
	wire _03882_;
	wire _03883_;
	wire _03884_;
	wire _03885_;
	wire _03886_;
	wire _03887_;
	wire _03888_;
	wire _03889_;
	wire _03890_;
	wire _03891_;
	wire _03892_;
	wire _03893_;
	wire _03894_;
	wire _03895_;
	wire _03896_;
	wire _03897_;
	wire _03898_;
	wire _03899_;
	wire _03900_;
	wire _03901_;
	wire _03902_;
	wire _03903_;
	wire _03904_;
	wire _03905_;
	wire _03906_;
	wire _03907_;
	wire _03908_;
	wire _03909_;
	wire _03910_;
	wire _03911_;
	wire _03912_;
	wire _03913_;
	wire _03914_;
	wire _03915_;
	wire _03916_;
	wire _03917_;
	wire _03918_;
	wire _03919_;
	wire _03920_;
	wire _03921_;
	wire _03922_;
	wire _03923_;
	wire _03924_;
	wire _03925_;
	wire _03926_;
	wire _03927_;
	wire _03928_;
	wire _03929_;
	wire _03930_;
	wire _03931_;
	wire _03932_;
	wire _03933_;
	wire _03934_;
	wire _03935_;
	wire _03936_;
	wire _03937_;
	wire _03938_;
	wire _03939_;
	wire _03940_;
	wire _03941_;
	wire _03942_;
	wire _03943_;
	wire _03944_;
	wire _03945_;
	wire _03946_;
	wire _03947_;
	wire _03948_;
	wire _03949_;
	wire _03950_;
	wire _03951_;
	wire _03952_;
	wire _03953_;
	wire _03954_;
	wire _03955_;
	wire _03956_;
	wire _03957_;
	wire _03958_;
	wire _03959_;
	wire _03960_;
	wire _03961_;
	wire _03962_;
	wire _03963_;
	wire _03964_;
	wire _03965_;
	wire _03966_;
	wire _03967_;
	wire _03968_;
	wire _03969_;
	wire _03970_;
	wire _03971_;
	wire _03972_;
	wire _03973_;
	wire _03974_;
	wire _03975_;
	wire _03976_;
	wire _03977_;
	wire _03978_;
	wire _03979_;
	wire _03980_;
	wire _03981_;
	wire _03982_;
	wire _03983_;
	wire _03984_;
	wire _03985_;
	wire _03986_;
	wire _03987_;
	wire _03988_;
	wire _03989_;
	wire _03990_;
	wire _03991_;
	wire _03992_;
	wire _03993_;
	wire _03994_;
	wire _03995_;
	wire _03996_;
	wire _03997_;
	wire _03998_;
	wire _03999_;
	wire _04000_;
	wire _04001_;
	wire _04002_;
	wire _04003_;
	wire _04004_;
	wire _04005_;
	wire _04006_;
	wire _04007_;
	wire _04008_;
	wire _04009_;
	wire _04010_;
	wire _04011_;
	wire _04012_;
	wire _04013_;
	wire _04014_;
	wire _04015_;
	wire _04016_;
	wire _04017_;
	wire _04018_;
	wire _04019_;
	wire _04020_;
	wire _04021_;
	wire _04022_;
	wire _04023_;
	wire _04024_;
	wire _04025_;
	wire _04026_;
	wire _04027_;
	wire _04028_;
	wire _04029_;
	wire _04030_;
	wire _04031_;
	wire _04032_;
	wire _04033_;
	wire _04034_;
	wire _04035_;
	wire _04036_;
	wire _04037_;
	wire _04038_;
	wire _04039_;
	wire _04040_;
	wire _04041_;
	wire _04042_;
	wire _04043_;
	wire _04044_;
	wire _04045_;
	wire _04046_;
	wire _04047_;
	wire _04048_;
	wire _04049_;
	wire _04050_;
	wire _04051_;
	wire _04052_;
	wire _04053_;
	wire _04054_;
	wire _04055_;
	wire _04056_;
	wire _04057_;
	wire _04058_;
	wire _04059_;
	wire _04060_;
	wire _04061_;
	wire _04062_;
	wire _04063_;
	wire _04064_;
	wire _04065_;
	wire _04066_;
	wire _04067_;
	wire _04068_;
	wire _04069_;
	wire _04070_;
	wire _04071_;
	wire _04072_;
	wire _04073_;
	wire _04074_;
	wire _04075_;
	wire _04076_;
	wire _04077_;
	wire _04078_;
	wire _04079_;
	wire _04080_;
	wire _04081_;
	wire _04082_;
	wire _04083_;
	wire _04084_;
	wire _04085_;
	wire _04086_;
	wire _04087_;
	wire _04088_;
	wire _04089_;
	wire _04090_;
	wire _04091_;
	wire _04092_;
	wire _04093_;
	wire _04094_;
	wire _04095_;
	wire _04096_;
	wire _04097_;
	wire _04098_;
	wire _04099_;
	wire _04100_;
	wire _04101_;
	wire _04102_;
	wire _04103_;
	wire _04104_;
	wire _04105_;
	wire _04106_;
	wire _04107_;
	wire _04108_;
	wire _04109_;
	wire _04110_;
	wire _04111_;
	wire _04112_;
	wire _04113_;
	wire _04114_;
	wire _04115_;
	wire _04116_;
	wire _04117_;
	wire _04118_;
	wire _04119_;
	wire _04120_;
	wire _04121_;
	wire _04122_;
	wire _04123_;
	wire _04124_;
	wire _04125_;
	wire _04126_;
	wire _04127_;
	wire _04128_;
	wire _04129_;
	wire _04130_;
	wire _04131_;
	wire _04132_;
	wire _04133_;
	wire _04134_;
	wire _04135_;
	wire _04136_;
	wire _04137_;
	wire _04138_;
	wire _04139_;
	wire _04140_;
	wire _04141_;
	wire _04142_;
	wire _04143_;
	wire _04144_;
	wire _04145_;
	wire _04146_;
	wire _04147_;
	wire _04148_;
	wire _04149_;
	wire _04150_;
	wire _04151_;
	wire _04152_;
	wire _04153_;
	wire _04154_;
	wire _04155_;
	wire _04156_;
	wire _04157_;
	wire _04158_;
	wire _04159_;
	wire _04160_;
	wire _04161_;
	wire _04162_;
	wire _04163_;
	wire _04164_;
	wire _04165_;
	wire _04166_;
	wire _04167_;
	wire _04168_;
	wire _04169_;
	wire _04170_;
	wire _04171_;
	wire _04172_;
	wire _04173_;
	wire _04174_;
	wire _04175_;
	wire _04176_;
	wire _04177_;
	wire _04178_;
	wire _04179_;
	wire _04180_;
	wire _04181_;
	wire _04182_;
	wire _04183_;
	wire _04184_;
	wire _04185_;
	wire _04186_;
	wire _04187_;
	wire _04188_;
	wire _04189_;
	wire _04190_;
	wire _04191_;
	wire _04192_;
	wire _04193_;
	wire _04194_;
	wire _04195_;
	wire _04196_;
	wire _04197_;
	wire _04198_;
	wire _04199_;
	wire _04200_;
	wire _04201_;
	wire _04202_;
	wire _04203_;
	wire _04204_;
	wire _04205_;
	wire _04206_;
	wire _04207_;
	wire _04208_;
	wire _04209_;
	wire _04210_;
	wire _04211_;
	wire _04212_;
	wire _04213_;
	wire _04214_;
	wire _04215_;
	wire _04216_;
	wire _04217_;
	wire _04218_;
	wire _04219_;
	wire _04220_;
	wire _04221_;
	wire _04222_;
	wire _04223_;
	wire _04224_;
	wire _04225_;
	wire _04226_;
	wire _04227_;
	wire _04228_;
	wire _04229_;
	wire _04230_;
	wire _04231_;
	wire _04232_;
	wire _04233_;
	wire _04234_;
	wire _04235_;
	wire _04236_;
	wire _04237_;
	wire _04238_;
	wire _04239_;
	wire _04240_;
	wire _04241_;
	wire _04242_;
	wire _04243_;
	wire _04244_;
	wire _04245_;
	wire _04246_;
	wire _04247_;
	wire _04248_;
	wire _04249_;
	wire _04250_;
	wire _04251_;
	wire _04252_;
	wire _04253_;
	wire _04254_;
	wire _04255_;
	wire _04256_;
	wire _04257_;
	wire _04258_;
	wire _04259_;
	wire _04260_;
	wire _04261_;
	wire _04262_;
	wire _04263_;
	wire _04264_;
	wire _04265_;
	wire _04266_;
	wire _04267_;
	wire _04268_;
	wire _04269_;
	wire _04270_;
	wire _04271_;
	wire _04272_;
	wire _04273_;
	wire _04274_;
	wire _04275_;
	wire _04276_;
	wire _04277_;
	wire _04278_;
	wire _04279_;
	wire _04280_;
	wire _04281_;
	wire _04282_;
	wire _04283_;
	wire _04284_;
	wire _04285_;
	wire _04286_;
	wire _04287_;
	wire _04288_;
	wire _04289_;
	wire _04290_;
	wire _04291_;
	wire _04292_;
	wire _04293_;
	wire _04294_;
	wire _04295_;
	wire _04296_;
	wire _04297_;
	wire _04298_;
	wire _04299_;
	wire _04300_;
	wire _04301_;
	wire _04302_;
	wire _04303_;
	wire _04304_;
	wire _04305_;
	wire _04306_;
	wire _04307_;
	wire _04308_;
	wire _04309_;
	wire _04310_;
	wire _04311_;
	wire _04312_;
	wire _04313_;
	wire _04314_;
	wire _04315_;
	wire _04316_;
	wire _04317_;
	wire _04318_;
	wire _04319_;
	wire _04320_;
	wire _04321_;
	wire _04322_;
	wire _04323_;
	wire _04324_;
	wire _04325_;
	wire _04326_;
	wire _04327_;
	wire _04328_;
	wire _04329_;
	wire _04330_;
	wire _04331_;
	wire _04332_;
	wire _04333_;
	wire _04334_;
	wire _04335_;
	wire _04336_;
	wire _04337_;
	wire _04338_;
	wire _04339_;
	wire _04340_;
	wire _04341_;
	wire _04342_;
	wire _04343_;
	wire _04344_;
	wire _04345_;
	wire _04346_;
	wire _04347_;
	wire _04348_;
	wire _04349_;
	wire _04350_;
	wire _04351_;
	wire _04352_;
	wire _04353_;
	wire _04354_;
	wire _04355_;
	wire _04356_;
	wire _04357_;
	wire _04358_;
	wire _04359_;
	wire _04360_;
	wire _04361_;
	wire _04362_;
	wire _04363_;
	wire _04364_;
	wire _04365_;
	wire _04366_;
	wire _04367_;
	wire _04368_;
	wire _04369_;
	wire _04370_;
	wire _04371_;
	wire _04372_;
	wire _04373_;
	wire _04374_;
	wire _04375_;
	wire _04376_;
	wire _04377_;
	wire _04378_;
	wire _04379_;
	wire _04380_;
	wire _04381_;
	wire _04382_;
	wire _04383_;
	wire _04384_;
	wire _04385_;
	wire _04386_;
	wire _04387_;
	wire _04388_;
	wire _04389_;
	wire _04390_;
	wire _04391_;
	wire _04392_;
	wire _04393_;
	wire _04394_;
	wire _04395_;
	wire _04396_;
	wire _04397_;
	wire _04398_;
	wire _04399_;
	wire _04400_;
	wire _04401_;
	wire _04402_;
	wire _04403_;
	wire _04404_;
	wire _04405_;
	wire _04406_;
	wire _04407_;
	wire _04408_;
	wire _04409_;
	wire _04410_;
	wire _04411_;
	wire _04412_;
	wire _04413_;
	wire _04414_;
	wire _04415_;
	wire _04416_;
	wire _04417_;
	wire _04418_;
	wire _04419_;
	wire _04420_;
	wire _04421_;
	wire _04422_;
	wire _04423_;
	wire _04424_;
	wire _04425_;
	wire _04426_;
	wire _04427_;
	wire _04428_;
	wire _04429_;
	wire _04430_;
	wire _04431_;
	wire _04432_;
	wire _04433_;
	wire _04434_;
	wire _04435_;
	wire _04436_;
	wire _04437_;
	wire _04438_;
	wire _04439_;
	wire _04440_;
	wire _04441_;
	wire _04442_;
	wire _04443_;
	wire _04444_;
	wire _04445_;
	wire _04446_;
	wire _04447_;
	wire _04448_;
	wire _04449_;
	wire _04450_;
	wire _04451_;
	wire _04452_;
	wire _04453_;
	wire _04454_;
	wire _04455_;
	wire _04456_;
	wire _04457_;
	wire _04458_;
	wire _04459_;
	wire _04460_;
	wire _04461_;
	wire _04462_;
	wire _04463_;
	wire _04464_;
	wire _04465_;
	wire _04466_;
	wire _04467_;
	wire _04468_;
	wire _04469_;
	wire _04470_;
	wire _04471_;
	wire _04472_;
	wire _04473_;
	wire _04474_;
	wire _04475_;
	wire _04476_;
	wire _04477_;
	wire _04478_;
	wire _04479_;
	wire _04480_;
	wire _04481_;
	wire _04482_;
	wire _04483_;
	wire _04484_;
	wire _04485_;
	wire _04486_;
	wire _04487_;
	wire _04488_;
	wire _04489_;
	wire _04490_;
	wire _04491_;
	wire _04492_;
	wire _04493_;
	wire _04494_;
	wire _04495_;
	wire _04496_;
	wire _04497_;
	wire _04498_;
	wire _04499_;
	wire _04500_;
	wire _04501_;
	wire _04502_;
	wire _04503_;
	wire _04504_;
	wire _04505_;
	wire _04506_;
	wire _04507_;
	wire _04508_;
	wire _04509_;
	wire _04510_;
	wire _04511_;
	wire _04512_;
	wire _04513_;
	wire _04514_;
	wire _04515_;
	wire _04516_;
	wire _04517_;
	wire _04518_;
	wire _04519_;
	wire _04520_;
	wire _04521_;
	wire _04522_;
	wire _04523_;
	wire _04524_;
	wire _04525_;
	wire _04526_;
	wire _04527_;
	wire _04528_;
	wire _04529_;
	wire _04530_;
	wire _04531_;
	wire _04532_;
	wire _04533_;
	wire _04534_;
	wire _04535_;
	wire _04536_;
	wire _04537_;
	wire _04538_;
	wire _04539_;
	wire _04540_;
	wire _04541_;
	wire _04542_;
	wire _04543_;
	wire _04544_;
	wire _04545_;
	wire _04546_;
	wire _04547_;
	wire _04548_;
	wire _04549_;
	wire _04550_;
	wire _04551_;
	wire _04552_;
	wire _04553_;
	wire _04554_;
	wire _04555_;
	wire _04556_;
	wire _04557_;
	wire _04558_;
	wire _04559_;
	wire _04560_;
	wire _04561_;
	wire _04562_;
	wire _04563_;
	wire _04564_;
	wire _04565_;
	wire _04566_;
	wire _04567_;
	wire _04568_;
	wire _04569_;
	wire _04570_;
	wire _04571_;
	wire _04572_;
	wire _04573_;
	wire _04574_;
	wire _04575_;
	wire _04576_;
	wire _04577_;
	wire _04578_;
	wire _04579_;
	wire _04580_;
	wire _04581_;
	wire _04582_;
	wire _04583_;
	wire _04584_;
	wire _04585_;
	wire _04586_;
	wire _04587_;
	wire _04588_;
	wire _04589_;
	wire _04590_;
	wire _04591_;
	wire _04592_;
	wire _04593_;
	wire _04594_;
	wire _04595_;
	wire _04596_;
	wire _04597_;
	wire _04598_;
	wire _04599_;
	wire _04600_;
	wire _04601_;
	wire _04602_;
	wire _04603_;
	wire _04604_;
	wire _04605_;
	wire _04606_;
	wire _04607_;
	wire _04608_;
	wire _04609_;
	wire _04610_;
	wire _04611_;
	wire _04612_;
	wire _04613_;
	wire _04614_;
	wire _04615_;
	wire _04616_;
	wire _04617_;
	wire _04618_;
	wire _04619_;
	wire _04620_;
	wire _04621_;
	wire _04622_;
	wire _04623_;
	wire _04624_;
	wire _04625_;
	wire _04626_;
	wire _04627_;
	wire _04628_;
	wire _04629_;
	wire _04630_;
	wire _04631_;
	wire _04632_;
	wire _04633_;
	wire _04634_;
	wire _04635_;
	wire _04636_;
	wire _04637_;
	wire _04638_;
	wire _04639_;
	wire _04640_;
	wire _04641_;
	wire _04642_;
	wire _04643_;
	wire _04644_;
	wire _04645_;
	wire _04646_;
	wire _04647_;
	wire _04648_;
	wire _04649_;
	wire _04650_;
	wire _04651_;
	wire _04652_;
	wire _04653_;
	wire _04654_;
	wire _04655_;
	wire _04656_;
	wire _04657_;
	wire _04658_;
	wire _04659_;
	wire _04660_;
	wire _04661_;
	wire _04662_;
	wire _04663_;
	wire _04664_;
	wire _04665_;
	wire _04666_;
	wire _04667_;
	wire _04668_;
	wire _04669_;
	wire _04670_;
	wire _04671_;
	wire _04672_;
	wire _04673_;
	wire _04674_;
	wire _04675_;
	wire _04676_;
	wire _04677_;
	wire _04678_;
	wire _04679_;
	wire _04680_;
	wire _04681_;
	wire _04682_;
	wire _04683_;
	wire _04684_;
	wire _04685_;
	wire _04686_;
	wire _04687_;
	wire _04688_;
	wire _04689_;
	wire _04690_;
	wire _04691_;
	wire _04692_;
	wire _04693_;
	wire _04694_;
	wire _04695_;
	wire _04696_;
	wire _04697_;
	wire _04698_;
	wire _04699_;
	wire _04700_;
	wire _04701_;
	wire _04702_;
	wire _04703_;
	wire _04704_;
	wire _04705_;
	wire _04706_;
	wire _04707_;
	wire _04708_;
	wire _04709_;
	wire _04710_;
	wire _04711_;
	wire _04712_;
	wire _04713_;
	wire _04714_;
	wire _04715_;
	wire _04716_;
	wire _04717_;
	wire _04718_;
	wire _04719_;
	wire _04720_;
	wire _04721_;
	wire _04722_;
	wire _04723_;
	wire _04724_;
	wire _04725_;
	wire _04726_;
	wire _04727_;
	wire _04728_;
	wire _04729_;
	wire _04730_;
	wire _04731_;
	wire _04732_;
	wire _04733_;
	wire _04734_;
	wire _04735_;
	wire _04736_;
	wire _04737_;
	wire _04738_;
	wire _04739_;
	wire _04740_;
	wire _04741_;
	wire _04742_;
	wire _04743_;
	wire _04744_;
	wire _04745_;
	wire _04746_;
	wire _04747_;
	wire _04748_;
	wire _04749_;
	wire _04750_;
	wire _04751_;
	wire _04752_;
	wire _04753_;
	wire _04754_;
	wire _04755_;
	wire _04756_;
	wire _04757_;
	wire _04758_;
	wire _04759_;
	wire _04760_;
	wire _04761_;
	wire _04762_;
	wire _04763_;
	wire _04764_;
	wire _04765_;
	wire _04766_;
	wire _04767_;
	wire _04768_;
	wire _04769_;
	wire _04770_;
	wire _04771_;
	wire _04772_;
	wire _04773_;
	wire _04774_;
	wire _04775_;
	wire _04776_;
	wire _04777_;
	wire _04778_;
	wire _04779_;
	wire _04780_;
	wire _04781_;
	wire _04782_;
	wire _04783_;
	wire _04784_;
	wire _04785_;
	wire _04786_;
	wire _04787_;
	wire _04788_;
	wire _04789_;
	wire _04790_;
	wire _04791_;
	wire _04792_;
	wire _04793_;
	wire _04794_;
	wire _04795_;
	wire _04796_;
	wire _04797_;
	wire _04798_;
	wire _04799_;
	wire _04800_;
	wire _04801_;
	wire _04802_;
	wire _04803_;
	wire _04804_;
	wire _04805_;
	wire _04806_;
	wire _04807_;
	wire _04808_;
	wire _04809_;
	wire _04810_;
	wire _04811_;
	wire _04812_;
	wire _04813_;
	wire _04814_;
	wire _04815_;
	wire _04816_;
	wire _04817_;
	wire _04818_;
	wire _04819_;
	wire _04820_;
	wire _04821_;
	wire _04822_;
	wire _04823_;
	wire _04824_;
	wire _04825_;
	wire _04826_;
	wire _04827_;
	wire _04828_;
	wire _04829_;
	wire _04830_;
	wire _04831_;
	wire _04832_;
	wire _04833_;
	wire _04834_;
	wire _04835_;
	wire _04836_;
	wire _04837_;
	wire _04838_;
	wire _04839_;
	wire _04840_;
	wire _04841_;
	wire _04842_;
	wire _04843_;
	wire _04844_;
	wire _04845_;
	wire _04846_;
	wire _04847_;
	wire _04848_;
	wire _04849_;
	wire _04850_;
	wire _04851_;
	wire _04852_;
	wire _04853_;
	wire _04854_;
	wire _04855_;
	wire _04856_;
	wire _04857_;
	wire _04858_;
	wire _04859_;
	wire _04860_;
	wire _04861_;
	wire _04862_;
	wire _04863_;
	wire _04864_;
	wire _04865_;
	wire _04866_;
	wire _04867_;
	wire _04868_;
	wire _04869_;
	wire _04870_;
	wire _04871_;
	wire _04872_;
	wire _04873_;
	wire _04874_;
	wire _04875_;
	wire _04876_;
	wire _04877_;
	wire _04878_;
	wire _04879_;
	wire _04880_;
	wire _04881_;
	wire _04882_;
	wire _04883_;
	wire _04884_;
	wire _04885_;
	wire _04886_;
	wire _04887_;
	wire _04888_;
	wire _04889_;
	wire _04890_;
	wire _04891_;
	wire _04892_;
	wire _04893_;
	wire _04894_;
	wire _04895_;
	wire _04896_;
	wire _04897_;
	wire _04898_;
	wire _04899_;
	wire _04900_;
	wire _04901_;
	wire _04902_;
	wire _04903_;
	wire _04904_;
	wire _04905_;
	wire _04906_;
	wire _04907_;
	wire _04908_;
	wire _04909_;
	wire _04910_;
	wire _04911_;
	wire _04912_;
	wire _04913_;
	wire _04914_;
	wire _04915_;
	wire _04916_;
	wire _04917_;
	wire _04918_;
	wire _04919_;
	wire _04920_;
	wire _04921_;
	wire _04922_;
	wire _04923_;
	wire _04924_;
	wire _04925_;
	wire _04926_;
	wire _04927_;
	wire _04928_;
	wire _04929_;
	wire _04930_;
	wire _04931_;
	wire _04932_;
	wire _04933_;
	wire _04934_;
	wire _04935_;
	wire _04936_;
	wire _04937_;
	wire _04938_;
	wire _04939_;
	wire _04940_;
	wire _04941_;
	wire _04942_;
	wire _04943_;
	wire _04944_;
	wire _04945_;
	wire _04946_;
	wire _04947_;
	wire _04948_;
	wire _04949_;
	wire _04950_;
	wire _04951_;
	wire _04952_;
	wire _04953_;
	wire _04954_;
	wire _04955_;
	wire _04956_;
	wire _04957_;
	wire _04958_;
	wire _04959_;
	wire _04960_;
	wire _04961_;
	wire _04962_;
	wire _04963_;
	wire _04964_;
	wire _04965_;
	wire _04966_;
	wire _04967_;
	wire _04968_;
	wire _04969_;
	wire _04970_;
	wire _04971_;
	wire _04972_;
	wire _04973_;
	wire _04974_;
	wire _04975_;
	wire _04976_;
	wire _04977_;
	wire _04978_;
	wire _04979_;
	wire _04980_;
	wire _04981_;
	wire _04982_;
	wire _04983_;
	wire _04984_;
	wire _04985_;
	wire _04986_;
	wire _04987_;
	wire _04988_;
	wire _04989_;
	wire _04990_;
	wire _04991_;
	wire _04992_;
	wire _04993_;
	wire _04994_;
	wire _04995_;
	wire _04996_;
	wire _04997_;
	wire _04998_;
	wire _04999_;
	wire _05000_;
	wire _05001_;
	wire _05002_;
	wire _05003_;
	wire _05004_;
	wire _05005_;
	wire _05006_;
	wire _05007_;
	wire _05008_;
	wire _05009_;
	wire _05010_;
	wire _05011_;
	wire _05012_;
	wire _05013_;
	wire _05014_;
	wire _05015_;
	wire _05016_;
	wire _05017_;
	wire _05018_;
	wire _05019_;
	wire _05020_;
	wire _05021_;
	wire _05022_;
	wire _05023_;
	wire _05024_;
	wire _05025_;
	wire _05026_;
	wire _05027_;
	wire _05028_;
	wire _05029_;
	wire _05030_;
	wire _05031_;
	wire _05032_;
	wire _05033_;
	wire _05034_;
	wire _05035_;
	wire _05036_;
	wire _05037_;
	wire _05038_;
	wire _05039_;
	wire _05040_;
	wire _05041_;
	wire _05042_;
	wire _05043_;
	wire _05044_;
	wire _05045_;
	wire _05046_;
	wire _05047_;
	wire _05048_;
	wire _05049_;
	wire _05050_;
	wire _05051_;
	wire _05052_;
	wire _05053_;
	wire _05054_;
	wire _05055_;
	wire _05056_;
	wire _05057_;
	wire _05058_;
	wire _05059_;
	wire _05060_;
	wire _05061_;
	wire _05062_;
	wire _05063_;
	wire _05064_;
	wire _05065_;
	wire _05066_;
	wire _05067_;
	wire _05068_;
	wire _05069_;
	wire _05070_;
	wire _05071_;
	wire _05072_;
	wire _05073_;
	wire _05074_;
	wire _05075_;
	wire _05076_;
	wire _05077_;
	wire _05078_;
	wire _05079_;
	wire _05080_;
	wire _05081_;
	wire _05082_;
	wire _05083_;
	wire _05084_;
	wire _05085_;
	wire _05086_;
	wire _05087_;
	wire _05088_;
	wire _05089_;
	wire _05090_;
	wire _05091_;
	wire _05092_;
	wire _05093_;
	wire _05094_;
	wire _05095_;
	wire _05096_;
	wire _05097_;
	wire _05098_;
	wire _05099_;
	wire _05100_;
	wire _05101_;
	wire _05102_;
	wire _05103_;
	wire _05104_;
	wire _05105_;
	wire _05106_;
	wire _05107_;
	wire _05108_;
	wire _05109_;
	wire _05110_;
	wire _05111_;
	wire _05112_;
	wire _05113_;
	wire _05114_;
	wire _05115_;
	wire _05116_;
	wire _05117_;
	wire _05118_;
	wire _05119_;
	wire _05120_;
	wire _05121_;
	wire _05122_;
	wire _05123_;
	wire _05124_;
	wire _05125_;
	wire _05126_;
	wire _05127_;
	wire _05128_;
	wire _05129_;
	wire _05130_;
	wire _05131_;
	wire _05132_;
	wire _05133_;
	wire _05134_;
	wire _05135_;
	wire _05136_;
	wire _05137_;
	wire _05138_;
	wire _05139_;
	wire _05140_;
	wire _05141_;
	wire _05142_;
	wire _05143_;
	wire _05144_;
	wire _05145_;
	wire _05146_;
	wire _05147_;
	wire _05148_;
	wire _05149_;
	wire _05150_;
	wire _05151_;
	wire _05152_;
	wire _05153_;
	wire _05154_;
	wire _05155_;
	wire _05156_;
	wire _05157_;
	wire _05158_;
	wire _05159_;
	wire _05160_;
	wire _05161_;
	wire _05162_;
	wire _05163_;
	wire _05164_;
	wire _05165_;
	wire _05166_;
	wire _05167_;
	wire _05168_;
	wire _05169_;
	wire _05170_;
	wire _05171_;
	wire _05172_;
	wire _05173_;
	wire _05174_;
	wire _05175_;
	wire _05176_;
	wire _05177_;
	wire _05178_;
	wire _05179_;
	wire _05180_;
	wire _05181_;
	wire _05182_;
	wire _05183_;
	wire _05184_;
	wire _05185_;
	wire _05186_;
	wire _05187_;
	wire _05188_;
	wire _05189_;
	wire _05190_;
	wire _05191_;
	wire _05192_;
	wire _05193_;
	wire _05194_;
	wire _05195_;
	wire _05196_;
	wire _05197_;
	wire _05198_;
	wire _05199_;
	wire _05200_;
	wire _05201_;
	wire _05202_;
	wire _05203_;
	wire _05204_;
	wire _05205_;
	wire _05206_;
	wire _05207_;
	wire _05208_;
	wire _05209_;
	wire _05210_;
	wire _05211_;
	wire _05212_;
	wire _05213_;
	wire _05214_;
	wire _05215_;
	wire _05216_;
	wire _05217_;
	wire _05218_;
	wire _05219_;
	wire _05220_;
	wire _05221_;
	wire _05222_;
	wire _05223_;
	wire _05224_;
	wire _05225_;
	wire _05226_;
	wire _05227_;
	wire _05228_;
	wire _05229_;
	wire _05230_;
	wire _05231_;
	wire _05232_;
	wire _05233_;
	wire _05234_;
	wire _05235_;
	wire _05236_;
	wire _05237_;
	wire _05238_;
	wire _05239_;
	wire _05240_;
	wire _05241_;
	wire _05242_;
	wire _05243_;
	wire _05244_;
	wire _05245_;
	wire _05246_;
	wire _05247_;
	wire _05248_;
	wire _05249_;
	wire _05250_;
	wire _05251_;
	wire _05252_;
	wire _05253_;
	wire _05254_;
	wire _05255_;
	wire _05256_;
	wire _05257_;
	wire _05258_;
	wire _05259_;
	wire _05260_;
	wire _05261_;
	wire _05262_;
	wire _05263_;
	wire _05264_;
	wire _05265_;
	wire _05266_;
	wire _05267_;
	wire _05268_;
	wire _05269_;
	wire _05270_;
	wire _05271_;
	wire _05272_;
	wire _05273_;
	wire _05274_;
	wire _05275_;
	wire _05276_;
	wire _05277_;
	wire _05278_;
	wire _05279_;
	wire _05280_;
	wire _05281_;
	wire _05282_;
	wire _05283_;
	wire _05284_;
	wire _05285_;
	wire _05286_;
	wire _05287_;
	wire _05288_;
	wire _05289_;
	wire _05290_;
	wire _05291_;
	wire _05292_;
	wire _05293_;
	wire _05294_;
	wire _05295_;
	wire _05296_;
	wire _05297_;
	wire _05298_;
	wire _05299_;
	wire _05300_;
	wire _05301_;
	wire _05302_;
	wire _05303_;
	wire _05304_;
	wire _05305_;
	wire _05306_;
	wire _05307_;
	wire _05308_;
	wire _05309_;
	wire _05310_;
	wire _05311_;
	wire _05312_;
	wire _05313_;
	wire _05314_;
	wire _05315_;
	wire _05316_;
	wire _05317_;
	wire _05318_;
	wire _05319_;
	wire _05320_;
	wire _05321_;
	wire _05322_;
	wire _05323_;
	wire _05324_;
	wire _05325_;
	wire _05326_;
	wire _05327_;
	wire _05328_;
	wire _05329_;
	wire _05330_;
	wire _05331_;
	wire _05332_;
	wire _05333_;
	wire _05334_;
	wire _05335_;
	wire _05336_;
	wire _05337_;
	wire _05338_;
	wire _05339_;
	wire _05340_;
	wire _05341_;
	wire _05342_;
	wire _05343_;
	wire _05344_;
	wire _05345_;
	wire _05346_;
	wire _05347_;
	wire _05348_;
	wire _05349_;
	wire _05350_;
	wire _05351_;
	wire _05352_;
	wire _05353_;
	wire _05354_;
	wire _05355_;
	wire _05356_;
	wire _05357_;
	wire _05358_;
	wire _05359_;
	wire _05360_;
	wire _05361_;
	wire _05362_;
	wire _05363_;
	wire _05364_;
	wire _05365_;
	wire _05366_;
	wire _05367_;
	wire _05368_;
	wire _05369_;
	wire _05370_;
	wire _05371_;
	wire _05372_;
	wire _05373_;
	wire _05374_;
	wire _05375_;
	wire _05376_;
	wire _05377_;
	wire _05378_;
	wire _05379_;
	wire _05380_;
	wire _05381_;
	wire _05382_;
	wire _05383_;
	wire _05384_;
	wire _05385_;
	wire _05386_;
	wire _05387_;
	wire _05388_;
	wire _05389_;
	wire _05390_;
	wire _05391_;
	wire _05392_;
	wire _05393_;
	wire _05394_;
	wire _05395_;
	wire _05396_;
	wire _05397_;
	wire _05398_;
	wire _05399_;
	wire _05400_;
	wire _05401_;
	wire _05402_;
	wire _05403_;
	wire _05404_;
	wire _05405_;
	wire _05406_;
	wire _05407_;
	wire _05408_;
	wire _05409_;
	wire _05410_;
	wire _05411_;
	wire _05412_;
	wire _05413_;
	wire _05414_;
	wire _05415_;
	wire _05416_;
	wire _05417_;
	wire _05418_;
	wire _05419_;
	wire _05420_;
	wire _05421_;
	wire _05422_;
	wire _05423_;
	wire _05424_;
	wire _05425_;
	wire _05426_;
	wire _05427_;
	wire _05428_;
	wire _05429_;
	wire _05430_;
	wire _05431_;
	wire _05432_;
	wire _05433_;
	wire _05434_;
	wire _05435_;
	wire _05436_;
	wire _05437_;
	wire _05438_;
	wire _05439_;
	wire _05440_;
	wire _05441_;
	wire _05442_;
	wire _05443_;
	wire _05444_;
	wire _05445_;
	wire _05446_;
	wire _05447_;
	wire _05448_;
	wire _05449_;
	wire _05450_;
	wire _05451_;
	wire _05452_;
	wire _05453_;
	wire _05454_;
	wire _05455_;
	wire _05456_;
	wire _05457_;
	wire _05458_;
	wire _05459_;
	wire _05460_;
	wire _05461_;
	wire _05462_;
	wire _05463_;
	wire _05464_;
	wire _05465_;
	wire _05466_;
	wire _05467_;
	wire _05468_;
	wire _05469_;
	wire _05470_;
	wire _05471_;
	wire _05472_;
	wire _05473_;
	wire _05474_;
	wire _05475_;
	wire _05476_;
	wire _05477_;
	wire _05478_;
	wire _05479_;
	wire _05480_;
	wire _05481_;
	wire _05482_;
	wire _05483_;
	wire _05484_;
	wire _05485_;
	wire _05486_;
	wire _05487_;
	wire _05488_;
	wire _05489_;
	wire _05490_;
	wire _05491_;
	wire _05492_;
	wire _05493_;
	wire _05494_;
	wire _05495_;
	wire _05496_;
	wire _05497_;
	wire _05498_;
	wire _05499_;
	wire _05500_;
	wire _05501_;
	wire _05502_;
	wire _05503_;
	wire _05504_;
	wire _05505_;
	wire _05506_;
	wire _05507_;
	wire _05508_;
	wire _05509_;
	wire _05510_;
	wire _05511_;
	wire _05512_;
	wire _05513_;
	wire _05514_;
	wire _05515_;
	wire _05516_;
	wire _05517_;
	wire _05518_;
	wire _05519_;
	wire _05520_;
	wire _05521_;
	wire _05522_;
	wire _05523_;
	wire _05524_;
	wire _05525_;
	wire _05526_;
	wire _05527_;
	wire _05528_;
	wire _05529_;
	wire _05530_;
	wire _05531_;
	wire _05532_;
	wire _05533_;
	wire _05534_;
	wire _05535_;
	wire _05536_;
	wire _05537_;
	wire _05538_;
	wire _05539_;
	wire _05540_;
	wire _05541_;
	wire _05542_;
	wire _05543_;
	wire _05544_;
	wire _05545_;
	wire _05546_;
	wire _05547_;
	wire _05548_;
	wire _05549_;
	wire _05550_;
	wire _05551_;
	wire _05552_;
	wire _05553_;
	wire _05554_;
	wire _05555_;
	wire _05556_;
	wire _05557_;
	wire _05558_;
	wire _05559_;
	wire _05560_;
	wire _05561_;
	wire _05562_;
	wire _05563_;
	wire _05564_;
	wire _05565_;
	wire _05566_;
	wire _05567_;
	wire _05568_;
	wire _05569_;
	wire _05570_;
	wire _05571_;
	wire _05572_;
	wire _05573_;
	wire _05574_;
	wire _05575_;
	wire _05576_;
	wire _05577_;
	wire _05578_;
	wire _05579_;
	wire _05580_;
	wire _05581_;
	wire _05582_;
	wire _05583_;
	wire _05584_;
	wire _05585_;
	wire _05586_;
	wire _05587_;
	wire _05588_;
	wire _05589_;
	wire _05590_;
	wire _05591_;
	wire _05592_;
	wire _05593_;
	wire _05594_;
	wire _05595_;
	wire _05596_;
	wire _05597_;
	wire _05598_;
	wire _05599_;
	wire _05600_;
	wire _05601_;
	wire _05602_;
	wire _05603_;
	wire _05604_;
	wire _05605_;
	wire _05606_;
	wire _05607_;
	wire _05608_;
	wire _05609_;
	wire _05610_;
	wire _05611_;
	wire _05612_;
	wire _05613_;
	wire _05614_;
	wire _05615_;
	wire _05616_;
	wire _05617_;
	wire _05618_;
	wire _05619_;
	wire _05620_;
	wire _05621_;
	wire _05622_;
	wire _05623_;
	wire _05624_;
	wire _05625_;
	wire _05626_;
	wire _05627_;
	wire _05628_;
	wire _05629_;
	wire _05630_;
	wire _05631_;
	wire _05632_;
	wire _05633_;
	wire _05634_;
	wire _05635_;
	wire _05636_;
	wire _05637_;
	wire _05638_;
	wire _05639_;
	wire _05640_;
	wire _05641_;
	wire _05642_;
	wire _05643_;
	wire _05644_;
	wire _05645_;
	wire _05646_;
	wire _05647_;
	wire _05648_;
	wire _05649_;
	wire _05650_;
	wire _05651_;
	wire _05652_;
	wire _05653_;
	wire _05654_;
	wire _05655_;
	wire _05656_;
	wire _05657_;
	wire _05658_;
	wire _05659_;
	wire _05660_;
	wire _05661_;
	wire _05662_;
	wire _05663_;
	wire _05664_;
	wire _05665_;
	wire _05666_;
	wire _05667_;
	wire _05668_;
	wire _05669_;
	wire _05670_;
	wire _05671_;
	wire _05672_;
	wire _05673_;
	wire _05674_;
	wire _05675_;
	wire _05676_;
	wire _05677_;
	wire _05678_;
	wire _05679_;
	wire _05680_;
	wire _05681_;
	wire _05682_;
	wire _05683_;
	wire _05684_;
	wire _05685_;
	wire _05686_;
	wire _05687_;
	wire _05688_;
	wire _05689_;
	wire _05690_;
	wire _05691_;
	wire _05692_;
	wire _05693_;
	wire _05694_;
	wire _05695_;
	wire _05696_;
	wire _05697_;
	wire _05698_;
	wire _05699_;
	wire _05700_;
	wire _05701_;
	wire _05702_;
	wire _05703_;
	wire _05704_;
	wire _05705_;
	wire _05706_;
	wire _05707_;
	wire _05708_;
	wire _05709_;
	wire _05710_;
	wire _05711_;
	wire _05712_;
	wire _05713_;
	wire _05714_;
	wire _05715_;
	wire _05716_;
	wire _05717_;
	wire _05718_;
	wire _05719_;
	wire _05720_;
	wire _05721_;
	wire _05722_;
	wire _05723_;
	wire _05724_;
	wire _05725_;
	wire _05726_;
	wire _05727_;
	wire _05728_;
	wire _05729_;
	wire _05730_;
	wire _05731_;
	wire _05732_;
	wire _05733_;
	wire _05734_;
	wire _05735_;
	wire _05736_;
	wire _05737_;
	wire _05738_;
	wire _05739_;
	wire _05740_;
	wire _05741_;
	wire _05742_;
	wire _05743_;
	wire _05744_;
	wire _05745_;
	wire _05746_;
	wire _05747_;
	wire _05748_;
	wire _05749_;
	wire _05750_;
	wire _05751_;
	wire _05752_;
	wire _05753_;
	wire _05754_;
	wire _05755_;
	wire _05756_;
	wire _05757_;
	wire _05758_;
	wire _05759_;
	wire _05760_;
	wire _05761_;
	wire _05762_;
	wire _05763_;
	wire _05764_;
	wire _05765_;
	wire _05766_;
	wire _05767_;
	wire _05768_;
	wire _05769_;
	wire _05770_;
	wire _05771_;
	wire _05772_;
	wire _05773_;
	wire _05774_;
	wire _05775_;
	wire _05776_;
	wire _05777_;
	wire _05778_;
	wire _05779_;
	wire _05780_;
	wire _05781_;
	wire _05782_;
	wire _05783_;
	wire _05784_;
	wire _05785_;
	wire _05786_;
	wire _05787_;
	wire _05788_;
	wire _05789_;
	wire _05790_;
	wire _05791_;
	wire _05792_;
	wire _05793_;
	wire _05794_;
	wire _05795_;
	wire _05796_;
	wire _05797_;
	wire _05798_;
	wire _05799_;
	wire _05800_;
	wire _05801_;
	wire _05802_;
	wire _05803_;
	wire _05804_;
	wire _05805_;
	wire _05806_;
	wire _05807_;
	wire _05808_;
	wire _05809_;
	wire _05810_;
	wire _05811_;
	wire _05812_;
	wire _05813_;
	wire _05814_;
	wire _05815_;
	wire _05816_;
	wire _05817_;
	wire _05818_;
	wire _05819_;
	wire _05820_;
	wire _05821_;
	wire _05822_;
	wire _05823_;
	wire _05824_;
	wire _05825_;
	wire _05826_;
	wire _05827_;
	wire _05828_;
	wire _05829_;
	wire _05830_;
	wire _05831_;
	wire _05832_;
	wire _05833_;
	wire _05834_;
	wire _05835_;
	wire _05836_;
	wire _05837_;
	wire _05838_;
	wire _05839_;
	wire _05840_;
	wire _05841_;
	wire _05842_;
	wire _05843_;
	wire _05844_;
	wire _05845_;
	wire _05846_;
	wire _05847_;
	wire _05848_;
	wire _05849_;
	wire _05850_;
	wire _05851_;
	wire _05852_;
	wire _05853_;
	wire _05854_;
	wire _05855_;
	wire _05856_;
	wire _05857_;
	wire _05858_;
	wire _05859_;
	wire _05860_;
	wire _05861_;
	wire _05862_;
	wire _05863_;
	wire _05864_;
	wire _05865_;
	wire _05866_;
	wire _05867_;
	wire _05868_;
	wire _05869_;
	wire _05870_;
	wire _05871_;
	wire _05872_;
	wire _05873_;
	wire _05874_;
	wire _05875_;
	wire _05876_;
	wire _05877_;
	wire _05878_;
	wire _05879_;
	wire _05880_;
	wire _05881_;
	wire _05882_;
	wire _05883_;
	wire _05884_;
	wire _05885_;
	wire _05886_;
	wire _05887_;
	wire _05888_;
	wire _05889_;
	wire _05890_;
	wire _05891_;
	wire _05892_;
	wire _05893_;
	wire _05894_;
	wire _05895_;
	wire _05896_;
	wire _05897_;
	wire _05898_;
	wire _05899_;
	wire _05900_;
	wire _05901_;
	wire _05902_;
	wire _05903_;
	wire _05904_;
	wire _05905_;
	wire _05906_;
	wire _05907_;
	wire _05908_;
	wire _05909_;
	wire _05910_;
	wire _05911_;
	wire _05912_;
	wire _05913_;
	wire _05914_;
	wire _05915_;
	wire _05916_;
	wire _05917_;
	wire _05918_;
	wire _05919_;
	wire _05920_;
	wire _05921_;
	wire _05922_;
	wire _05923_;
	wire _05924_;
	wire _05925_;
	wire _05926_;
	wire _05927_;
	wire _05928_;
	wire _05929_;
	wire _05930_;
	wire _05931_;
	wire _05932_;
	wire _05933_;
	wire _05934_;
	wire _05935_;
	wire _05936_;
	wire _05937_;
	wire _05938_;
	wire _05939_;
	wire _05940_;
	wire _05941_;
	wire _05942_;
	wire _05943_;
	wire _05944_;
	wire _05945_;
	wire _05946_;
	wire _05947_;
	wire _05948_;
	wire _05949_;
	wire _05950_;
	wire _05951_;
	wire _05952_;
	wire _05953_;
	wire _05954_;
	wire _05955_;
	wire _05956_;
	wire _05957_;
	wire _05958_;
	wire _05959_;
	wire _05960_;
	wire _05961_;
	wire _05962_;
	wire _05963_;
	wire _05964_;
	wire _05965_;
	wire _05966_;
	wire _05967_;
	wire _05968_;
	wire _05969_;
	wire _05970_;
	wire _05971_;
	wire _05972_;
	wire _05973_;
	wire _05974_;
	wire _05975_;
	wire _05976_;
	wire _05977_;
	wire _05978_;
	wire _05979_;
	wire _05980_;
	wire _05981_;
	wire _05982_;
	wire _05983_;
	wire _05984_;
	wire _05985_;
	wire _05986_;
	wire _05987_;
	wire _05988_;
	wire _05989_;
	wire _05990_;
	wire _05991_;
	wire _05992_;
	wire _05993_;
	wire _05994_;
	wire _05995_;
	wire _05996_;
	wire _05997_;
	wire _05998_;
	wire _05999_;
	wire _06000_;
	wire _06001_;
	wire _06002_;
	wire _06003_;
	wire _06004_;
	wire _06005_;
	wire _06006_;
	wire _06007_;
	wire _06008_;
	wire _06009_;
	wire _06010_;
	wire _06011_;
	wire _06012_;
	wire _06013_;
	wire _06014_;
	wire _06015_;
	wire _06016_;
	wire _06017_;
	wire _06018_;
	wire _06019_;
	wire _06020_;
	wire _06021_;
	wire _06022_;
	wire _06023_;
	wire _06024_;
	wire _06025_;
	wire _06026_;
	wire _06027_;
	wire _06028_;
	wire _06029_;
	wire _06030_;
	wire _06031_;
	wire _06032_;
	wire _06033_;
	wire _06034_;
	wire _06035_;
	wire _06036_;
	wire _06037_;
	wire _06038_;
	wire _06039_;
	wire _06040_;
	wire _06041_;
	wire _06042_;
	wire _06043_;
	wire _06044_;
	wire _06045_;
	wire _06046_;
	wire _06047_;
	wire _06048_;
	wire _06049_;
	wire _06050_;
	wire _06051_;
	wire _06052_;
	wire _06053_;
	wire _06054_;
	wire _06055_;
	wire _06056_;
	wire _06057_;
	wire _06058_;
	wire _06059_;
	wire _06060_;
	wire [9:0] _06061_;
	wire [22:0] _06062_;
	wire [22:0] _06063_;
	wire [22:0] _06064_;
	wire [22:0] _06065_;
	wire [9:0] _06066_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire \mchip.design.HS ;
	wire [1:0] \mchip.design.VGA_Blue ;
	wire [1:0] \mchip.design.VGA_Green ;
	wire [1:0] \mchip.design.VGA_Red ;
	wire \mchip.design.VS ;
	wire \mchip.design.blank ;
	wire [9:0] \mchip.design.board.col ;
	wire \mchip.design.board.is_board ;
	wire [8:0] \mchip.design.board.level_0_H.high ;
	wire [8:0] \mchip.design.board.level_0_H.low ;
	wire [8:0] \mchip.design.board.level_0_H.val ;
	wire [9:0] \mchip.design.board.level_0_V.high ;
	wire [9:0] \mchip.design.board.level_0_V.low ;
	wire [9:0] \mchip.design.board.level_0_V.val ;
	wire [8:0] \mchip.design.board.level_1_H.high ;
	wire [8:0] \mchip.design.board.level_1_H.low ;
	wire [8:0] \mchip.design.board.level_1_H.val ;
	wire [9:0] \mchip.design.board.level_1_V.high ;
	wire [9:0] \mchip.design.board.level_1_V.low ;
	wire [9:0] \mchip.design.board.level_1_V.val ;
	wire [8:0] \mchip.design.board.level_2_H.high ;
	wire [8:0] \mchip.design.board.level_2_H.low ;
	wire [8:0] \mchip.design.board.level_2_H.val ;
	wire [9:0] \mchip.design.board.level_2_V.high ;
	wire [9:0] \mchip.design.board.level_2_V.low ;
	wire [9:0] \mchip.design.board.level_2_V.val ;
	wire [8:0] \mchip.design.board.level_3_H.high ;
	wire [8:0] \mchip.design.board.level_3_H.low ;
	wire [8:0] \mchip.design.board.level_3_H.val ;
	wire [9:0] \mchip.design.board.level_3_V.high ;
	wire [9:0] \mchip.design.board.level_3_V.low ;
	wire [9:0] \mchip.design.board.level_3_V.val ;
	wire [8:0] \mchip.design.board.level_4_H.high ;
	wire [8:0] \mchip.design.board.level_4_H.low ;
	wire [8:0] \mchip.design.board.level_4_H.val ;
	wire [9:0] \mchip.design.board.level_4_V.high ;
	wire [9:0] \mchip.design.board.level_4_V.low ;
	wire [9:0] \mchip.design.board.level_4_V.val ;
	wire [8:0] \mchip.design.board.level_5_H.high ;
	wire [8:0] \mchip.design.board.level_5_H.low ;
	wire [8:0] \mchip.design.board.level_5_H.val ;
	wire [9:0] \mchip.design.board.level_5_V.high ;
	wire [9:0] \mchip.design.board.level_5_V.low ;
	wire [9:0] \mchip.design.board.level_5_V.val ;
	wire [8:0] \mchip.design.board.level_6_H.high ;
	wire [8:0] \mchip.design.board.level_6_H.low ;
	wire [8:0] \mchip.design.board.level_6_H.val ;
	wire [9:0] \mchip.design.board.level_6_V.high ;
	wire [9:0] \mchip.design.board.level_6_V.low ;
	wire [9:0] \mchip.design.board.level_6_V.val ;
	wire [9:0] \mchip.design.board.level_7_V.high ;
	wire [9:0] \mchip.design.board.level_7_V.low ;
	wire [9:0] \mchip.design.board.level_7_V.val ;
	wire [8:0] \mchip.design.board.row ;
	wire \mchip.design.bot_confirm ;
	wire \mchip.design.clock ;
	wire [9:0] \mchip.design.colFromVGA ;
	wire [9:0] \mchip.design.colToModule ;
	wire [1:0] \mchip.design.colors.blue ;
	wire \mchip.design.colors.clock ;
	wire [6:0] \mchip.design.colors.currentTokenCol ;
	wire [5:0] \mchip.design.colors.currentTokenRow ;
	wire [1:0] \mchip.design.colors.green ;
	wire \mchip.design.colors.is_board ;
	wire [1:0] \mchip.design.colors.red ;
	wire \mchip.design.colors.reset ;
	wire [83:0] \mchip.design.colors.tokens ;
	reg [2:0] \mchip.design.currStateConfirm ;
	wire \mchip.design.debounceClear ;
	reg [22:0] \mchip.design.debounceCount ;
	wire \mchip.design.debounceCountEn ;
	wire [22:0] \mchip.design.debounceLimit ;
	wire \mchip.design.inputChangeDebug ;
	wire \mchip.design.inputConfirm ;
	reg \mchip.design.inputConfirmHalf ;
	wire \mchip.design.inputConfirmLimited ;
	reg \mchip.design.inputConfirmSync ;
	wire [6:0] \mchip.design.inputMoves ;
	reg [6:0] \mchip.design.inputMovesHalf ;
	reg [6:0] \mchip.design.inputMovesSync ;
	wire \mchip.design.inputNewGame ;
	reg \mchip.design.inputNewGameHalf ;
	reg \mchip.design.inputNewGameSync ;
	wire \mchip.design.inputSwitchPVP ;
	reg \mchip.design.inputSwitchPVPHalf ;
	reg \mchip.design.inputSwitchPVPSync ;
	wire \mchip.design.inputSwitchPlayer ;
	reg \mchip.design.inputSwitchPlayerHalf ;
	reg \mchip.design.inputSwitchPlayerSync ;
	wire \mchip.design.is_board ;
	wire [11:0] \mchip.design.outputs ;
	wire \mchip.design.owner.clock ;
	wire \mchip.design.owner.currentPlayer ;
	wire \mchip.design.owner.fsm.clock ;
	reg \mchip.design.owner.fsm.currState ;
	wire \mchip.design.owner.fsm.currentPlayer ;
	wire \mchip.design.owner.fsm.nextState ;
	wire \mchip.design.owner.fsm.reset ;
	wire \mchip.design.owner.fsm.switchTurn ;
	wire [6:0] \mchip.design.owner.move ;
	wire \mchip.design.owner.newGame ;
	wire \mchip.design.owner.player_1_confirm ;
	wire [6:0] \mchip.design.owner.player_1_input ;
	wire \mchip.design.owner.reset ;
	wire \mchip.design.owner.switchTurn ;
	reg [83:0] \mchip.design.owner.tokens ;
	wire \mchip.design.pve.bot_confirm ;
	wire \mchip.design.pve.bot_turn ;
	wire \mchip.design.pve.clock ;
	wire \mchip.design.pve.fsm.bot_confirm ;
	wire \mchip.design.pve.fsm.bot_turn ;
	wire \mchip.design.pve.fsm.clock ;
	reg [2:0] \mchip.design.pve.fsm.currState ;
	wire \mchip.design.pve.fsm.reset ;
	wire [6:0] \mchip.design.pve.fsm.selectedMove ;
	reg [22:0] \mchip.design.pve.fsm.timeOut ;
	wire [22:0] \mchip.design.pve.fsm.timeOutDelay ;
	wire \mchip.design.pve.fsm.timeOutEn ;
	wire \mchip.design.pve.rand0.clock ;
	wire [3:0] \mchip.design.pve.rand0.inputFF ;
	reg [3:0] \mchip.design.pve.rand0.outputFF ;
	wire \mchip.design.pve.rand0.randomOut ;
	wire \mchip.design.pve.rand0.reset ;
	wire \mchip.design.pve.rand1.clock ;
	wire [3:0] \mchip.design.pve.rand1.inputFF ;
	reg [3:0] \mchip.design.pve.rand1.outputFF ;
	wire \mchip.design.pve.rand1.randomOut ;
	wire \mchip.design.pve.rand1.reset ;
	wire \mchip.design.pve.rand2.clock ;
	wire [3:0] \mchip.design.pve.rand2.inputFF ;
	reg [3:0] \mchip.design.pve.rand2.outputFF ;
	wire \mchip.design.pve.rand2.randomOut ;
	wire \mchip.design.pve.rand2.reset ;
	wire \mchip.design.pve.rand3.clock ;
	wire [3:0] \mchip.design.pve.rand3.inputFF ;
	reg [3:0] \mchip.design.pve.rand3.outputFF ;
	wire \mchip.design.pve.rand3.randomOut ;
	wire \mchip.design.pve.rand3.reset ;
	wire \mchip.design.pve.rand4.clock ;
	wire [3:0] \mchip.design.pve.rand4.inputFF ;
	reg [3:0] \mchip.design.pve.rand4.outputFF ;
	wire \mchip.design.pve.rand4.randomOut ;
	wire \mchip.design.pve.rand4.reset ;
	wire \mchip.design.pve.rand5.clock ;
	wire [3:0] \mchip.design.pve.rand5.inputFF ;
	reg [3:0] \mchip.design.pve.rand5.outputFF ;
	wire \mchip.design.pve.rand5.randomOut ;
	wire \mchip.design.pve.rand5.reset ;
	wire \mchip.design.pve.rand6.clock ;
	wire [3:0] \mchip.design.pve.rand6.inputFF ;
	reg [3:0] \mchip.design.pve.rand6.outputFF ;
	wire \mchip.design.pve.rand6.randomOut ;
	wire \mchip.design.pve.rand6.reset ;
	wire [6:0] \mchip.design.pve.random ;
	wire \mchip.design.pve.reset ;
	wire [83:0] \mchip.design.pve.tokens ;
	wire \mchip.design.reset ;
	wire [8:0] \mchip.design.rowFromVGA ;
	wire [8:0] \mchip.design.rowToModule ;
	wire [9:0] \mchip.design.token.col ;
	wire [9:0] \mchip.design.token.level_0_H_0.high ;
	wire [9:0] \mchip.design.token.level_0_H_0.low ;
	wire [9:0] \mchip.design.token.level_0_H_0.val ;
	wire [9:0] \mchip.design.token.level_0_H_14.high ;
	wire [9:0] \mchip.design.token.level_0_H_14.low ;
	wire [9:0] \mchip.design.token.level_0_H_14.val ;
	wire [9:0] \mchip.design.token.level_0_H_21.high ;
	wire [9:0] \mchip.design.token.level_0_H_21.low ;
	wire [9:0] \mchip.design.token.level_0_H_21.val ;
	wire [9:0] \mchip.design.token.level_0_H_28.high ;
	wire [9:0] \mchip.design.token.level_0_H_28.low ;
	wire [9:0] \mchip.design.token.level_0_H_28.val ;
	wire [9:0] \mchip.design.token.level_0_H_35.high ;
	wire [9:0] \mchip.design.token.level_0_H_35.low ;
	wire [9:0] \mchip.design.token.level_0_H_35.val ;
	wire [9:0] \mchip.design.token.level_0_H_7.high ;
	wire [9:0] \mchip.design.token.level_0_H_7.low ;
	wire [9:0] \mchip.design.token.level_0_H_7.val ;
	wire [8:0] \mchip.design.token.level_0_V_0.high ;
	wire [8:0] \mchip.design.token.level_0_V_0.low ;
	wire [8:0] \mchip.design.token.level_0_V_0.val ;
	wire [8:0] \mchip.design.token.level_0_V_1.high ;
	wire [8:0] \mchip.design.token.level_0_V_1.low ;
	wire [8:0] \mchip.design.token.level_0_V_1.val ;
	wire [8:0] \mchip.design.token.level_0_V_2.high ;
	wire [8:0] \mchip.design.token.level_0_V_2.low ;
	wire [8:0] \mchip.design.token.level_0_V_2.val ;
	wire [8:0] \mchip.design.token.level_0_V_3.high ;
	wire [8:0] \mchip.design.token.level_0_V_3.low ;
	wire [8:0] \mchip.design.token.level_0_V_3.val ;
	wire [8:0] \mchip.design.token.level_0_V_4.high ;
	wire [8:0] \mchip.design.token.level_0_V_4.low ;
	wire [8:0] \mchip.design.token.level_0_V_4.val ;
	wire [8:0] \mchip.design.token.level_0_V_5.high ;
	wire [8:0] \mchip.design.token.level_0_V_5.low ;
	wire [8:0] \mchip.design.token.level_0_V_5.val ;
	wire [8:0] \mchip.design.token.level_0_V_6.high ;
	wire [8:0] \mchip.design.token.level_0_V_6.low ;
	wire [8:0] \mchip.design.token.level_0_V_6.val ;
	wire [9:0] \mchip.design.token.level_1_H_1.high ;
	wire [9:0] \mchip.design.token.level_1_H_1.low ;
	wire [9:0] \mchip.design.token.level_1_H_1.val ;
	wire [9:0] \mchip.design.token.level_1_H_15.high ;
	wire [9:0] \mchip.design.token.level_1_H_15.low ;
	wire [9:0] \mchip.design.token.level_1_H_15.val ;
	wire [9:0] \mchip.design.token.level_1_H_22.high ;
	wire [9:0] \mchip.design.token.level_1_H_22.low ;
	wire [9:0] \mchip.design.token.level_1_H_22.val ;
	wire [9:0] \mchip.design.token.level_1_H_29.high ;
	wire [9:0] \mchip.design.token.level_1_H_29.low ;
	wire [9:0] \mchip.design.token.level_1_H_29.val ;
	wire [9:0] \mchip.design.token.level_1_H_36.high ;
	wire [9:0] \mchip.design.token.level_1_H_36.low ;
	wire [9:0] \mchip.design.token.level_1_H_36.val ;
	wire [9:0] \mchip.design.token.level_1_H_8.high ;
	wire [9:0] \mchip.design.token.level_1_H_8.low ;
	wire [9:0] \mchip.design.token.level_1_H_8.val ;
	wire [8:0] \mchip.design.token.level_1_V_10.high ;
	wire [8:0] \mchip.design.token.level_1_V_10.low ;
	wire [8:0] \mchip.design.token.level_1_V_10.val ;
	wire [8:0] \mchip.design.token.level_1_V_11.high ;
	wire [8:0] \mchip.design.token.level_1_V_11.low ;
	wire [8:0] \mchip.design.token.level_1_V_11.val ;
	wire [8:0] \mchip.design.token.level_1_V_12.high ;
	wire [8:0] \mchip.design.token.level_1_V_12.low ;
	wire [8:0] \mchip.design.token.level_1_V_12.val ;
	wire [8:0] \mchip.design.token.level_1_V_13.high ;
	wire [8:0] \mchip.design.token.level_1_V_13.low ;
	wire [8:0] \mchip.design.token.level_1_V_13.val ;
	wire [8:0] \mchip.design.token.level_1_V_7.high ;
	wire [8:0] \mchip.design.token.level_1_V_7.low ;
	wire [8:0] \mchip.design.token.level_1_V_7.val ;
	wire [8:0] \mchip.design.token.level_1_V_8.high ;
	wire [8:0] \mchip.design.token.level_1_V_8.low ;
	wire [8:0] \mchip.design.token.level_1_V_8.val ;
	wire [8:0] \mchip.design.token.level_1_V_9.high ;
	wire [8:0] \mchip.design.token.level_1_V_9.low ;
	wire [8:0] \mchip.design.token.level_1_V_9.val ;
	wire [9:0] \mchip.design.token.level_2_H_16.high ;
	wire [9:0] \mchip.design.token.level_2_H_16.low ;
	wire [9:0] \mchip.design.token.level_2_H_16.val ;
	wire [9:0] \mchip.design.token.level_2_H_2.high ;
	wire [9:0] \mchip.design.token.level_2_H_2.low ;
	wire [9:0] \mchip.design.token.level_2_H_2.val ;
	wire [9:0] \mchip.design.token.level_2_H_23.high ;
	wire [9:0] \mchip.design.token.level_2_H_23.low ;
	wire [9:0] \mchip.design.token.level_2_H_23.val ;
	wire [9:0] \mchip.design.token.level_2_H_30.high ;
	wire [9:0] \mchip.design.token.level_2_H_30.low ;
	wire [9:0] \mchip.design.token.level_2_H_30.val ;
	wire [9:0] \mchip.design.token.level_2_H_37.high ;
	wire [9:0] \mchip.design.token.level_2_H_37.low ;
	wire [9:0] \mchip.design.token.level_2_H_37.val ;
	wire [9:0] \mchip.design.token.level_2_H_9.high ;
	wire [9:0] \mchip.design.token.level_2_H_9.low ;
	wire [9:0] \mchip.design.token.level_2_H_9.val ;
	wire [8:0] \mchip.design.token.level_2_V_14.high ;
	wire [8:0] \mchip.design.token.level_2_V_14.low ;
	wire [8:0] \mchip.design.token.level_2_V_14.val ;
	wire [8:0] \mchip.design.token.level_2_V_15.high ;
	wire [8:0] \mchip.design.token.level_2_V_15.low ;
	wire [8:0] \mchip.design.token.level_2_V_15.val ;
	wire [8:0] \mchip.design.token.level_2_V_16.high ;
	wire [8:0] \mchip.design.token.level_2_V_16.low ;
	wire [8:0] \mchip.design.token.level_2_V_16.val ;
	wire [8:0] \mchip.design.token.level_2_V_17.high ;
	wire [8:0] \mchip.design.token.level_2_V_17.low ;
	wire [8:0] \mchip.design.token.level_2_V_17.val ;
	wire [8:0] \mchip.design.token.level_2_V_18.high ;
	wire [8:0] \mchip.design.token.level_2_V_18.low ;
	wire [8:0] \mchip.design.token.level_2_V_18.val ;
	wire [8:0] \mchip.design.token.level_2_V_19.high ;
	wire [8:0] \mchip.design.token.level_2_V_19.low ;
	wire [8:0] \mchip.design.token.level_2_V_19.val ;
	wire [8:0] \mchip.design.token.level_2_V_20.high ;
	wire [8:0] \mchip.design.token.level_2_V_20.low ;
	wire [8:0] \mchip.design.token.level_2_V_20.val ;
	wire [9:0] \mchip.design.token.level_3_H_10.high ;
	wire [9:0] \mchip.design.token.level_3_H_10.low ;
	wire [9:0] \mchip.design.token.level_3_H_10.val ;
	wire [9:0] \mchip.design.token.level_3_H_17.high ;
	wire [9:0] \mchip.design.token.level_3_H_17.low ;
	wire [9:0] \mchip.design.token.level_3_H_17.val ;
	wire [9:0] \mchip.design.token.level_3_H_24.high ;
	wire [9:0] \mchip.design.token.level_3_H_24.low ;
	wire [9:0] \mchip.design.token.level_3_H_24.val ;
	wire [9:0] \mchip.design.token.level_3_H_3.high ;
	wire [9:0] \mchip.design.token.level_3_H_3.low ;
	wire [9:0] \mchip.design.token.level_3_H_3.val ;
	wire [9:0] \mchip.design.token.level_3_H_31.high ;
	wire [9:0] \mchip.design.token.level_3_H_31.low ;
	wire [9:0] \mchip.design.token.level_3_H_31.val ;
	wire [9:0] \mchip.design.token.level_3_H_38.high ;
	wire [9:0] \mchip.design.token.level_3_H_38.low ;
	wire [9:0] \mchip.design.token.level_3_H_38.val ;
	wire [8:0] \mchip.design.token.level_3_V_21.high ;
	wire [8:0] \mchip.design.token.level_3_V_21.low ;
	wire [8:0] \mchip.design.token.level_3_V_21.val ;
	wire [8:0] \mchip.design.token.level_3_V_22.high ;
	wire [8:0] \mchip.design.token.level_3_V_22.low ;
	wire [8:0] \mchip.design.token.level_3_V_22.val ;
	wire [8:0] \mchip.design.token.level_3_V_23.high ;
	wire [8:0] \mchip.design.token.level_3_V_23.low ;
	wire [8:0] \mchip.design.token.level_3_V_23.val ;
	wire [8:0] \mchip.design.token.level_3_V_24.high ;
	wire [8:0] \mchip.design.token.level_3_V_24.low ;
	wire [8:0] \mchip.design.token.level_3_V_24.val ;
	wire [8:0] \mchip.design.token.level_3_V_25.high ;
	wire [8:0] \mchip.design.token.level_3_V_25.low ;
	wire [8:0] \mchip.design.token.level_3_V_25.val ;
	wire [8:0] \mchip.design.token.level_3_V_26.high ;
	wire [8:0] \mchip.design.token.level_3_V_26.low ;
	wire [8:0] \mchip.design.token.level_3_V_26.val ;
	wire [8:0] \mchip.design.token.level_3_V_27.high ;
	wire [8:0] \mchip.design.token.level_3_V_27.low ;
	wire [8:0] \mchip.design.token.level_3_V_27.val ;
	wire [9:0] \mchip.design.token.level_4_H_11.high ;
	wire [9:0] \mchip.design.token.level_4_H_11.low ;
	wire [9:0] \mchip.design.token.level_4_H_11.val ;
	wire [9:0] \mchip.design.token.level_4_H_18.high ;
	wire [9:0] \mchip.design.token.level_4_H_18.low ;
	wire [9:0] \mchip.design.token.level_4_H_18.val ;
	wire [9:0] \mchip.design.token.level_4_H_25.high ;
	wire [9:0] \mchip.design.token.level_4_H_25.low ;
	wire [9:0] \mchip.design.token.level_4_H_25.val ;
	wire [9:0] \mchip.design.token.level_4_H_32.high ;
	wire [9:0] \mchip.design.token.level_4_H_32.low ;
	wire [9:0] \mchip.design.token.level_4_H_32.val ;
	wire [9:0] \mchip.design.token.level_4_H_39.high ;
	wire [9:0] \mchip.design.token.level_4_H_39.low ;
	wire [9:0] \mchip.design.token.level_4_H_39.val ;
	wire [9:0] \mchip.design.token.level_4_H_4.high ;
	wire [9:0] \mchip.design.token.level_4_H_4.low ;
	wire [9:0] \mchip.design.token.level_4_H_4.val ;
	wire [8:0] \mchip.design.token.level_4_V_28.high ;
	wire [8:0] \mchip.design.token.level_4_V_28.low ;
	wire [8:0] \mchip.design.token.level_4_V_28.val ;
	wire [8:0] \mchip.design.token.level_4_V_29.high ;
	wire [8:0] \mchip.design.token.level_4_V_29.low ;
	wire [8:0] \mchip.design.token.level_4_V_29.val ;
	wire [8:0] \mchip.design.token.level_4_V_30.high ;
	wire [8:0] \mchip.design.token.level_4_V_30.low ;
	wire [8:0] \mchip.design.token.level_4_V_30.val ;
	wire [8:0] \mchip.design.token.level_4_V_31.high ;
	wire [8:0] \mchip.design.token.level_4_V_31.low ;
	wire [8:0] \mchip.design.token.level_4_V_31.val ;
	wire [8:0] \mchip.design.token.level_4_V_32.high ;
	wire [8:0] \mchip.design.token.level_4_V_32.low ;
	wire [8:0] \mchip.design.token.level_4_V_32.val ;
	wire [8:0] \mchip.design.token.level_4_V_33.high ;
	wire [8:0] \mchip.design.token.level_4_V_33.low ;
	wire [8:0] \mchip.design.token.level_4_V_33.val ;
	wire [8:0] \mchip.design.token.level_4_V_34.high ;
	wire [8:0] \mchip.design.token.level_4_V_34.low ;
	wire [8:0] \mchip.design.token.level_4_V_34.val ;
	wire [9:0] \mchip.design.token.level_5_H_12.high ;
	wire [9:0] \mchip.design.token.level_5_H_12.low ;
	wire [9:0] \mchip.design.token.level_5_H_12.val ;
	wire [9:0] \mchip.design.token.level_5_H_19.high ;
	wire [9:0] \mchip.design.token.level_5_H_19.low ;
	wire [9:0] \mchip.design.token.level_5_H_19.val ;
	wire [9:0] \mchip.design.token.level_5_H_26.high ;
	wire [9:0] \mchip.design.token.level_5_H_26.low ;
	wire [9:0] \mchip.design.token.level_5_H_26.val ;
	wire [9:0] \mchip.design.token.level_5_H_33.high ;
	wire [9:0] \mchip.design.token.level_5_H_33.low ;
	wire [9:0] \mchip.design.token.level_5_H_33.val ;
	wire [9:0] \mchip.design.token.level_5_H_40.high ;
	wire [9:0] \mchip.design.token.level_5_H_40.low ;
	wire [9:0] \mchip.design.token.level_5_H_40.val ;
	wire [9:0] \mchip.design.token.level_5_H_5.high ;
	wire [9:0] \mchip.design.token.level_5_H_5.low ;
	wire [9:0] \mchip.design.token.level_5_H_5.val ;
	wire [8:0] \mchip.design.token.level_5_V_35.high ;
	wire [8:0] \mchip.design.token.level_5_V_35.low ;
	wire [8:0] \mchip.design.token.level_5_V_35.val ;
	wire [8:0] \mchip.design.token.level_5_V_36.high ;
	wire [8:0] \mchip.design.token.level_5_V_36.low ;
	wire [8:0] \mchip.design.token.level_5_V_36.val ;
	wire [8:0] \mchip.design.token.level_5_V_37.high ;
	wire [8:0] \mchip.design.token.level_5_V_37.low ;
	wire [8:0] \mchip.design.token.level_5_V_37.val ;
	wire [8:0] \mchip.design.token.level_5_V_38.high ;
	wire [8:0] \mchip.design.token.level_5_V_38.low ;
	wire [8:0] \mchip.design.token.level_5_V_38.val ;
	wire [8:0] \mchip.design.token.level_5_V_39.high ;
	wire [8:0] \mchip.design.token.level_5_V_39.low ;
	wire [8:0] \mchip.design.token.level_5_V_39.val ;
	wire [8:0] \mchip.design.token.level_5_V_40.high ;
	wire [8:0] \mchip.design.token.level_5_V_40.low ;
	wire [8:0] \mchip.design.token.level_5_V_40.val ;
	wire [8:0] \mchip.design.token.level_5_V_41.high ;
	wire [8:0] \mchip.design.token.level_5_V_41.low ;
	wire [8:0] \mchip.design.token.level_5_V_41.val ;
	wire [9:0] \mchip.design.token.level_6_H_13.high ;
	wire [9:0] \mchip.design.token.level_6_H_13.low ;
	wire [9:0] \mchip.design.token.level_6_H_13.val ;
	wire [9:0] \mchip.design.token.level_6_H_20.high ;
	wire [9:0] \mchip.design.token.level_6_H_20.low ;
	wire [9:0] \mchip.design.token.level_6_H_20.val ;
	wire [9:0] \mchip.design.token.level_6_H_27.high ;
	wire [9:0] \mchip.design.token.level_6_H_27.low ;
	wire [9:0] \mchip.design.token.level_6_H_27.val ;
	wire [9:0] \mchip.design.token.level_6_H_34.high ;
	wire [9:0] \mchip.design.token.level_6_H_34.low ;
	wire [9:0] \mchip.design.token.level_6_H_34.val ;
	wire [9:0] \mchip.design.token.level_6_H_41.high ;
	wire [9:0] \mchip.design.token.level_6_H_41.low ;
	wire [9:0] \mchip.design.token.level_6_H_41.val ;
	wire [9:0] \mchip.design.token.level_6_H_6.high ;
	wire [9:0] \mchip.design.token.level_6_H_6.low ;
	wire [9:0] \mchip.design.token.level_6_H_6.val ;
	wire [8:0] \mchip.design.token.row ;
	wire [83:0] \mchip.design.tokens ;
	wire \mchip.design.vga.clk ;
	reg [9:0] \mchip.design.vga.h_idx ;
	reg \mchip.design.vga.hsync ;
	wire \mchip.design.vga.rst ;
	reg [9:0] \mchip.design.vga.v_idx ;
	wire \mchip.design.vga.valid ;
	reg \mchip.design.vga.vsync ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _06064_[0] = ~\mchip.design.pve.fsm.timeOut [0];
	assign _02661_ = ~\mchip.design.inputSwitchPlayerSync ;
	assign _02671_ = \mchip.design.pve.fsm.timeOut [20] & ~\mchip.design.pve.fsm.timeOut [21];
	assign _02682_ = ~(_02671_ & \mchip.design.pve.fsm.timeOut [22]);
	assign _02693_ = \mchip.design.pve.fsm.timeOut [16] & \mchip.design.pve.fsm.timeOut [17];
	assign _02704_ = \mchip.design.pve.fsm.timeOut [18] & \mchip.design.pve.fsm.timeOut [19];
	assign _02715_ = ~(_02704_ & _02693_);
	assign _02726_ = _02715_ | _02682_;
	assign _02737_ = \mchip.design.pve.fsm.timeOut [10] & \mchip.design.pve.fsm.timeOut [11];
	assign _02747_ = \mchip.design.pve.fsm.timeOut [8] | ~\mchip.design.pve.fsm.timeOut [9];
	assign _02758_ = _02737_ & ~_02747_;
	assign _02769_ = \mchip.design.pve.fsm.timeOut [13] | ~\mchip.design.pve.fsm.timeOut [12];
	assign _02780_ = \mchip.design.pve.fsm.timeOut [15] | ~\mchip.design.pve.fsm.timeOut [14];
	assign _02790_ = _02780_ | _02769_;
	assign _02801_ = _02790_ | ~_02758_;
	assign _02812_ = \mchip.design.pve.fsm.timeOut [4] & ~\mchip.design.pve.fsm.timeOut [5];
	assign _02823_ = ~(\mchip.design.pve.fsm.timeOut [6] | \mchip.design.pve.fsm.timeOut [7]);
	assign _02834_ = ~(_02823_ & _02812_);
	assign _02845_ = \mchip.design.pve.fsm.timeOut [2] | \mchip.design.pve.fsm.timeOut [3];
	assign _02855_ = \mchip.design.pve.fsm.timeOut [1] | \mchip.design.pve.fsm.timeOut [0];
	assign _02866_ = _02855_ | _02845_;
	assign _02877_ = _02866_ | _02834_;
	assign _02888_ = _02877_ | _02801_;
	assign _02899_ = _02888_ | _02726_;
	assign _02909_ = _02780_ | ~\mchip.design.pve.fsm.timeOut [13];
	assign _02920_ = _02909_ & ~\mchip.design.pve.fsm.timeOut [15];
	assign _02931_ = _02920_ | _02715_;
	assign _02942_ = ~(_02790_ | _02715_);
	assign _02953_ = ~(\mchip.design.pve.fsm.timeOut [9] & \mchip.design.pve.fsm.timeOut [8]);
	assign _02964_ = _02953_ | ~_02737_;
	assign _02974_ = \mchip.design.pve.fsm.timeOut [5] | \mchip.design.pve.fsm.timeOut [4];
	assign _02985_ = _02823_ & ~_02974_;
	assign _02996_ = _02758_ & ~_02985_;
	assign _03007_ = _02964_ & ~_02996_;
	assign _03017_ = _02942_ & ~_03007_;
	assign _03028_ = _02931_ & ~_03017_;
	assign _03039_ = _03028_ | ~_02671_;
	assign _03050_ = _03039_ & ~\mchip.design.pve.fsm.timeOut [21];
	assign _03061_ = \mchip.design.pve.fsm.timeOut [22] & ~_03050_;
	assign _03072_ = _02899_ & ~_03061_;
	assign _03083_ = _02661_ & ~_03072_;
	assign _03093_ = _03083_ | io_in[13];
	assign _03104_ = \mchip.design.pve.fsm.currState [1] & ~_03093_;
	assign _03115_ = \mchip.design.pve.fsm.currState [2] & ~io_in[13];
	assign _00005_ = _03115_ | _03104_;
	assign _03135_ = io_in[13] | ~_03083_;
	assign _03146_ = \mchip.design.pve.fsm.currState [1] & ~_03135_;
	assign _03157_ = \mchip.design.inputSwitchPlayerSync  | io_in[13];
	assign _03168_ = \mchip.design.pve.fsm.currState [0] & ~_03157_;
	assign _03179_ = _03168_ | _03146_;
	assign _03190_ = ~(\mchip.design.owner.tokens [76] | \mchip.design.owner.tokens [77]);
	assign _03200_ = ~(_03190_ & \mchip.design.pve.rand3.outputFF [3]);
	assign _03211_ = \mchip.design.inputSwitchPlayerSync  & ~_03200_;
	assign _03222_ = ~_03211_;
	assign _03233_ = ~(\mchip.design.owner.tokens [74] | \mchip.design.owner.tokens [75]);
	assign _03243_ = ~(_03233_ & \mchip.design.pve.rand4.outputFF [3]);
	assign _03254_ = _03243_ | _02661_;
	assign _03265_ = ~(\mchip.design.owner.tokens [70] | \mchip.design.owner.tokens [71]);
	assign _03276_ = ~(_03265_ & \mchip.design.pve.rand6.outputFF [3]);
	assign _03287_ = \mchip.design.inputSwitchPlayerSync  & ~_03276_;
	assign _03298_ = ~(\mchip.design.owner.tokens [82] | \mchip.design.owner.tokens [83]);
	assign _03309_ = ~(_03298_ & \mchip.design.pve.rand0.outputFF [3]);
	assign _03319_ = \mchip.design.inputSwitchPlayerSync  & ~_03309_;
	assign _03330_ = _03319_ | _03287_;
	assign _03341_ = ~(\mchip.design.owner.tokens [80] | \mchip.design.owner.tokens [81]);
	assign _03352_ = ~(_03341_ & \mchip.design.pve.rand1.outputFF [3]);
	assign _03362_ = \mchip.design.inputSwitchPlayerSync  & ~_03352_;
	assign _03373_ = ~(_03362_ | _03330_);
	assign _03384_ = ~(\mchip.design.owner.tokens [72] | \mchip.design.owner.tokens [73]);
	assign _03395_ = ~(_03384_ & \mchip.design.pve.rand5.outputFF [3]);
	assign _03406_ = _03395_ | _02661_;
	assign _03417_ = ~(_03406_ & _03373_);
	assign _03427_ = ~(\mchip.design.owner.tokens [78] | \mchip.design.owner.tokens [79]);
	assign _03438_ = ~(_03427_ & \mchip.design.pve.rand2.outputFF [3]);
	assign _03449_ = \mchip.design.inputSwitchPlayerSync  & ~_03438_;
	assign _03460_ = _03449_ | _03417_;
	assign _03471_ = _03460_ | ~_03254_;
	assign _03481_ = _03222_ & ~_03471_;
	assign _03492_ = ~_03449_;
	assign _03503_ = _03319_ & ~_03287_;
	assign _03514_ = _03503_ | _03362_;
	assign _03525_ = _03406_ & ~_03514_;
	assign _03535_ = _03492_ & ~_03525_;
	assign _03546_ = _03254_ & ~_03535_;
	assign _03557_ = _03222_ & ~_03546_;
	assign _03567_ = _03406_ & ~_03362_;
	assign _03578_ = _03567_ | _03449_;
	assign _03589_ = _03254_ & ~_03578_;
	assign _03600_ = _03589_ | _03211_;
	assign _03611_ = _03557_ | ~_03600_;
	assign _03622_ = _03287_ & ~_03362_;
	assign _03632_ = _03406_ & ~_03622_;
	assign _03643_ = _03492_ & ~_03632_;
	assign _03654_ = _03254_ & ~_03643_;
	assign _03664_ = _03654_ | _03211_;
	assign _03675_ = ~(_03664_ | _03611_);
	assign _03686_ = ~(_03675_ | _03481_);
	assign _03697_ = io_in[13] | ~\mchip.design.inputSwitchPlayerSync ;
	assign _03708_ = _03697_ | _03686_;
	assign _03718_ = \mchip.design.pve.fsm.currState [0] & ~_03708_;
	assign _03729_ = _03718_ | io_in[13];
	assign _00004_ = _03729_ | _03179_;
	assign _03750_ = \mchip.design.vga.h_idx [9] & \mchip.design.vga.h_idx [8];
	assign _03760_ = \mchip.design.vga.h_idx [6] | \mchip.design.vga.h_idx [7];
	assign _03771_ = \mchip.design.vga.h_idx [4] | ~\mchip.design.vga.h_idx [5];
	assign _03782_ = _03771_ | _03760_;
	assign _03793_ = \mchip.design.vga.h_idx [2] | \mchip.design.vga.h_idx [3];
	assign _03804_ = \mchip.design.vga.h_idx [0] | \mchip.design.vga.h_idx [1];
	assign _03814_ = _03804_ | _03793_;
	assign _03825_ = _03814_ | _03782_;
	assign _03836_ = _03750_ & ~_03825_;
	assign _03847_ = \mchip.design.vga.h_idx [8] & \mchip.design.vga.h_idx [7];
	assign _03857_ = \mchip.design.vga.h_idx [8] & ~\mchip.design.vga.h_idx [7];
	assign _03868_ = ~(\mchip.design.vga.h_idx [5] | \mchip.design.vga.h_idx [6]);
	assign _03879_ = _03868_ | ~_03857_;
	assign _03890_ = _03879_ & ~_03847_;
	assign _03901_ = \mchip.design.vga.h_idx [9] & ~_03890_;
	assign _03911_ = _03901_ & ~_03836_;
	assign _03922_ = _03911_ | io_in[13];
	assign _00007_ = _03922_ | _03836_;
	assign _00011_ = _03901_ | _03836_;
	assign _00010_ = io_in[13] | ~\mchip.design.currStateConfirm [2];
	assign _00009_ = \mchip.design.inputNewGameSync  | io_in[13];
	assign _00008_ = io_in[13] | ~\mchip.design.pve.fsm.currState [1];
	assign _03992_ = \mchip.design.inputMovesSync [1] | \mchip.design.inputMovesSync [0];
	assign _04002_ = \mchip.design.inputMovesSync [3] | \mchip.design.inputMovesSync [2];
	assign _04013_ = ~(_04002_ | _03992_);
	assign _04024_ = \mchip.design.inputMovesSync [4] | ~\mchip.design.inputMovesSync [5];
	assign _04034_ = _04024_ | \mchip.design.inputMovesSync [6];
	assign _04045_ = _04013_ & ~_04034_;
	assign _04056_ = ~\mchip.design.inputMovesSync [6];
	assign _04067_ = \mchip.design.inputMovesSync [5] | \mchip.design.inputMovesSync [4];
	assign _04078_ = _04067_ | _04056_;
	assign _04089_ = _04013_ & ~_04078_;
	assign _04099_ = ~(_04089_ | _04045_);
	assign _04110_ = \mchip.design.inputMovesSync [5] | ~\mchip.design.inputMovesSync [4];
	assign _04121_ = _04110_ | \mchip.design.inputMovesSync [6];
	assign _04131_ = _04013_ & ~_04121_;
	assign _04142_ = _04099_ & ~_04131_;
	assign _04153_ = ~_04142_;
	assign _04164_ = ~\mchip.design.inputMovesSync [3];
	assign _04175_ = _03557_ & ~_03600_;
	assign _04185_ = _04175_ & _03664_;
	assign _04196_ = _04185_ ^ _03481_;
	assign _04207_ = ~(_04175_ ^ _03664_);
	assign _04218_ = _04207_ | _03611_;
	assign _04228_ = ~(_04218_ | _04196_);
	assign _04239_ = \mchip.design.pve.fsm.currState [2] & ~_04228_;
	assign _04250_ = (\mchip.design.inputSwitchPVPSync  ? _04164_ : _04239_);
	assign _04261_ = _03600_ | _03557_;
	assign _04272_ = _04261_ | _04207_;
	assign _04282_ = _04272_ | _04196_;
	assign _04293_ = \mchip.design.pve.fsm.currState [2] & ~_04282_;
	assign _04304_ = (\mchip.design.inputSwitchPVPSync  ? \mchip.design.inputMovesSync [2] : _04293_);
	assign _04315_ = _04304_ | ~_04250_;
	assign _04325_ = ~(_03600_ & _03557_);
	assign _04336_ = _04325_ | _04207_;
	assign _04347_ = _04336_ | _04196_;
	assign _04358_ = \mchip.design.pve.fsm.currState [2] & ~_04347_;
	assign _04369_ = (\mchip.design.inputSwitchPVPSync  ? \mchip.design.inputMovesSync [1] : _04358_);
	assign _04379_ = ~(_04325_ & _04261_);
	assign _04390_ = _03481_ | ~_03664_;
	assign _04401_ = _04175_ & ~_04390_;
	assign _04412_ = _03600_ | ~_04401_;
	assign _04422_ = _04412_ | _04379_;
	assign _04433_ = _04422_ | ~_04207_;
	assign _04444_ = _04433_ | ~_04196_;
	assign _04455_ = ~(_04444_ & \mchip.design.pve.fsm.currState [2]);
	assign _04466_ = (\mchip.design.inputSwitchPVPSync  ? \mchip.design.inputMovesSync [0] : _04455_);
	assign _04476_ = _04466_ | _04369_;
	assign _04487_ = ~(_04476_ | _04315_);
	assign _04498_ = _04261_ | ~_04207_;
	assign _04508_ = _04498_ | _04196_;
	assign _04519_ = \mchip.design.pve.fsm.currState [2] & ~_04508_;
	assign _04530_ = (\mchip.design.inputSwitchPVPSync  ? \mchip.design.inputMovesSync [6] : _04519_);
	assign _04541_ = _04325_ | ~_04207_;
	assign _04552_ = _04541_ | _04196_;
	assign _04563_ = \mchip.design.pve.fsm.currState [2] & ~_04552_;
	assign _04573_ = (\mchip.design.inputSwitchPVPSync  ? \mchip.design.inputMovesSync [5] : _04563_);
	assign _04584_ = _04401_ | _03600_;
	assign _04595_ = _04584_ | _04379_;
	assign _04605_ = _04595_ | _04207_;
	assign _04616_ = _04605_ | _04196_;
	assign _04627_ = \mchip.design.pve.fsm.currState [2] & ~_04616_;
	assign _04638_ = (\mchip.design.inputSwitchPVPSync  ? \mchip.design.inputMovesSync [4] : _04627_);
	assign _04649_ = _04638_ | ~_04573_;
	assign _04659_ = _04649_ | _04530_;
	assign _04670_ = _04487_ & ~_04659_;
	assign _04681_ = _04638_ | _04573_;
	assign _04692_ = _04681_ | ~_04530_;
	assign _04702_ = _04487_ & ~_04692_;
	assign _04713_ = _04702_ | _04670_;
	assign _04724_ = _04573_ | ~_04638_;
	assign _04735_ = _04724_ | _04530_;
	assign _04746_ = _04487_ & ~_04735_;
	assign _04756_ = _04746_ | _04713_;
	assign _04767_ = (\mchip.design.owner.fsm.currState  ? _04756_ : _04153_);
	assign _04778_ = _04056_ & ~_04067_;
	assign _04789_ = \mchip.design.inputMovesSync [2] | ~\mchip.design.inputMovesSync [3];
	assign _04799_ = _04789_ | _03992_;
	assign _04810_ = _04778_ & ~_04799_;
	assign _04821_ = _04810_ | _04131_;
	assign _04832_ = _04099_ & ~_04821_;
	assign _04843_ = \mchip.design.inputMovesSync [1] | ~\mchip.design.inputMovesSync [0];
	assign _04853_ = _04843_ | _04002_;
	assign _04864_ = _04778_ & ~_04853_;
	assign _04875_ = \mchip.design.inputMovesSync [0] | ~\mchip.design.inputMovesSync [1];
	assign _04886_ = _04875_ | _04002_;
	assign _04896_ = _04778_ & ~_04886_;
	assign _04907_ = \mchip.design.inputMovesSync [3] | ~\mchip.design.inputMovesSync [2];
	assign _04918_ = _04907_ | _03992_;
	assign _04929_ = _04778_ & ~_04918_;
	assign _04940_ = _04929_ | _04896_;
	assign _04950_ = _04940_ | _04864_;
	assign _04961_ = _04832_ & ~_04950_;
	assign _04972_ = ~(_04681_ | _04530_);
	assign _04982_ = _04369_ | ~_04466_;
	assign _04993_ = _04982_ | _04315_;
	assign _05004_ = _04993_ | ~_04972_;
	assign _05015_ = ~(_04304_ & _04250_);
	assign _05025_ = _05015_ | _04476_;
	assign _05036_ = _05025_ | ~_04972_;
	assign _05047_ = _04466_ | ~_04369_;
	assign _05057_ = _05047_ | _04315_;
	assign _05068_ = _04972_ & ~_05057_;
	assign _05079_ = _05068_ | ~_05036_;
	assign _05090_ = _05004_ & ~_05079_;
	assign _05100_ = _04304_ | _04250_;
	assign _05111_ = _05100_ | _04476_;
	assign _05122_ = _04972_ & ~_05111_;
	assign _05132_ = _05122_ | _04746_;
	assign _05143_ = _05132_ | _04713_;
	assign _05154_ = _05090_ & ~_05143_;
	assign _05165_ = (\mchip.design.owner.fsm.currState  ? _05154_ : _04961_);
	assign _01343_ = _05165_ | _04767_;
	assign _05185_ = _04810_ | _04045_;
	assign _05196_ = _05185_ | _04896_;
	assign _05206_ = ~(_05196_ | _04961_);
	assign _05217_ = _05143_ | ~_05090_;
	assign _05228_ = _05122_ | _04670_;
	assign _05239_ = _05228_ | _05068_;
	assign _05249_ = _05217_ & ~_05239_;
	assign _05260_ = (\mchip.design.owner.fsm.currState  ? _05249_ : _05206_);
	assign _05271_ = _04810_ | _04089_;
	assign _05281_ = _05271_ | _04929_;
	assign _05292_ = _05281_ & ~_04961_;
	assign _05303_ = _05122_ | _04702_;
	assign _05314_ = _05036_ & ~_05303_;
	assign _05324_ = _05217_ & ~_05314_;
	assign _05335_ = (\mchip.design.owner.fsm.currState  ? _05324_ : _05292_);
	assign _05346_ = _05260_ | ~_05335_;
	assign _05356_ = _05165_ | ~_04767_;
	assign _05367_ = _05346_ & ~_05356_;
	assign _05378_ = _01343_ & ~_05367_;
	assign _05389_ = ~\mchip.design.owner.tokens [28];
	assign _05399_ = ~\mchip.design.owner.tokens [30];
	assign _05410_ = (_05260_ ? _05389_ : _05399_);
	assign _05421_ = _05335_ | _05260_;
	assign _05431_ = ~(_05335_ & _05260_);
	assign _05442_ = _05431_ & _05421_;
	assign _05453_ = ~\mchip.design.owner.tokens [24];
	assign _05464_ = ~\mchip.design.owner.tokens [26];
	assign _05474_ = (_05260_ ? _05453_ : _05464_);
	assign _05485_ = (_05442_ ? _05410_ : _05474_);
	assign _01309_ = _05346_ ^ _04767_;
	assign _05505_ = ~\mchip.design.owner.tokens [20];
	assign _05516_ = ~\mchip.design.owner.tokens [22];
	assign _05527_ = (_05260_ ? _05505_ : _05516_);
	assign _05538_ = ~\mchip.design.owner.tokens [16];
	assign _05548_ = ~\mchip.design.owner.tokens [18];
	assign _05559_ = (_05260_ ? _05538_ : _05548_);
	assign _05570_ = (_05442_ ? _05527_ : _05559_);
	assign _05580_ = (_01309_ ? _05485_ : _05570_);
	assign _05591_ = _04767_ & ~_05346_;
	assign _05602_ = _05591_ ^ _05165_;
	assign _05613_ = ~\mchip.design.owner.tokens [12];
	assign _05623_ = ~\mchip.design.owner.tokens [14];
	assign _05634_ = (_05260_ ? _05613_ : _05623_);
	assign _05645_ = ~\mchip.design.owner.tokens [8];
	assign _05654_ = ~\mchip.design.owner.tokens [10];
	assign _05665_ = (_05260_ ? _05645_ : _05654_);
	assign _05675_ = (_05442_ ? _05634_ : _05665_);
	assign _05684_ = ~\mchip.design.owner.tokens [4];
	assign _05691_ = ~\mchip.design.owner.tokens [6];
	assign _05698_ = (_05260_ ? _05684_ : _05691_);
	assign _05705_ = ~\mchip.design.owner.tokens [0];
	assign _05712_ = ~\mchip.design.owner.tokens [2];
	assign _05719_ = (_05260_ ? _05705_ : _05712_);
	assign _05724_ = (_05442_ ? _05698_ : _05719_);
	assign _05728_ = (_01309_ ? _05675_ : _05724_);
	assign _05734_ = (_05602_ ? _05580_ : _05728_);
	assign _05742_ = ~\mchip.design.owner.tokens [82];
	assign _05748_ = ~\mchip.design.owner.tokens [80];
	assign _05756_ = (_05260_ ? _05748_ : _05742_);
	assign _05763_ = ~\mchip.design.owner.tokens [78];
	assign _05764_ = ~\mchip.design.owner.tokens [76];
	assign _05765_ = (_05260_ ? _05764_ : _05763_);
	assign _05766_ = ~\mchip.design.owner.tokens [72];
	assign _05767_ = ~\mchip.design.owner.tokens [74];
	assign _05768_ = (_05260_ ? _05766_ : _05767_);
	assign _05769_ = (_05442_ ? _05765_ : _05768_);
	assign _05770_ = ~\mchip.design.owner.tokens [70];
	assign _05771_ = ~\mchip.design.owner.tokens [68];
	assign _05772_ = (_05260_ ? _05771_ : _05770_);
	assign _05773_ = ~\mchip.design.owner.tokens [64];
	assign _05774_ = ~\mchip.design.owner.tokens [66];
	assign _05775_ = (_05260_ ? _05773_ : _05774_);
	assign _05776_ = (_05442_ ? _05772_ : _05775_);
	assign _05777_ = ~(_05734_ | _05378_);
	assign _05778_ = ~\mchip.design.owner.tokens [29];
	assign _05779_ = ~\mchip.design.owner.tokens [31];
	assign _05780_ = (_05260_ ? _05778_ : _05779_);
	assign _05781_ = ~\mchip.design.owner.tokens [25];
	assign _05782_ = ~\mchip.design.owner.tokens [27];
	assign _05783_ = (_05260_ ? _05781_ : _05782_);
	assign _05784_ = (_05442_ ? _05780_ : _05783_);
	assign _05785_ = ~\mchip.design.owner.tokens [21];
	assign _05786_ = ~\mchip.design.owner.tokens [23];
	assign _05787_ = (_05260_ ? _05785_ : _05786_);
	assign _05788_ = ~\mchip.design.owner.tokens [17];
	assign _05789_ = ~\mchip.design.owner.tokens [19];
	assign _05790_ = (_05260_ ? _05788_ : _05789_);
	assign _05791_ = (_05442_ ? _05787_ : _05790_);
	assign _05792_ = (_01309_ ? _05784_ : _05791_);
	assign _05793_ = ~\mchip.design.owner.tokens [13];
	assign _05794_ = ~\mchip.design.owner.tokens [15];
	assign _05795_ = (_05260_ ? _05793_ : _05794_);
	assign _05796_ = ~\mchip.design.owner.tokens [9];
	assign _05797_ = ~\mchip.design.owner.tokens [11];
	assign _05798_ = (_05260_ ? _05796_ : _05797_);
	assign _05799_ = (_05442_ ? _05795_ : _05798_);
	assign _05800_ = ~\mchip.design.owner.tokens [5];
	assign _05801_ = ~\mchip.design.owner.tokens [7];
	assign _05802_ = (_05260_ ? _05800_ : _05801_);
	assign _05803_ = ~\mchip.design.owner.tokens [1];
	assign _05804_ = ~\mchip.design.owner.tokens [3];
	assign _05805_ = (_05260_ ? _05803_ : _05804_);
	assign _05806_ = (_05442_ ? _05802_ : _05805_);
	assign _05807_ = (_01309_ ? _05799_ : _05806_);
	assign _05808_ = (_05602_ ? _05792_ : _05807_);
	assign _05809_ = ~\mchip.design.owner.tokens [83];
	assign _05810_ = ~\mchip.design.owner.tokens [81];
	assign _05811_ = (_05260_ ? _05810_ : _05809_);
	assign _05812_ = ~\mchip.design.owner.tokens [79];
	assign _05813_ = ~\mchip.design.owner.tokens [77];
	assign _05814_ = (_05260_ ? _05813_ : _05812_);
	assign _05815_ = ~\mchip.design.owner.tokens [73];
	assign _05816_ = ~\mchip.design.owner.tokens [75];
	assign _05817_ = (_05260_ ? _05815_ : _05816_);
	assign _05818_ = (_05442_ ? _05814_ : _05817_);
	assign _05819_ = ~\mchip.design.owner.tokens [71];
	assign _05820_ = ~\mchip.design.owner.tokens [69];
	assign _05821_ = (_05260_ ? _05820_ : _05819_);
	assign _05822_ = ~\mchip.design.owner.tokens [65];
	assign _05823_ = ~\mchip.design.owner.tokens [67];
	assign _05824_ = (_05260_ ? _05822_ : _05823_);
	assign _05825_ = (_05442_ ? _05821_ : _05824_);
	assign _05826_ = ~(_05808_ | _05378_);
	assign _05827_ = _05826_ | _05777_;
	assign _05828_ = _01309_ | ~_05602_;
	assign _05829_ = _05828_ | ~_05431_;
	assign _05830_ = ~(_05602_ & _01309_);
	assign _05831_ = ~(_05830_ & _05829_);
	assign _05832_ = _05378_ & ~_05831_;
	assign _05833_ = ~\mchip.design.owner.tokens [60];
	assign _05834_ = ~\mchip.design.owner.tokens [62];
	assign _05835_ = (_05260_ ? _05834_ : _05833_);
	assign _05836_ = ~(_05431_ & _05346_);
	assign _05837_ = ~\mchip.design.owner.tokens [56];
	assign _05838_ = ~\mchip.design.owner.tokens [58];
	assign _05839_ = (_05260_ ? _05838_ : _05837_);
	assign _05840_ = (_05836_ ? _05835_ : _05839_);
	assign _05841_ = ~(_01309_ ^ _05431_);
	assign _05842_ = ~\mchip.design.owner.tokens [52];
	assign _05843_ = ~\mchip.design.owner.tokens [54];
	assign _05844_ = (_05260_ ? _05843_ : _05842_);
	assign _05845_ = ~\mchip.design.owner.tokens [48];
	assign _05846_ = ~\mchip.design.owner.tokens [50];
	assign _05847_ = (_05260_ ? _05846_ : _05845_);
	assign _05848_ = (_05836_ ? _05844_ : _05847_);
	assign _05849_ = (_05841_ ? _05840_ : _05848_);
	assign _05850_ = ~(_01309_ | _05431_);
	assign _05851_ = ~(_05850_ ^ _05602_);
	assign _05852_ = ~\mchip.design.owner.tokens [44];
	assign _05853_ = ~\mchip.design.owner.tokens [46];
	assign _05854_ = (_05260_ ? _05853_ : _05852_);
	assign _05855_ = ~\mchip.design.owner.tokens [40];
	assign _05856_ = ~\mchip.design.owner.tokens [42];
	assign _05857_ = (_05260_ ? _05856_ : _05855_);
	assign _05858_ = (_05836_ ? _05854_ : _05857_);
	assign _05859_ = ~\mchip.design.owner.tokens [36];
	assign _05860_ = ~\mchip.design.owner.tokens [38];
	assign _05861_ = (_05260_ ? _05860_ : _05859_);
	assign _05862_ = ~\mchip.design.owner.tokens [32];
	assign _05863_ = ~\mchip.design.owner.tokens [34];
	assign _05864_ = (_05260_ ? _05863_ : _05862_);
	assign _05865_ = (_05836_ ? _05861_ : _05864_);
	assign _05866_ = (_05841_ ? _05858_ : _05865_);
	assign _05867_ = (_05851_ ? _05849_ : _05866_);
	assign _05868_ = _05831_ ^ _05378_;
	assign _05869_ = (_05260_ ? _05399_ : _05389_);
	assign _05870_ = (_05260_ ? _05464_ : _05453_);
	assign _05871_ = (_05836_ ? _05869_ : _05870_);
	assign _05872_ = (_05260_ ? _05516_ : _05505_);
	assign _05873_ = (_05260_ ? _05548_ : _05538_);
	assign _05874_ = (_05836_ ? _05872_ : _05873_);
	assign _05875_ = (_05841_ ? _05871_ : _05874_);
	assign _05876_ = (_05260_ ? _05623_ : _05613_);
	assign _05877_ = (_05260_ ? _05654_ : _05645_);
	assign _05878_ = (_05836_ ? _05876_ : _05877_);
	assign _05879_ = (_05260_ ? _05691_ : _05684_);
	assign _05880_ = (_05260_ ? _05712_ : _05705_);
	assign _05881_ = (_05836_ ? _05879_ : _05880_);
	assign _05882_ = (_05841_ ? _05878_ : _05881_);
	assign _05883_ = (_05851_ ? _05875_ : _05882_);
	assign _05884_ = (_05868_ ? _05867_ : _05883_);
	assign _05885_ = ~(_05884_ | _05832_);
	assign _05886_ = ~\mchip.design.owner.tokens [61];
	assign _05887_ = ~\mchip.design.owner.tokens [63];
	assign _05888_ = (_05260_ ? _05887_ : _05886_);
	assign _05889_ = ~\mchip.design.owner.tokens [57];
	assign _05890_ = ~\mchip.design.owner.tokens [59];
	assign _05891_ = (_05260_ ? _05890_ : _05889_);
	assign _05892_ = (_05836_ ? _05888_ : _05891_);
	assign _05893_ = ~\mchip.design.owner.tokens [53];
	assign _05894_ = ~\mchip.design.owner.tokens [55];
	assign _05895_ = (_05260_ ? _05894_ : _05893_);
	assign _05896_ = ~\mchip.design.owner.tokens [49];
	assign _05897_ = ~\mchip.design.owner.tokens [51];
	assign _05898_ = (_05260_ ? _05897_ : _05896_);
	assign _05899_ = (_05836_ ? _05895_ : _05898_);
	assign _05900_ = (_05841_ ? _05892_ : _05899_);
	assign _05901_ = ~\mchip.design.owner.tokens [45];
	assign _05902_ = ~\mchip.design.owner.tokens [47];
	assign _05903_ = (_05260_ ? _05902_ : _05901_);
	assign _05904_ = ~\mchip.design.owner.tokens [41];
	assign _05905_ = ~\mchip.design.owner.tokens [43];
	assign _05906_ = (_05260_ ? _05905_ : _05904_);
	assign _05907_ = (_05836_ ? _05903_ : _05906_);
	assign _05908_ = ~\mchip.design.owner.tokens [37];
	assign _05909_ = ~\mchip.design.owner.tokens [39];
	assign _05910_ = (_05260_ ? _05909_ : _05908_);
	assign _05911_ = ~\mchip.design.owner.tokens [33];
	assign _05912_ = ~\mchip.design.owner.tokens [35];
	assign _05913_ = (_05260_ ? _05912_ : _05911_);
	assign _05914_ = (_05836_ ? _05910_ : _05913_);
	assign _05915_ = (_05841_ ? _05907_ : _05914_);
	assign _05916_ = (_05851_ ? _05900_ : _05915_);
	assign _05917_ = (_05260_ ? _05779_ : _05778_);
	assign _05918_ = (_05260_ ? _05782_ : _05781_);
	assign _05919_ = (_05836_ ? _05917_ : _05918_);
	assign _05920_ = (_05260_ ? _05786_ : _05785_);
	assign _05921_ = (_05260_ ? _05789_ : _05788_);
	assign _05922_ = (_05836_ ? _05920_ : _05921_);
	assign _05923_ = (_05841_ ? _05919_ : _05922_);
	assign _05924_ = (_05260_ ? _05794_ : _05793_);
	assign _05925_ = (_05260_ ? _05797_ : _05796_);
	assign _05926_ = (_05836_ ? _05924_ : _05925_);
	assign _05927_ = (_05260_ ? _05801_ : _05800_);
	assign _05928_ = (_05260_ ? _05804_ : _05803_);
	assign _05929_ = (_05836_ ? _05927_ : _05928_);
	assign _05930_ = (_05841_ ? _05926_ : _05929_);
	assign _05931_ = (_05851_ ? _05923_ : _05930_);
	assign _05932_ = (_05868_ ? _05916_ : _05931_);
	assign _05933_ = ~(_05932_ | _05832_);
	assign _05934_ = _05933_ | _05885_;
	assign _05935_ = ~(_05934_ & _05827_);
	assign _05936_ = ~(_05602_ & _05378_);
	assign _05937_ = _05378_ & ~_05602_;
	assign _05938_ = ~(_01309_ | _05442_);
	assign _05939_ = _05937_ & ~_05938_;
	assign _05940_ = _05936_ & ~_05939_;
	assign _05941_ = _05940_ & _05378_;
	assign _05942_ = _05811_ | ~_05442_;
	assign _05943_ = _01309_ | ~_05442_;
	assign _05944_ = _05442_ | ~_01309_;
	assign _05945_ = _05944_ & _05943_;
	assign _05946_ = _05945_ | _05942_;
	assign _05947_ = _05938_ ^ _05602_;
	assign _05948_ = (_05442_ ? _05817_ : _05814_);
	assign _05949_ = (_05442_ ? _05824_ : _05821_);
	assign _05950_ = (_05945_ ? _05948_ : _05949_);
	assign _05951_ = (_05947_ ? _05946_ : _05950_);
	assign _05952_ = _05938_ & ~_05602_;
	assign _05953_ = ~(_05952_ ^ _05378_);
	assign _05954_ = _05953_ | _05951_;
	assign _05955_ = ~(_05940_ ^ _05378_);
	assign _05956_ = (_05442_ ? _05783_ : _05780_);
	assign _05957_ = (_05442_ ? _05790_ : _05787_);
	assign _05958_ = (_05945_ ? _05956_ : _05957_);
	assign _05959_ = (_05442_ ? _05798_ : _05795_);
	assign _05960_ = (_05442_ ? _05805_ : _05802_);
	assign _05961_ = (_05945_ ? _05959_ : _05960_);
	assign _05962_ = (_05947_ ? _05958_ : _05961_);
	assign _05963_ = (_05260_ ? _05889_ : _05890_);
	assign _05964_ = (_05260_ ? _05886_ : _05887_);
	assign _05965_ = (_05442_ ? _05963_ : _05964_);
	assign _05966_ = (_05260_ ? _05896_ : _05897_);
	assign _05967_ = (_05260_ ? _05893_ : _05894_);
	assign _05968_ = (_05442_ ? _05966_ : _05967_);
	assign _05969_ = (_05945_ ? _05965_ : _05968_);
	assign _05970_ = (_05260_ ? _05904_ : _05905_);
	assign _05971_ = (_05260_ ? _05901_ : _05902_);
	assign _05972_ = (_05442_ ? _05970_ : _05971_);
	assign _05973_ = (_05260_ ? _05911_ : _05912_);
	assign _05974_ = (_05260_ ? _05908_ : _05909_);
	assign _05975_ = (_05442_ ? _05973_ : _05974_);
	assign _05976_ = (_05945_ ? _05972_ : _05975_);
	assign _05977_ = (_05947_ ? _05969_ : _05976_);
	assign _05978_ = (_05953_ ? _05977_ : _05962_);
	assign _05979_ = (_05955_ ? _05954_ : _05978_);
	assign _05980_ = ~(_05979_ | _05941_);
	assign _05981_ = _05756_ | ~_05442_;
	assign _05982_ = _05981_ | _05945_;
	assign _05983_ = (_05442_ ? _05768_ : _05765_);
	assign _05984_ = (_05442_ ? _05775_ : _05772_);
	assign _05985_ = (_05945_ ? _05983_ : _05984_);
	assign _05986_ = (_05947_ ? _05982_ : _05985_);
	assign _05987_ = _05986_ | _05953_;
	assign _05988_ = (_05442_ ? _05474_ : _05410_);
	assign _05989_ = (_05442_ ? _05559_ : _05527_);
	assign _05990_ = (_05945_ ? _05988_ : _05989_);
	assign _05991_ = (_05442_ ? _05665_ : _05634_);
	assign _05992_ = (_05442_ ? _05719_ : _05698_);
	assign _05993_ = (_05945_ ? _05991_ : _05992_);
	assign _05994_ = (_05947_ ? _05990_ : _05993_);
	assign _00146_ = (_05260_ ? _05837_ : _05838_);
	assign _00145_ = (_05260_ ? _05833_ : _05834_);
	assign _05995_ = (_05442_ ? _00146_ : _00145_);
	assign _00143_ = (_05260_ ? _05845_ : _05846_);
	assign _00142_ = (_05260_ ? _05842_ : _05843_);
	assign _05996_ = (_05442_ ? _00143_ : _00142_);
	assign _05997_ = (_05945_ ? _05995_ : _05996_);
	assign _00153_ = (_05260_ ? _05855_ : _05856_);
	assign _00152_ = (_05260_ ? _05852_ : _05853_);
	assign _05998_ = (_05442_ ? _00153_ : _00152_);
	assign _00150_ = (_05260_ ? _05862_ : _05863_);
	assign _00149_ = (_05260_ ? _05859_ : _05860_);
	assign _05999_ = (_05442_ ? _00150_ : _00149_);
	assign _06000_ = (_05945_ ? _05998_ : _05999_);
	assign _06001_ = (_05947_ ? _05997_ : _06000_);
	assign _06002_ = (_05953_ ? _06001_ : _05994_);
	assign _06003_ = (_05955_ ? _05987_ : _06002_);
	assign _06004_ = ~(_06003_ | _05941_);
	assign _06005_ = _06004_ | _05980_;
	assign _06006_ = ~(_05828_ | _05346_);
	assign _06007_ = _05830_ & ~_06006_;
	assign _06008_ = ~(_06007_ | _05378_);
	assign _06009_ = (_05260_ ? _05742_ : _05748_);
	assign _06010_ = ~(_05442_ ^ _05260_);
	assign _06011_ = _06010_ | _06009_;
	assign _06012_ = ~_05260_;
	assign _06013_ = _04767_ | _06011_;
	assign _01341_ = ~(_05165_ ^ _04767_);
	assign _06014_ = (_05260_ ? _05763_ : _05764_);
	assign _06015_ = (_05260_ ? _05767_ : _05766_);
	assign _06016_ = (_06010_ ? _06014_ : _06015_);
	assign _06017_ = (_05260_ ? _05770_ : _05771_);
	assign _06018_ = (_05260_ ? _05774_ : _05773_);
	assign _06019_ = (_06010_ ? _06017_ : _06018_);
	assign _06020_ = (_04767_ ? _06016_ : _06019_);
	assign _06021_ = (_01341_ ? _06013_ : _06020_);
	assign _06022_ = ~(_05165_ & _04767_);
	assign _06023_ = _06022_ | _06021_;
	assign _06024_ = (_06010_ ? _05835_ : _05839_);
	assign _06025_ = (_06010_ ? _05844_ : _05847_);
	assign _06026_ = (_04767_ ? _06024_ : _06025_);
	assign _06027_ = (_06010_ ? _05854_ : _05857_);
	assign _06028_ = (_06010_ ? _05861_ : _05864_);
	assign _06029_ = (_04767_ ? _06027_ : _06028_);
	assign _06030_ = (_01341_ ? _06026_ : _06029_);
	assign _06031_ = (_06010_ ? _05869_ : _05870_);
	assign _06032_ = (_06010_ ? _05872_ : _05873_);
	assign _06033_ = (_04767_ ? _06031_ : _06032_);
	assign _06034_ = (_06010_ ? _05876_ : _05877_);
	assign _06035_ = (_06010_ ? _05879_ : _05880_);
	assign _06036_ = (_04767_ ? _06034_ : _06035_);
	assign _06037_ = (_01341_ ? _06033_ : _06036_);
	assign _06038_ = (_06022_ ? _06030_ : _06037_);
	assign _06039_ = (_06008_ ? _06023_ : _06038_);
	assign _06040_ = (_05260_ ? _05809_ : _05810_);
	assign _06041_ = _06040_ | _06010_;
	assign _06042_ = _06041_ | _04767_;
	assign _06043_ = (_05260_ ? _05812_ : _05813_);
	assign _06044_ = (_05260_ ? _05816_ : _05815_);
	assign _06045_ = (_06010_ ? _06043_ : _06044_);
	assign _06046_ = (_05260_ ? _05819_ : _05820_);
	assign _06047_ = (_05260_ ? _05823_ : _05822_);
	assign _06048_ = (_06010_ ? _06046_ : _06047_);
	assign _06049_ = (_04767_ ? _06045_ : _06048_);
	assign _06050_ = (_01341_ ? _06042_ : _06049_);
	assign _06051_ = ~(_06050_ | _06022_);
	assign _06052_ = (_05260_ ? \mchip.design.owner.tokens [63] : \mchip.design.owner.tokens [61]);
	assign _06053_ = (_05260_ ? \mchip.design.owner.tokens [59] : \mchip.design.owner.tokens [57]);
	assign _06054_ = (_06010_ ? _06052_ : _06053_);
	assign _06055_ = (_05260_ ? \mchip.design.owner.tokens [55] : \mchip.design.owner.tokens [53]);
	assign _06056_ = (_05260_ ? \mchip.design.owner.tokens [51] : \mchip.design.owner.tokens [49]);
	assign _06057_ = (_06010_ ? _06055_ : _06056_);
	assign _06058_ = (_04767_ ? _06054_ : _06057_);
	assign _06059_ = (_05260_ ? \mchip.design.owner.tokens [47] : \mchip.design.owner.tokens [45]);
	assign _06060_ = (_05260_ ? \mchip.design.owner.tokens [43] : \mchip.design.owner.tokens [41]);
	assign _00108_ = (_06010_ ? _06059_ : _06060_);
	assign _00109_ = (_05260_ ? \mchip.design.owner.tokens [39] : \mchip.design.owner.tokens [37]);
	assign _00110_ = (_05260_ ? \mchip.design.owner.tokens [35] : \mchip.design.owner.tokens [33]);
	assign _00111_ = (_06010_ ? _00109_ : _00110_);
	assign _00112_ = (_04767_ ? _00108_ : _00111_);
	assign _00113_ = (_01341_ ? _06058_ : _00112_);
	assign _00114_ = (_05260_ ? \mchip.design.owner.tokens [31] : \mchip.design.owner.tokens [29]);
	assign _00115_ = (_05260_ ? \mchip.design.owner.tokens [27] : \mchip.design.owner.tokens [25]);
	assign _00116_ = (_06010_ ? _00114_ : _00115_);
	assign _00117_ = (_05260_ ? \mchip.design.owner.tokens [23] : \mchip.design.owner.tokens [21]);
	assign _00118_ = (_05260_ ? \mchip.design.owner.tokens [19] : \mchip.design.owner.tokens [17]);
	assign _00119_ = (_06010_ ? _00117_ : _00118_);
	assign _00120_ = (_04767_ ? _00116_ : _00119_);
	assign _00121_ = (_05260_ ? \mchip.design.owner.tokens [15] : \mchip.design.owner.tokens [13]);
	assign _00122_ = (_05260_ ? \mchip.design.owner.tokens [11] : \mchip.design.owner.tokens [9]);
	assign _00123_ = (_06010_ ? _00121_ : _00122_);
	assign _00124_ = (_05260_ ? \mchip.design.owner.tokens [7] : \mchip.design.owner.tokens [5]);
	assign _00125_ = (_05260_ ? \mchip.design.owner.tokens [3] : \mchip.design.owner.tokens [1]);
	assign _00126_ = (_06010_ ? _00124_ : _00125_);
	assign _00127_ = (_04767_ ? _00123_ : _00126_);
	assign _00128_ = (_01341_ ? _00120_ : _00127_);
	assign _00129_ = (_06022_ ? _00113_ : _00128_);
	assign _00130_ = (_06008_ ? _06051_ : _00129_);
	assign _00131_ = _00130_ | ~_06039_;
	assign _00132_ = ~(_00131_ & _06005_);
	assign _00133_ = ~(_05602_ | _01309_);
	assign _00134_ = ~(_00133_ | _05378_);
	assign _00135_ = _05756_ | _05442_;
	assign _00136_ = _00135_ | ~_01309_;
	assign _00137_ = ~(_05602_ ^ _01309_);
	assign _00138_ = (_01309_ ? _05776_ : _05769_);
	assign _00139_ = (_00137_ ? _00136_ : _00138_);
	assign _00140_ = _00133_ ^ _05378_;
	assign _00141_ = _00140_ | _00139_;
	assign _00144_ = (_05442_ ? _00142_ : _00143_);
	assign _00147_ = (_05442_ ? _00145_ : _00146_);
	assign _00148_ = (_01309_ ? _00144_ : _00147_);
	assign _00151_ = (_05442_ ? _00149_ : _00150_);
	assign _00154_ = (_05442_ ? _00152_ : _00153_);
	assign _00155_ = (_01309_ ? _00151_ : _00154_);
	assign _00156_ = (_00137_ ? _00148_ : _00155_);
	assign _00157_ = (_01309_ ? _05570_ : _05485_);
	assign _00158_ = (_01309_ ? _05724_ : _05675_);
	assign _00159_ = (_00137_ ? _00157_ : _00158_);
	assign _00160_ = (_00140_ ? _00156_ : _00159_);
	assign _00161_ = (_00134_ ? _00141_ : _00160_);
	assign _00162_ = _05811_ | _05442_;
	assign _00163_ = _00162_ | ~_01309_;
	assign _00164_ = (_01309_ ? _05825_ : _05818_);
	assign _00165_ = (_00137_ ? _00163_ : _00164_);
	assign _00166_ = ~(_00165_ | _00140_);
	assign _00167_ = ~_05966_;
	assign _00168_ = ~_05967_;
	assign _00169_ = (_05442_ ? _00168_ : _00167_);
	assign _00170_ = ~_05963_;
	assign _00171_ = ~_05964_;
	assign _00172_ = (_05442_ ? _00171_ : _00170_);
	assign _00173_ = (_01309_ ? _00169_ : _00172_);
	assign _00174_ = ~_05973_;
	assign _00175_ = ~_05974_;
	assign _00176_ = (_05442_ ? _00175_ : _00174_);
	assign _00177_ = ~_05970_;
	assign _00178_ = ~_05971_;
	assign _00179_ = (_05442_ ? _00178_ : _00177_);
	assign _00180_ = (_01309_ ? _00176_ : _00179_);
	assign _00181_ = (_00137_ ? _00173_ : _00180_);
	assign _00182_ = ~_05790_;
	assign _00183_ = ~_05787_;
	assign _00184_ = (_05442_ ? _00183_ : _00182_);
	assign _00185_ = ~_05783_;
	assign _00186_ = ~_05780_;
	assign _00187_ = (_05442_ ? _00186_ : _00185_);
	assign _00188_ = (_01309_ ? _00184_ : _00187_);
	assign _00189_ = ~_05805_;
	assign _00190_ = ~_05802_;
	assign _00191_ = (_05442_ ? _00190_ : _00189_);
	assign _00192_ = ~_05798_;
	assign _00193_ = ~_05795_;
	assign _00194_ = (_05442_ ? _00193_ : _00192_);
	assign _00195_ = (_01309_ ? _00191_ : _00194_);
	assign _00196_ = (_00137_ ? _00188_ : _00195_);
	assign _00197_ = (_00140_ ? _00181_ : _00196_);
	assign _00198_ = (_00134_ ? _00166_ : _00197_);
	assign _00199_ = _00198_ | ~_00161_;
	assign _00200_ = _06009_ | _05836_;
	assign _00201_ = _01309_ & _05431_;
	assign _00202_ = ~(_00201_ | _05850_);
	assign _00203_ = _00202_ | _00200_;
	assign _00204_ = _00201_ ^ _05602_;
	assign _00205_ = (_05836_ ? _06014_ : _06015_);
	assign _00206_ = (_05836_ ? _06017_ : _06018_);
	assign _00207_ = (_00202_ ? _00205_ : _00206_);
	assign _00208_ = (_00204_ ? _00203_ : _00207_);
	assign _00209_ = _05431_ & ~_05830_;
	assign _00210_ = _00209_ ^ _05378_;
	assign _00211_ = _00210_ | _00208_;
	assign _00212_ = _00209_ | ~_05378_;
	assign _00213_ = (_00202_ ? _05840_ : _05848_);
	assign _00214_ = (_00202_ ? _05858_ : _05865_);
	assign _00215_ = (_00204_ ? _00213_ : _00214_);
	assign _00216_ = (_00202_ ? _05871_ : _05874_);
	assign _00217_ = (_00202_ ? _05878_ : _05881_);
	assign _00218_ = (_00204_ ? _00216_ : _00217_);
	assign _00219_ = (_00210_ ? _00215_ : _00218_);
	assign _00220_ = (_00212_ ? _00211_ : _00219_);
	assign _00221_ = _06040_ | _05836_;
	assign _00222_ = _00221_ | _00202_;
	assign _00223_ = (_05836_ ? _06043_ : _06044_);
	assign _00224_ = (_05836_ ? _06046_ : _06047_);
	assign _00225_ = (_00202_ ? _00223_ : _00224_);
	assign _00226_ = (_00204_ ? _00222_ : _00225_);
	assign _00227_ = ~(_00226_ | _00210_);
	assign _00228_ = (_05836_ ? _06052_ : _06053_);
	assign _00229_ = (_05836_ ? _06055_ : _06056_);
	assign _00230_ = (_00202_ ? _00228_ : _00229_);
	assign _00231_ = (_05836_ ? _06059_ : _06060_);
	assign _00232_ = (_05836_ ? _00109_ : _00110_);
	assign _00233_ = (_00202_ ? _00231_ : _00232_);
	assign _00234_ = (_00204_ ? _00230_ : _00233_);
	assign _00235_ = (_05836_ ? _00114_ : _00115_);
	assign _00236_ = (_05836_ ? _00117_ : _00118_);
	assign _00237_ = (_00202_ ? _00235_ : _00236_);
	assign _00238_ = (_05836_ ? _00121_ : _00122_);
	assign _00239_ = (_05836_ ? _00124_ : _00125_);
	assign _00240_ = (_00202_ ? _00238_ : _00239_);
	assign _00241_ = (_00204_ ? _00237_ : _00240_);
	assign _00242_ = (_00210_ ? _00234_ : _00241_);
	assign _00243_ = (_00212_ ? _00227_ : _00242_);
	assign _00244_ = _00220_ & ~_00243_;
	assign _00245_ = _00244_ | ~_00199_;
	assign _00246_ = _00245_ | _00132_;
	assign _00247_ = ~(_00246_ | _05935_);
	assign _00248_ = (\mchip.design.inputSwitchPVPSync  ? \mchip.design.currStateConfirm [1] : \mchip.design.pve.fsm.currState [2]);
	assign _00249_ = (\mchip.design.owner.fsm.currState  ? _00248_ : \mchip.design.currStateConfirm [1]);
	assign _00006_ = _00249_ & ~_00247_;
	assign _00250_ = \mchip.design.debounceCount [20] & ~\mchip.design.debounceCount [21];
	assign _00251_ = ~(_00250_ & \mchip.design.debounceCount [22]);
	assign _00252_ = \mchip.design.debounceCount [16] & \mchip.design.debounceCount [17];
	assign _00253_ = \mchip.design.debounceCount [18] & \mchip.design.debounceCount [19];
	assign _00254_ = ~(_00253_ & _00252_);
	assign _00255_ = _00254_ | _00251_;
	assign _00256_ = \mchip.design.debounceCount [10] & \mchip.design.debounceCount [11];
	assign _00257_ = \mchip.design.debounceCount [8] | ~\mchip.design.debounceCount [9];
	assign _00258_ = _00256_ & ~_00257_;
	assign _00259_ = \mchip.design.debounceCount [13] | ~\mchip.design.debounceCount [12];
	assign _00260_ = \mchip.design.debounceCount [15] | ~\mchip.design.debounceCount [14];
	assign _00261_ = _00260_ | _00259_;
	assign _00262_ = _00261_ | ~_00258_;
	assign _00263_ = \mchip.design.debounceCount [4] & ~\mchip.design.debounceCount [5];
	assign _00264_ = ~(\mchip.design.debounceCount [6] | \mchip.design.debounceCount [7]);
	assign _00265_ = ~(_00264_ & _00263_);
	assign _00266_ = \mchip.design.debounceCount [2] | \mchip.design.debounceCount [3];
	assign _00267_ = \mchip.design.debounceCount [0] | \mchip.design.debounceCount [1];
	assign _00268_ = _00267_ | _00266_;
	assign _00269_ = _00268_ | _00265_;
	assign _00270_ = _00269_ | _00262_;
	assign _00271_ = _00270_ | _00255_;
	assign _00272_ = _00260_ | ~\mchip.design.debounceCount [13];
	assign _00273_ = _00272_ & ~\mchip.design.debounceCount [15];
	assign _00274_ = _00273_ | _00254_;
	assign _00275_ = ~(_00261_ | _00254_);
	assign _00276_ = ~(\mchip.design.debounceCount [9] & \mchip.design.debounceCount [8]);
	assign _00277_ = _00276_ | ~_00256_;
	assign _00278_ = \mchip.design.debounceCount [5] | \mchip.design.debounceCount [4];
	assign _00279_ = _00264_ & ~_00278_;
	assign _00280_ = _00258_ & ~_00279_;
	assign _00281_ = _00277_ & ~_00280_;
	assign _00282_ = _00275_ & ~_00281_;
	assign _00283_ = _00274_ & ~_00282_;
	assign _00284_ = _00283_ | ~_00250_;
	assign _00285_ = _00284_ & ~\mchip.design.debounceCount [21];
	assign _00286_ = \mchip.design.debounceCount [22] & ~_00285_;
	assign _00287_ = _00271_ & ~_00286_;
	assign _00288_ = ~(_00287_ | \mchip.design.inputConfirmSync );
	assign _00289_ = _00288_ | io_in[13];
	assign _00290_ = \mchip.design.currStateConfirm [2] & ~_00289_;
	assign _00291_ = \mchip.design.currStateConfirm [1] & ~io_in[13];
	assign _00003_ = _00291_ | _00290_;
	assign _06062_[0] = ~\mchip.design.debounceCount [0];
	assign _00292_ = \mchip.design.inputConfirmSync  | io_in[13];
	assign _00293_ = \mchip.design.currStateConfirm [0] & ~_00292_;
	assign _00294_ = io_in[13] | ~_00288_;
	assign _00295_ = \mchip.design.currStateConfirm [2] & ~_00294_;
	assign _00296_ = _00295_ | io_in[13];
	assign _00002_ = _00296_ | _00293_;
	assign _00297_ = \mchip.design.vga.v_idx [8] & ~\mchip.design.vga.v_idx [9];
	assign _00298_ = \mchip.design.vga.v_idx [0] | \mchip.design.vga.v_idx [1];
	assign _00299_ = \mchip.design.vga.v_idx [2] | \mchip.design.vga.v_idx [3];
	assign _00300_ = _00299_ | _00298_;
	assign _00301_ = \mchip.design.vga.v_idx [6] & \mchip.design.vga.v_idx [7];
	assign _00302_ = \mchip.design.vga.v_idx [5] & ~\mchip.design.vga.v_idx [4];
	assign _00303_ = ~(_00302_ & _00301_);
	assign _00304_ = _00303_ | _00300_;
	assign _00305_ = ~(_00301_ & \mchip.design.vga.v_idx [5]);
	assign _00306_ = _00304_ & ~_00305_;
	assign _00307_ = _00297_ & ~_00306_;
	assign _00308_ = ~(\mchip.design.vga.v_idx [8] | \mchip.design.vga.v_idx [9]);
	assign _00309_ = _00308_ | _00307_;
	assign _00310_ = _00297_ & ~_00304_;
	assign _00311_ = _00309_ & ~_00310_;
	assign _00312_ = ~(\mchip.design.vga.h_idx [8] | \mchip.design.vga.h_idx [7]);
	assign _00313_ = \mchip.design.vga.h_idx [9] & ~_00312_;
	assign \mchip.design.blank  = _00311_ & ~_00313_;
	assign _00314_ = \mchip.design.vga.v_idx [1] | ~\mchip.design.vga.v_idx [0];
	assign _00315_ = \mchip.design.vga.v_idx [2] & \mchip.design.vga.v_idx [3];
	assign _00316_ = _00314_ | ~_00315_;
	assign _00317_ = \mchip.design.vga.v_idx [4] | \mchip.design.vga.v_idx [5];
	assign _00318_ = \mchip.design.vga.v_idx [6] | \mchip.design.vga.v_idx [7];
	assign _00319_ = _00318_ | _00317_;
	assign _00320_ = ~(_00319_ | _00316_);
	assign _00321_ = \mchip.design.vga.v_idx [9] & ~\mchip.design.vga.v_idx [8];
	assign _00322_ = ~(_00321_ & _00320_);
	assign _00323_ = ~(_00318_ | _00317_);
	assign _00324_ = _00315_ & _00298_;
	assign _00325_ = _00324_ & ~_00319_;
	assign _00326_ = _00323_ & ~_00325_;
	assign _00327_ = _00321_ & ~_00326_;
	assign _00328_ = \mchip.design.vga.v_idx [8] & \mchip.design.vga.v_idx [9];
	assign _00329_ = _00328_ | _00327_;
	assign _00330_ = _00322_ & ~_00329_;
	assign _00097_ = _00330_ & ~\mchip.design.vga.v_idx [0];
	assign _00331_ = \mchip.design.vga.v_idx [0] | ~\mchip.design.vga.v_idx [1];
	assign _00332_ = _00331_ & _00314_;
	assign _00098_ = _00330_ & ~_00332_;
	assign _00333_ = ~(\mchip.design.vga.v_idx [0] & \mchip.design.vga.v_idx [1]);
	assign _00334_ = _00333_ ^ \mchip.design.vga.v_idx [2];
	assign _00099_ = _00330_ & ~_00334_;
	assign _00335_ = ~\mchip.design.vga.v_idx [3];
	assign _00336_ = \mchip.design.vga.v_idx [2] & ~_00333_;
	assign _00337_ = _00336_ ^ _00335_;
	assign _00100_ = _00330_ & ~_00337_;
	assign _00338_ = ~\mchip.design.vga.v_idx [4];
	assign _00339_ = _00315_ & ~_00333_;
	assign _00340_ = _00339_ ^ _00338_;
	assign _00101_ = _00330_ & ~_00340_;
	assign _00341_ = ~\mchip.design.vga.v_idx [5];
	assign _00342_ = _00339_ & ~_00338_;
	assign _00343_ = _00342_ ^ _00341_;
	assign _00102_ = _00330_ & ~_00343_;
	assign _00344_ = ~\mchip.design.vga.v_idx [6];
	assign _00345_ = \mchip.design.vga.v_idx [4] & \mchip.design.vga.v_idx [5];
	assign _00346_ = ~_00345_;
	assign _00347_ = _00339_ & ~_00346_;
	assign _00348_ = _00347_ ^ _00344_;
	assign _00103_ = _00330_ & ~_00348_;
	assign _00349_ = ~\mchip.design.vga.v_idx [7];
	assign _00350_ = _00347_ & ~_00344_;
	assign _00351_ = _00350_ ^ _00349_;
	assign _00104_ = _00330_ & ~_00351_;
	assign _00352_ = ~\mchip.design.vga.v_idx [8];
	assign _00353_ = _00345_ & _00301_;
	assign _00354_ = _00353_ & _00339_;
	assign _00355_ = _00354_ & ~_00352_;
	assign _00356_ = _00352_ & ~_00354_;
	assign _00357_ = _00356_ | _00355_;
	assign _00105_ = _00330_ & ~_00357_;
	assign _00358_ = ~(_00355_ ^ \mchip.design.vga.v_idx [9]);
	assign _00106_ = _00330_ & ~_00358_;
	assign _00359_ = \mchip.design.vga.v_idx [5] | \mchip.design.vga.v_idx [6];
	assign _00360_ = ~(\mchip.design.vga.v_idx [7] | \mchip.design.vga.v_idx [8]);
	assign _00361_ = _00360_ & ~_00359_;
	assign _00362_ = \mchip.design.vga.v_idx [3] & \mchip.design.vga.v_idx [4];
	assign _00363_ = ~(\mchip.design.vga.v_idx [1] & \mchip.design.vga.v_idx [2]);
	assign _00364_ = _00362_ & ~_00363_;
	assign _00365_ = _00361_ & ~_00364_;
	assign _00366_ = \mchip.design.vga.v_idx [5] | ~\mchip.design.vga.v_idx [4];
	assign _00367_ = _00366_ | _00318_;
	assign _00368_ = _00367_ | _00316_;
	assign _00369_ = _00352_ & ~_00368_;
	assign _00370_ = ~(_00369_ | _00365_);
	assign _00371_ = ~(_00317_ | _00315_);
	assign _00372_ = \mchip.design.vga.v_idx [7] | ~\mchip.design.vga.v_idx [6];
	assign _00373_ = _00371_ & ~_00372_;
	assign _00374_ = _00318_ & ~_00373_;
	assign _00375_ = _00374_ | \mchip.design.vga.v_idx [8];
	assign _00376_ = ~(_00372_ | _00317_);
	assign _00377_ = \mchip.design.vga.v_idx [2] | ~\mchip.design.vga.v_idx [3];
	assign _00378_ = ~(_00377_ | _00333_);
	assign _00379_ = ~(_00378_ & _00376_);
	assign _00380_ = _00352_ & ~_00379_;
	assign _00381_ = _00380_ | _00375_;
	assign _00382_ = _00372_ | ~_00302_;
	assign _00383_ = ~(_00377_ | _00298_);
	assign _00384_ = _00382_ | ~_00383_;
	assign _00385_ = _00384_ | \mchip.design.vga.v_idx [8];
	assign _00386_ = _00341_ & ~_00372_;
	assign _00387_ = _00318_ & ~_00386_;
	assign _00388_ = _00383_ | _00335_;
	assign _00389_ = _00388_ & ~_00382_;
	assign _00390_ = _00387_ & ~_00389_;
	assign _00391_ = _00352_ & ~_00390_;
	assign _00392_ = _00385_ & ~_00391_;
	assign _00393_ = _00381_ & ~_00392_;
	assign _00394_ = _00370_ & ~_00393_;
	assign _00395_ = \mchip.design.vga.v_idx [6] | ~\mchip.design.vga.v_idx [7];
	assign _00396_ = ~(_00395_ | _00317_);
	assign _00397_ = \mchip.design.vga.v_idx [7] & ~_00396_;
	assign _00398_ = ~(_00395_ | _00366_);
	assign _00399_ = \mchip.design.vga.v_idx [3] | ~\mchip.design.vga.v_idx [2];
	assign _00400_ = _00333_ & ~_00399_;
	assign _00401_ = _00299_ & ~_00400_;
	assign _00402_ = _00398_ & ~_00401_;
	assign _00403_ = _00397_ & ~_00402_;
	assign _00404_ = _00403_ | \mchip.design.vga.v_idx [8];
	assign _00405_ = _00399_ | _00331_;
	assign _00406_ = _00405_ | ~_00398_;
	assign _00407_ = _00352_ & ~_00406_;
	assign _00408_ = _00407_ | _00404_;
	assign _00409_ = _00395_ | ~_00345_;
	assign _00410_ = _00333_ | _00299_;
	assign _00411_ = _00410_ | _00409_;
	assign _00412_ = _00411_ | \mchip.design.vga.v_idx [8];
	assign _00413_ = ~(_00345_ & _00299_);
	assign _00414_ = _00413_ & ~_00395_;
	assign _00415_ = \mchip.design.vga.v_idx [7] & ~_00414_;
	assign _00416_ = _00352_ & ~_00415_;
	assign _00417_ = _00412_ & ~_00416_;
	assign _00418_ = _00408_ & ~_00417_;
	assign _00419_ = _00394_ & ~_00418_;
	assign _00420_ = _00314_ | _00299_;
	assign _00421_ = _00420_ | _00303_;
	assign _00422_ = _00352_ & ~_00421_;
	assign _00423_ = ~_00360_;
	assign _00424_ = \mchip.design.vga.v_idx [5] & \mchip.design.vga.v_idx [6];
	assign _00425_ = \mchip.design.vga.v_idx [8] | ~\mchip.design.vga.v_idx [7];
	assign _00426_ = ~(_00425_ | _00424_);
	assign _00427_ = _00423_ & ~_00426_;
	assign _00428_ = _00424_ & ~_00425_;
	assign _00429_ = \mchip.design.vga.v_idx [3] | \mchip.design.vga.v_idx [4];
	assign _00430_ = ~(\mchip.design.vga.v_idx [1] | \mchip.design.vga.v_idx [2]);
	assign _00431_ = _00429_ | ~_00430_;
	assign _00432_ = _00428_ & ~_00431_;
	assign _00433_ = _00427_ & ~_00432_;
	assign _00434_ = _00433_ | _00422_;
	assign _00435_ = _00331_ | ~_00315_;
	assign _00436_ = _00435_ | ~_00353_;
	assign _00437_ = _00436_ | \mchip.design.vga.v_idx [8];
	assign _00438_ = _00353_ & ~_00339_;
	assign _00439_ = _00353_ & ~_00438_;
	assign _00440_ = _00352_ & ~_00439_;
	assign _00441_ = _00437_ & ~_00440_;
	assign _00442_ = _00434_ & ~_00441_;
	assign _00443_ = _00419_ & ~_00442_;
	assign _00444_ = _00315_ & _00302_;
	assign _00445_ = _00346_ & ~_00444_;
	assign _00446_ = _00445_ & ~_00318_;
	assign _00447_ = \mchip.design.vga.v_idx [8] & ~_00446_;
	assign _00448_ = _00302_ & ~_00318_;
	assign _00449_ = _00298_ | ~_00315_;
	assign _00450_ = _00449_ | ~_00448_;
	assign _00451_ = \mchip.design.vga.v_idx [8] & ~_00450_;
	assign _00452_ = _00451_ | _00447_;
	assign _00453_ = _00317_ & ~_00372_;
	assign _00454_ = _00349_ & ~_00453_;
	assign _00455_ = ~_00315_;
	assign _00456_ = _00298_ & ~_00377_;
	assign _00457_ = _00455_ & ~_00456_;
	assign _00458_ = _00376_ & ~_00457_;
	assign _00459_ = _00454_ & ~_00458_;
	assign _00460_ = \mchip.design.vga.v_idx [8] & ~_00459_;
	assign _00461_ = _00377_ | _00314_;
	assign _00462_ = _00461_ | ~_00376_;
	assign _00463_ = \mchip.design.vga.v_idx [8] & ~_00462_;
	assign _00464_ = _00460_ & ~_00463_;
	assign _00465_ = _00452_ & ~_00464_;
	assign _00466_ = _00443_ & ~_00465_;
	assign _00467_ = ~(_00399_ | _00333_);
	assign _00468_ = _00467_ | \mchip.design.vga.v_idx [3];
	assign _00469_ = _00372_ | ~_00345_;
	assign _00470_ = _00468_ & ~_00469_;
	assign _00471_ = _00349_ & ~_00470_;
	assign _00472_ = \mchip.design.vga.v_idx [8] & ~_00471_;
	assign _00473_ = _00469_ | ~_00467_;
	assign _00474_ = \mchip.design.vga.v_idx [8] & ~_00473_;
	assign _00475_ = _00474_ | _00472_;
	assign _00476_ = _00399_ | _00298_;
	assign _00477_ = _00476_ | ~_00398_;
	assign _00478_ = _00477_ | _00352_;
	assign _00479_ = ~_00301_;
	assign _00480_ = _00299_ & ~_00366_;
	assign _00481_ = _00341_ & ~_00480_;
	assign _00482_ = ~(_00481_ | _00395_);
	assign _00483_ = _00479_ & ~_00482_;
	assign _00484_ = _00483_ | _00352_;
	assign _00485_ = _00478_ & ~_00484_;
	assign _00486_ = _00475_ & ~_00485_;
	assign _00487_ = _00466_ & ~_00486_;
	assign _00488_ = ~(_00331_ | _00299_);
	assign _00489_ = _00301_ & ~_00317_;
	assign _00490_ = ~(_00489_ & _00488_);
	assign _00491_ = \mchip.design.vga.v_idx [8] & ~_00490_;
	assign _00492_ = _00299_ | ~_00333_;
	assign _00493_ = _00489_ & ~_00492_;
	assign _00494_ = _00493_ | _00479_;
	assign _00495_ = \mchip.design.vga.v_idx [8] & ~_00494_;
	assign _00496_ = _00495_ | _00491_;
	assign _00497_ = _00366_ | ~_00301_;
	assign _00498_ = _00339_ & ~_00497_;
	assign _00499_ = _00305_ & ~_00498_;
	assign _00500_ = \mchip.design.vga.v_idx [8] & ~_00499_;
	assign _00501_ = _00498_ & ~_00352_;
	assign _00502_ = _00500_ & ~_00501_;
	assign _00503_ = _00496_ & ~_00502_;
	assign _00504_ = _00487_ & ~_00503_;
	assign _00505_ = \mchip.design.vga.h_idx [9] & ~\mchip.design.vga.h_idx [8];
	assign _00506_ = \mchip.design.vga.h_idx [6] & ~\mchip.design.vga.h_idx [7];
	assign _00507_ = ~(_00506_ & \mchip.design.vga.h_idx [5]);
	assign _00508_ = _00507_ & ~\mchip.design.vga.h_idx [7];
	assign _00509_ = \mchip.design.vga.h_idx [5] | ~\mchip.design.vga.h_idx [4];
	assign _00510_ = _00506_ & ~_00509_;
	assign _00511_ = ~(\mchip.design.vga.h_idx [0] & \mchip.design.vga.h_idx [1]);
	assign _00512_ = _00511_ & ~_03793_;
	assign _00513_ = _00510_ & ~_00512_;
	assign _00514_ = _00508_ & ~_00513_;
	assign _00515_ = _00505_ & ~_00514_;
	assign _00516_ = _00515_ | _03750_;
	assign _00517_ = ~(_00511_ | _03793_);
	assign _00518_ = ~(_00517_ & _00510_);
	assign _00519_ = _00505_ & ~_00518_;
	assign _00520_ = _00519_ | _00516_;
	assign _00521_ = \mchip.design.vga.h_idx [5] & \mchip.design.vga.h_idx [4];
	assign _00522_ = _00521_ & _00506_;
	assign _00523_ = ~(\mchip.design.vga.h_idx [2] & \mchip.design.vga.h_idx [3]);
	assign _00524_ = ~(_00523_ | _00511_);
	assign _00525_ = ~(_00524_ & _00522_);
	assign _00526_ = _00505_ & ~_00525_;
	assign _00527_ = _00313_ & ~_00526_;
	assign _00528_ = _00520_ & ~_00527_;
	assign _00529_ = \mchip.design.vga.h_idx [8] & ~\mchip.design.vga.h_idx [9];
	assign _00530_ = \mchip.design.vga.h_idx [0] | ~\mchip.design.vga.h_idx [1];
	assign _00531_ = _00530_ | _00523_;
	assign _00532_ = ~(\mchip.design.vga.h_idx [6] & \mchip.design.vga.h_idx [7]);
	assign _00533_ = _00532_ | ~_00521_;
	assign _00534_ = _00533_ | _00531_;
	assign _00535_ = _00529_ & ~_00534_;
	assign _00536_ = ~(\mchip.design.vga.h_idx [9] | \mchip.design.vga.h_idx [8]);
	assign _00537_ = ~_00536_;
	assign _00538_ = _00521_ & ~_00532_;
	assign _00539_ = _00523_ | _00511_;
	assign _00540_ = _00539_ & ~_00533_;
	assign _00541_ = _00538_ & ~_00540_;
	assign _00542_ = _00529_ & ~_00541_;
	assign _00543_ = _00537_ & ~_00542_;
	assign _00544_ = _00543_ | _00535_;
	assign _00545_ = _00312_ & ~\mchip.design.vga.h_idx [6];
	assign _00546_ = \mchip.design.vga.h_idx [6] | ~\mchip.design.vga.h_idx [5];
	assign _00547_ = _00312_ & ~_00546_;
	assign _00548_ = ~\mchip.design.vga.h_idx [4];
	assign _00549_ = \mchip.design.vga.h_idx [1] | \mchip.design.vga.h_idx [2];
	assign _00550_ = \mchip.design.vga.h_idx [4] | ~\mchip.design.vga.h_idx [3];
	assign _00551_ = _00549_ & ~_00550_;
	assign _00552_ = _00548_ & ~_00551_;
	assign _00553_ = _00547_ & ~_00552_;
	assign _00554_ = _00545_ & ~_00553_;
	assign _00555_ = \mchip.design.vga.h_idx [9] & ~_00554_;
	assign _00556_ = \mchip.design.vga.h_idx [2] | ~\mchip.design.vga.h_idx [3];
	assign _00557_ = _00556_ | _00530_;
	assign _00558_ = _00557_ | _03782_;
	assign _00559_ = _00505_ & ~_00558_;
	assign _00560_ = _00555_ & ~_00559_;
	assign _00561_ = _00544_ & ~_00560_;
	assign _00562_ = \mchip.design.vga.h_idx [1] | ~\mchip.design.vga.h_idx [0];
	assign _00563_ = ~(_00562_ | _00556_);
	assign _00564_ = \mchip.design.vga.h_idx [6] | ~\mchip.design.vga.h_idx [7];
	assign _00565_ = ~(_00564_ | _03771_);
	assign _00566_ = ~(_00565_ & _00563_);
	assign _00567_ = _00529_ & ~_00566_;
	assign _00568_ = _03847_ & ~_03868_;
	assign _00569_ = _00550_ | _00549_;
	assign _00570_ = \mchip.design.vga.h_idx [4] | \mchip.design.vga.h_idx [3];
	assign _00571_ = ~(_00570_ & _00569_);
	assign _00572_ = _00546_ | ~_03847_;
	assign _00573_ = _00571_ & ~_00572_;
	assign _00574_ = _00568_ & ~_00573_;
	assign _00575_ = _00574_ | \mchip.design.vga.h_idx [9];
	assign _00576_ = _00575_ | _00567_;
	assign _00577_ = ~_00529_;
	assign _00578_ = _00532_ | _00509_;
	assign _00579_ = \mchip.design.vga.h_idx [3] | ~\mchip.design.vga.h_idx [2];
	assign _00580_ = _00579_ | _00562_;
	assign _00581_ = _00580_ | _00578_;
	assign _00582_ = _00581_ | _00577_;
	assign _00583_ = ~\mchip.design.vga.h_idx [9];
	assign _00584_ = _03847_ & \mchip.design.vga.h_idx [6];
	assign _00585_ = \mchip.design.vga.h_idx [5] | ~\mchip.design.vga.h_idx [6];
	assign _00586_ = _03847_ & ~_00585_;
	assign _00587_ = \mchip.design.vga.h_idx [1] & \mchip.design.vga.h_idx [2];
	assign _00588_ = \mchip.design.vga.h_idx [3] | ~\mchip.design.vga.h_idx [4];
	assign _00589_ = ~(_00588_ | _00587_);
	assign _00590_ = \mchip.design.vga.h_idx [4] & ~_00589_;
	assign _00591_ = _00586_ & ~_00590_;
	assign _00592_ = _00584_ & ~_00591_;
	assign _00593_ = _00583_ & ~_00592_;
	assign _00594_ = _00582_ & ~_00593_;
	assign _00595_ = _00576_ & ~_00594_;
	assign _00596_ = ~(_00579_ | _03804_);
	assign _00597_ = ~(_00596_ & _00510_);
	assign _00598_ = _00529_ & ~_00597_;
	assign _00599_ = ~(\mchip.design.vga.h_idx [5] | \mchip.design.vga.h_idx [4]);
	assign _00600_ = _00599_ & _00506_;
	assign _00601_ = _03760_ & ~_00600_;
	assign _00602_ = _03793_ & ~_00596_;
	assign _00603_ = _00510_ & ~_00602_;
	assign _00604_ = _00601_ & ~_00603_;
	assign _00605_ = _00529_ & ~_00604_;
	assign _00606_ = _00537_ & ~_00605_;
	assign _00607_ = _00606_ | _00598_;
	assign _00608_ = _00564_ | ~_00599_;
	assign _00609_ = ~(_00608_ | _03814_);
	assign _00610_ = ~(_00609_ & _00529_);
	assign _00611_ = \mchip.design.vga.h_idx [7] & ~_00609_;
	assign _00612_ = _00529_ & ~_00611_;
	assign _00613_ = _00612_ | _00536_;
	assign _00614_ = _00610_ & ~_00613_;
	assign _00615_ = _00607_ & ~_00614_;
	assign _00616_ = _00524_ & ~_00533_;
	assign _00617_ = _00616_ | _00537_;
	assign _00618_ = ~(\mchip.design.vga.h_idx [6] | \mchip.design.vga.h_idx [7]);
	assign _00619_ = _00618_ & ~_03771_;
	assign _00620_ = ~(_00556_ | _00511_);
	assign _00621_ = ~(_00620_ & _00619_);
	assign _00622_ = _00621_ | _00577_;
	assign _00623_ = _00529_ & ~_03760_;
	assign _00624_ = _00523_ & ~_03771_;
	assign _00625_ = \mchip.design.vga.h_idx [5] & ~_00624_;
	assign _00626_ = _00623_ & ~_00625_;
	assign _00627_ = _00626_ | _00536_;
	assign _00628_ = _00622_ & ~_00627_;
	assign _00629_ = _00617_ & ~_00628_;
	assign _00630_ = _00557_ | ~_00565_;
	assign _00631_ = _00536_ & ~_00630_;
	assign _00632_ = ~\mchip.design.vga.h_idx [5];
	assign _00633_ = _00632_ & ~_00564_;
	assign _00634_ = \mchip.design.vga.h_idx [7] & ~_00633_;
	assign _00635_ = _00511_ & ~_00556_;
	assign _00636_ = \mchip.design.vga.h_idx [3] & ~_00635_;
	assign _00637_ = _00565_ & ~_00636_;
	assign _00638_ = _00634_ & ~_00637_;
	assign _00639_ = _00638_ | _00537_;
	assign _00640_ = _00639_ | _00631_;
	assign _00641_ = _00579_ | _00530_;
	assign _00642_ = _00641_ | _00578_;
	assign _00643_ = _00642_ | ~_00536_;
	assign _00644_ = _00511_ & ~_00579_;
	assign _00645_ = _03793_ & ~_00644_;
	assign _00646_ = _00645_ | _00578_;
	assign _00647_ = _00599_ | _00532_;
	assign _00648_ = _00646_ & ~_00647_;
	assign _00649_ = _00536_ & ~_00648_;
	assign _00650_ = _00643_ & ~_00649_;
	assign _00651_ = _00640_ & ~_00650_;
	assign _00652_ = _00580_ | ~_00510_;
	assign _00653_ = _00536_ & ~_00652_;
	assign _00654_ = \mchip.design.vga.h_idx [6] | ~_00312_;
	assign _00655_ = _00312_ & ~_00585_;
	assign _00656_ = _00655_ & ~_00590_;
	assign _00657_ = _00654_ & ~_00656_;
	assign _00658_ = _00657_ | \mchip.design.vga.h_idx [9];
	assign _00659_ = _00658_ | _00653_;
	assign _00660_ = _00562_ | _03793_;
	assign _00661_ = _00660_ | _00608_;
	assign _00662_ = _00661_ | _00537_;
	assign _00663_ = ~_00312_;
	assign _00664_ = _00570_ | _00549_;
	assign _00665_ = \mchip.design.vga.h_idx [8] | ~\mchip.design.vga.h_idx [7];
	assign _00666_ = _03868_ & ~_00665_;
	assign _00667_ = _00666_ & ~_00664_;
	assign _00668_ = _00663_ & ~_00667_;
	assign _00669_ = _00583_ & ~_00668_;
	assign _00670_ = _00662_ & ~_00669_;
	assign _00671_ = _00659_ & ~_00670_;
	assign _00672_ = _03804_ & ~_00523_;
	assign _00673_ = _00672_ | _03782_;
	assign _00674_ = _00632_ & ~_03760_;
	assign _00675_ = _00673_ & ~_00674_;
	assign _00676_ = _00536_ & ~_00675_;
	assign _00677_ = _00523_ | _03804_;
	assign _00678_ = _00677_ | _03782_;
	assign _00679_ = _00536_ & ~_00678_;
	assign _00680_ = _00679_ | _00676_;
	assign _00681_ = _00680_ | _00671_;
	assign _00682_ = _00681_ | _00651_;
	assign _00683_ = _00682_ | _00629_;
	assign _00684_ = _00683_ | _00615_;
	assign _00685_ = _00684_ | _00595_;
	assign _00686_ = _00685_ | _00561_;
	assign _00687_ = _00686_ | _00528_;
	assign _00688_ = _00504_ & ~_00687_;
	assign \mchip.design.board.is_board  = ~_00688_;
	assign _00689_ = _00530_ | _03793_;
	assign _00690_ = _00689_ | _00608_;
	assign _00691_ = _00536_ & ~_00690_;
	assign _00692_ = _00512_ & ~_00608_;
	assign _00693_ = \mchip.design.vga.h_idx [7] & ~_00692_;
	assign _00694_ = _00693_ | _00537_;
	assign _00695_ = _00694_ | _00691_;
	assign _00696_ = _00566_ | _00537_;
	assign _00697_ = _00663_ & ~_00666_;
	assign _00698_ = _00665_ | _00546_;
	assign _00699_ = _00571_ & ~_00698_;
	assign _00700_ = _00697_ & ~_00699_;
	assign _00701_ = _00583_ & ~_00700_;
	assign _00702_ = _00696_ & ~_00701_;
	assign _00703_ = _00695_ & ~_00702_;
	assign _00704_ = _00424_ | ~_00360_;
	assign _00705_ = _00424_ & _00360_;
	assign _00706_ = \mchip.design.vga.v_idx [4] | ~\mchip.design.vga.v_idx [3];
	assign _00707_ = _00430_ & ~_00706_;
	assign _00708_ = _00429_ & ~_00707_;
	assign _00709_ = _00705_ & ~_00708_;
	assign _00710_ = _00704_ & ~_00709_;
	assign _00711_ = _00461_ | _00382_;
	assign _00712_ = _00352_ & ~_00711_;
	assign _00713_ = _00712_ | _00710_;
	assign _00714_ = ~(_00399_ | _00314_);
	assign _00715_ = ~(_00714_ & _00398_);
	assign _00716_ = _00715_ | \mchip.design.vga.v_idx [8];
	assign _00717_ = \mchip.design.vga.v_idx [3] | ~\mchip.design.vga.v_idx [4];
	assign _00718_ = _00363_ & ~_00717_;
	assign _00719_ = _00718_ | _00338_;
	assign _00720_ = _00425_ | _00359_;
	assign _00721_ = _00719_ & ~_00720_;
	assign _00722_ = _00721_ | _00360_;
	assign _00723_ = _00716_ & ~_00722_;
	assign _00724_ = _00713_ & ~_00723_;
	assign _00725_ = _00724_ & _00703_;
	assign _00726_ = ~(_00312_ & _03868_);
	assign _00727_ = ~(_00587_ | _00550_);
	assign _00728_ = _00570_ & ~_00727_;
	assign _00729_ = _00547_ & ~_00728_;
	assign _00730_ = _00726_ & ~_00729_;
	assign _00731_ = _00730_ | \mchip.design.vga.h_idx [9];
	assign _00732_ = _00562_ | _00523_;
	assign _00733_ = _00732_ | _03782_;
	assign _00734_ = _00536_ & ~_00733_;
	assign _00735_ = _00734_ | _00731_;
	assign _00736_ = _00597_ | _00537_;
	assign _00737_ = _00536_ & ~_00604_;
	assign _00738_ = _00736_ & ~_00737_;
	assign _00739_ = _00735_ & ~_00738_;
	assign _00740_ = _00739_ & _00724_;
	assign _00741_ = ~(_00740_ | _00725_);
	assign _00742_ = ~(\mchip.design.vga.h_idx [4] & \mchip.design.vga.h_idx [3]);
	assign _00743_ = _00742_ & ~_00585_;
	assign _00744_ = _00743_ | ~\mchip.design.vga.h_idx [6];
	assign _00745_ = _00744_ & ~_00665_;
	assign _00746_ = _00663_ & ~_00745_;
	assign _00747_ = _00746_ | \mchip.design.vga.h_idx [9];
	assign _00748_ = _00579_ | _00511_;
	assign _00749_ = _00748_ | _00578_;
	assign _00750_ = _00536_ & ~_00749_;
	assign _00751_ = _00750_ | _00747_;
	assign _00752_ = _00537_ | _00534_;
	assign _00753_ = _00536_ & ~_00541_;
	assign _00754_ = _00752_ & ~_00753_;
	assign _00755_ = _00751_ & ~_00754_;
	assign _00756_ = _00755_ & _00724_;
	assign _00757_ = _00741_ & ~_00756_;
	assign _00758_ = _00529_ & ~_00678_;
	assign _00759_ = _00529_ & ~_00675_;
	assign _00760_ = _00537_ & ~_00759_;
	assign _00761_ = _00760_ | _00758_;
	assign _00762_ = _00577_ | _00518_;
	assign _00763_ = _00529_ & _00506_;
	assign _00764_ = ~_00599_;
	assign _00765_ = ~(_00509_ | _03793_);
	assign _00766_ = _00764_ & ~_00765_;
	assign _00767_ = _00763_ & ~_00766_;
	assign _00768_ = _00623_ | _00536_;
	assign _00769_ = _00768_ | _00767_;
	assign _00770_ = _00762_ & ~_00769_;
	assign _00771_ = _00761_ & ~_00770_;
	assign _00772_ = _00771_ & _00724_;
	assign _00773_ = _00757_ & ~_00772_;
	assign _00774_ = _03868_ & _03847_;
	assign _00775_ = _00774_ & ~_00664_;
	assign _00776_ = _03847_ & ~_00775_;
	assign _00777_ = _00776_ | \mchip.design.vga.h_idx [9];
	assign _00778_ = _00529_ & ~_00661_;
	assign _00779_ = _00778_ | _00777_;
	assign _00780_ = ~(_00556_ | _03804_);
	assign _00781_ = ~(_00780_ & _00565_);
	assign _00782_ = _00781_ | _00577_;
	assign _00783_ = \mchip.design.vga.h_idx [3] & ~_00780_;
	assign _00784_ = _00565_ & ~_00783_;
	assign _00785_ = _00634_ & ~_00784_;
	assign _00786_ = _00529_ & ~_00785_;
	assign _00787_ = _00786_ | _00536_;
	assign _00788_ = _00782_ & ~_00787_;
	assign _00789_ = _00779_ & ~_00788_;
	assign _00790_ = _00789_ & _00724_;
	assign _00791_ = _00773_ & ~_00790_;
	assign _00792_ = _00529_ & ~_00642_;
	assign _00793_ = _00529_ & ~_00648_;
	assign _00794_ = _00537_ & ~_00793_;
	assign _00795_ = _00794_ | _00792_;
	assign _00796_ = _00732_ | _00533_;
	assign _00797_ = _00796_ | _00577_;
	assign _00798_ = ~(\mchip.design.vga.h_idx [5] & \mchip.design.vga.h_idx [6]);
	assign _00799_ = _03847_ & ~_00798_;
	assign _00800_ = _00587_ & ~_00742_;
	assign _00801_ = _00799_ & ~_00800_;
	assign _00802_ = _00799_ & ~_00801_;
	assign _00803_ = _00583_ & ~_00802_;
	assign _00804_ = _00797_ & ~_00803_;
	assign _00805_ = _00795_ & ~_00804_;
	assign _00806_ = _00805_ & _00724_;
	assign _00807_ = _00791_ & ~_00806_;
	assign _00808_ = _00618_ & ~_00521_;
	assign _00809_ = _00523_ & ~_00620_;
	assign _00810_ = _00619_ & ~_00809_;
	assign _00811_ = _00808_ & ~_00810_;
	assign _00812_ = _00505_ & ~_00811_;
	assign _00813_ = ~(_00812_ | _03750_);
	assign _00814_ = _00505_ & ~_00621_;
	assign _00815_ = _00814_ | ~_00813_;
	assign _00816_ = _00510_ & ~_00689_;
	assign _00817_ = ~(_00816_ & _00505_);
	assign _00818_ = _00798_ & _00312_;
	assign _00819_ = _00549_ & ~_00588_;
	assign _00820_ = _00742_ & ~_00819_;
	assign _00821_ = _00655_ & ~_00820_;
	assign _00822_ = _00818_ & ~_00821_;
	assign _00823_ = _00822_ | _00583_;
	assign _00824_ = _00817_ & ~_00823_;
	assign _00825_ = _00815_ & ~_00824_;
	assign _00826_ = _00825_ & _00724_;
	assign _00827_ = _00807_ & ~_00826_;
	assign _00828_ = _00377_ | _00331_;
	assign _00829_ = _00828_ | ~_00376_;
	assign _00830_ = _00829_ | \mchip.design.vga.v_idx [8];
	assign _00831_ = _00333_ & ~_00377_;
	assign _00832_ = \mchip.design.vga.v_idx [3] & ~_00831_;
	assign _00833_ = _00376_ & ~_00832_;
	assign _00834_ = _00833_ | ~_00318_;
	assign _00835_ = _00834_ & ~\mchip.design.vga.v_idx [8];
	assign _00836_ = _00830_ & ~_00835_;
	assign _00837_ = _00435_ | _00367_;
	assign _00838_ = _00837_ | \mchip.design.vga.v_idx [8];
	assign _00839_ = ~(_00339_ | _00367_);
	assign _00840_ = _00319_ & ~_00839_;
	assign _00841_ = _00840_ | \mchip.design.vga.v_idx [8];
	assign _00842_ = _00838_ & ~_00841_;
	assign _00843_ = _00842_ | _00836_;
	assign _00844_ = _00825_ & ~_00843_;
	assign _00845_ = _00805_ & ~_00843_;
	assign _00846_ = _00789_ & ~_00843_;
	assign _00847_ = _00771_ & ~_00843_;
	assign _00848_ = _00755_ & ~_00843_;
	assign _00849_ = _00703_ & ~_00843_;
	assign _00850_ = _00739_ & ~_00843_;
	assign _00851_ = _00850_ | _00849_;
	assign _00852_ = _00851_ | _00848_;
	assign _00853_ = _00852_ | _00847_;
	assign _00854_ = _00853_ | _00846_;
	assign _00855_ = _00854_ | _00845_;
	assign _00856_ = _00855_ | _00844_;
	assign _00857_ = _00827_ & ~_00856_;
	assign _00858_ = ~(_00448_ & _00378_);
	assign _00859_ = _00858_ | _00352_;
	assign _00860_ = ~(_00345_ | _00318_);
	assign _00861_ = _00455_ & ~_00378_;
	assign _00862_ = _00448_ & ~_00861_;
	assign _00863_ = _00860_ & ~_00862_;
	assign _00864_ = _00863_ | _00352_;
	assign _00865_ = _00859_ & ~_00864_;
	assign _00866_ = _00865_ | _00356_;
	assign _00867_ = _00825_ & ~_00866_;
	assign _00868_ = _00805_ & ~_00866_;
	assign _00869_ = _00789_ & ~_00866_;
	assign _00870_ = _00771_ & ~_00866_;
	assign _00871_ = _00755_ & ~_00866_;
	assign _00872_ = _00703_ & ~_00866_;
	assign _00873_ = _00739_ & ~_00866_;
	assign _00874_ = _00873_ | _00872_;
	assign _00875_ = _00874_ | _00871_;
	assign _00876_ = _00875_ | _00870_;
	assign _00877_ = _00876_ | _00869_;
	assign _00878_ = _00877_ | _00868_;
	assign _00879_ = _00878_ | _00867_;
	assign _00880_ = _00304_ | \mchip.design.vga.v_idx [8];
	assign _00881_ = _00352_ & ~_00306_;
	assign _00882_ = _00880_ & ~_00881_;
	assign _00883_ = _00476_ | _00409_;
	assign _00884_ = _00883_ | \mchip.design.vga.v_idx [8];
	assign _00885_ = ~(_00395_ | _00345_);
	assign _00886_ = \mchip.design.vga.v_idx [7] & ~_00885_;
	assign _00887_ = ~(_00476_ & _00299_);
	assign _00888_ = _00887_ & ~_00409_;
	assign _00889_ = _00886_ & ~_00888_;
	assign _00890_ = _00889_ | \mchip.design.vga.v_idx [8];
	assign _00891_ = _00884_ & ~_00890_;
	assign _00892_ = _00891_ | _00882_;
	assign _00893_ = _00825_ & ~_00892_;
	assign _00894_ = _00805_ & ~_00892_;
	assign _00895_ = _00789_ & ~_00892_;
	assign _00896_ = _00771_ & ~_00892_;
	assign _00897_ = _00755_ & ~_00892_;
	assign _00898_ = _00703_ & ~_00892_;
	assign _00899_ = _00739_ & ~_00892_;
	assign _00900_ = _00899_ | _00898_;
	assign _00901_ = _00900_ | _00897_;
	assign _00902_ = _00901_ | _00896_;
	assign _00903_ = _00902_ | _00895_;
	assign _00904_ = _00903_ | _00894_;
	assign _00905_ = _00904_ | _00893_;
	assign _00906_ = _00879_ | ~_00905_;
	assign _00907_ = ~(_00317_ & _00301_);
	assign _00908_ = ~(_00299_ | _00298_);
	assign _00909_ = _00489_ & ~_00908_;
	assign _00910_ = _00907_ & ~_00909_;
	assign _00911_ = \mchip.design.vga.v_idx [8] & ~_00910_;
	assign _00912_ = _00420_ | ~_00489_;
	assign _00913_ = \mchip.design.vga.v_idx [8] & ~_00912_;
	assign _00914_ = _00911_ & ~_00913_;
	assign _00915_ = _00715_ | _00352_;
	assign _00916_ = \mchip.design.vga.v_idx [5] & ~_00395_;
	assign _00917_ = _00479_ & ~_00916_;
	assign _00918_ = _00298_ & ~_00399_;
	assign _00919_ = _00335_ & ~_00918_;
	assign _00920_ = _00398_ & ~_00919_;
	assign _00921_ = _00917_ & ~_00920_;
	assign _00922_ = \mchip.design.vga.v_idx [8] & ~_00921_;
	assign _00923_ = _00915_ & ~_00922_;
	assign _00924_ = _00923_ | _00914_;
	assign _00925_ = _00825_ & ~_00924_;
	assign _00926_ = _00805_ & ~_00924_;
	assign _00927_ = _00789_ & ~_00924_;
	assign _00928_ = _00771_ & ~_00924_;
	assign _00929_ = _00755_ & ~_00924_;
	assign _00930_ = _00703_ & ~_00924_;
	assign _00931_ = _00739_ & ~_00924_;
	assign _00932_ = _00931_ | _00930_;
	assign _00933_ = _00932_ | _00929_;
	assign _00934_ = _00933_ | _00928_;
	assign _00935_ = _00934_ | _00927_;
	assign _00936_ = _00935_ | _00926_;
	assign _00937_ = ~(_00936_ | _00925_);
	assign _00938_ = \mchip.design.vga.v_idx [7] | ~\mchip.design.vga.v_idx [8];
	assign _00939_ = _00424_ & ~_00938_;
	assign _00940_ = _00717_ | _00363_;
	assign _00941_ = _00940_ & ~_00362_;
	assign _00942_ = _00939_ & ~_00941_;
	assign _00943_ = \mchip.design.vga.v_idx [7] & \mchip.design.vga.v_idx [8];
	assign _00944_ = _00943_ | _00942_;
	assign _00945_ = _00469_ | _00405_;
	assign _00946_ = \mchip.design.vga.v_idx [8] & ~_00945_;
	assign _00947_ = _00944_ & ~_00946_;
	assign _00948_ = _00829_ | _00352_;
	assign _00949_ = \mchip.design.vga.v_idx [8] & ~_00834_;
	assign _00950_ = _00948_ & ~_00949_;
	assign _00951_ = _00950_ | _00947_;
	assign _00952_ = _00825_ & ~_00951_;
	assign _00953_ = _00805_ & ~_00951_;
	assign _00954_ = _00789_ & ~_00951_;
	assign _00955_ = _00771_ & ~_00951_;
	assign _00956_ = _00755_ & ~_00951_;
	assign _00957_ = _00703_ & ~_00951_;
	assign _00958_ = _00739_ & ~_00951_;
	assign _00959_ = _00958_ | _00957_;
	assign _00960_ = _00959_ | _00956_;
	assign _00961_ = _00960_ | _00955_;
	assign _00962_ = _00961_ | _00954_;
	assign _00963_ = _00962_ | _00953_;
	assign _00964_ = _00963_ | _00952_;
	assign _00965_ = _00964_ | ~_00937_;
	assign _00966_ = _00965_ | _00906_;
	assign _00967_ = _00966_ | ~_00857_;
	assign _00968_ = _00905_ | ~_00879_;
	assign _00969_ = _00968_ | _00965_;
	assign _00970_ = _00857_ & ~_00969_;
	assign _00971_ = _00970_ | ~_00967_;
	assign _00972_ = ~(_00964_ & _00937_);
	assign _00973_ = _00905_ | _00879_;
	assign _00974_ = _00973_ | _00972_;
	assign _00975_ = _00974_ | ~_00857_;
	assign _00976_ = _00964_ | _00937_;
	assign _00977_ = _00976_ | _00973_;
	assign _00978_ = _00857_ & ~_00977_;
	assign _00979_ = _00975_ & ~_00978_;
	assign _00980_ = _00971_ & ~_00979_;
	assign _00981_ = _00848_ | _00756_;
	assign _00982_ = _00981_ | _00897_;
	assign _00983_ = _00982_ | _00871_;
	assign _00984_ = _00983_ | _00956_;
	assign _00985_ = ~(_00984_ | _00929_);
	assign _00986_ = _00849_ | _00725_;
	assign _00987_ = _00986_ | _00898_;
	assign _00988_ = _00987_ | _00872_;
	assign _00989_ = _00988_ | _00957_;
	assign _00990_ = _00989_ | _00930_;
	assign _00991_ = _00985_ & ~_00990_;
	assign _00992_ = _00850_ | _00740_;
	assign _00993_ = _00992_ | _00899_;
	assign _00994_ = _00993_ | _00873_;
	assign _00995_ = _00994_ | _00958_;
	assign _00996_ = _00995_ | _00931_;
	assign _00997_ = _00991_ & ~_00996_;
	assign _00998_ = _00847_ | _00772_;
	assign _00999_ = _00998_ | _00896_;
	assign _01000_ = _00999_ | _00870_;
	assign _01001_ = _01000_ | _00955_;
	assign _01002_ = _01001_ | _00928_;
	assign _01003_ = _00846_ | _00790_;
	assign _01004_ = _01003_ | _00895_;
	assign _01005_ = _01004_ | _00869_;
	assign _01006_ = _01005_ | _00954_;
	assign _01007_ = _01006_ | _00927_;
	assign _01008_ = _01002_ | ~_01007_;
	assign _01009_ = _00845_ | _00806_;
	assign _01010_ = _01009_ | _00894_;
	assign _01011_ = _01010_ | _00868_;
	assign _01012_ = _01011_ | _00953_;
	assign _01013_ = ~(_01012_ | _00926_);
	assign _01014_ = _00844_ | _00826_;
	assign _01015_ = _01014_ | _00893_;
	assign _01016_ = _01015_ | _00867_;
	assign _01017_ = _01016_ | _00952_;
	assign _01018_ = _01017_ | _00925_;
	assign _01019_ = _01018_ | ~_01013_;
	assign _01020_ = _01019_ | _01008_;
	assign _01021_ = _00997_ & ~_01020_;
	assign _01022_ = _01018_ | _01013_;
	assign _01023_ = _01007_ | _01002_;
	assign _01024_ = _01023_ | _01022_;
	assign _01025_ = _00997_ & ~_01024_;
	assign _01026_ = ~(_01018_ & _01013_);
	assign _01027_ = _01026_ | _01023_;
	assign _01028_ = _00997_ & ~_01027_;
	assign _01029_ = _01028_ | _01025_;
	assign _01030_ = ~(_01029_ | _01021_);
	assign _01031_ = ~(_01023_ | _01019_);
	assign _01032_ = ~(_00990_ & _00985_);
	assign _01033_ = ~(_01032_ | _00996_);
	assign _01034_ = ~(_01033_ & _01031_);
	assign _01035_ = _00990_ | _00985_;
	assign _01036_ = _01035_ | _00996_;
	assign _01037_ = _01031_ & ~_01036_;
	assign _01038_ = _01034_ & ~_01037_;
	assign _01039_ = _01007_ | ~_01002_;
	assign _01040_ = _01039_ | _01019_;
	assign _01041_ = _00997_ & ~_01040_;
	assign _01042_ = _01041_ | _01021_;
	assign _01043_ = _01042_ | _01029_;
	assign _01044_ = _01043_ | ~_01038_;
	assign _01045_ = _01041_ | _01025_;
	assign _01046_ = _01034_ & ~_01045_;
	assign _01047_ = _01044_ & ~_01046_;
	assign _01048_ = _01041_ | _01028_;
	assign _01049_ = ~(_01048_ | _01037_);
	assign _01050_ = _01049_ | ~_01044_;
	assign _01051_ = _01047_ & ~_01050_;
	assign _01052_ = _01051_ & ~_01030_;
	assign _01053_ = _01052_ ^ _00980_;
	assign _01054_ = ~_00980_;
	assign _01055_ = ~(_01052_ & _00980_);
	assign _01056_ = _00979_ ^ _00971_;
	assign _01057_ = _01056_ & _01053_;
	assign _01058_ = _01055_ & ~_01057_;
	assign _01059_ = (_01053_ ? _01058_ : _01054_);
	assign _01060_ = _01053_ ^ _00980_;
	assign _01061_ = _01059_ | ~_01060_;
	assign _01062_ = ~(_01060_ ^ _01059_);
	assign _01063_ = ~(_00973_ | _00965_);
	assign _01064_ = _00856_ | _00827_;
	assign _01065_ = _01063_ & ~_01064_;
	assign _01066_ = _00971_ & _01053_;
	assign _01067_ = _01055_ & ~_01066_;
	assign _01068_ = ~(_01056_ ^ _01053_);
	assign _01069_ = _01068_ | _01067_;
	assign _01070_ = _01068_ ^ _01067_;
	assign _01071_ = _01070_ & ~_01054_;
	assign _01072_ = _01069_ & ~_01071_;
	assign _01073_ = _01053_ ^ _01054_;
	assign _01074_ = _01073_ ^ _01058_;
	assign _01075_ = _01074_ ^ _00980_;
	assign _01076_ = _01072_ | ~_01075_;
	assign _01077_ = ~(_01075_ ^ _01072_);
	assign _01078_ = _01051_ ^ _01030_;
	assign _01079_ = ~(_01078_ & _01056_);
	assign _01080_ = _00979_ & ~_00971_;
	assign _01081_ = _01065_ | ~_01080_;
	assign _01082_ = _00978_ | _00970_;
	assign _01083_ = ~(_01082_ | _01065_);
	assign _01084_ = _01081_ & ~_01083_;
	assign _01085_ = _01078_ ^ _01056_;
	assign _01086_ = _01085_ & ~_01084_;
	assign _01087_ = _01079_ & ~_01086_;
	assign _01088_ = ~(_00971_ ^ _01053_);
	assign _01089_ = _01088_ | _01087_;
	assign _01090_ = _01088_ ^ _01087_;
	assign _01091_ = _01090_ & _01056_;
	assign _01092_ = _01089_ & ~_01091_;
	assign _01093_ = _01070_ ^ _00980_;
	assign _01094_ = _01092_ | ~_01093_;
	assign _01095_ = _01077_ & ~_01094_;
	assign _01096_ = _01076_ & ~_01095_;
	assign _01097_ = _01093_ ^ _01092_;
	assign _01098_ = _01077_ & ~_01097_;
	assign _01099_ = ~(_01085_ ^ _01084_);
	assign _01100_ = ~(_01050_ ^ _01047_);
	assign _01101_ = _00971_ & ~_01100_;
	assign _01102_ = ~(_01101_ & _01099_);
	assign _01103_ = _01101_ ^ _01099_;
	assign _01104_ = _01103_ & _00971_;
	assign _01105_ = _01104_ | ~_01102_;
	assign _01106_ = _01090_ ^ _01056_;
	assign _01107_ = ~(_01106_ & _01105_);
	assign _01108_ = _01106_ ^ _01105_;
	assign _01109_ = ~(_01100_ ^ _00971_);
	assign _01110_ = _01047_ & ~_01084_;
	assign _01111_ = _01110_ & _01109_;
	assign _01112_ = _01110_ ^ _01109_;
	assign _01113_ = _01112_ & ~_01084_;
	assign _01114_ = _01113_ | _01111_;
	assign _01115_ = ~(_01103_ ^ _00971_);
	assign _01116_ = _01115_ | ~_01114_;
	assign _01117_ = _01108_ & ~_01116_;
	assign _01118_ = _01107_ & ~_01117_;
	assign _01119_ = _01098_ & ~_01118_;
	assign _01120_ = _01096_ & ~_01119_;
	assign _01121_ = _01062_ & ~_01120_;
	assign _01122_ = _01061_ & ~_01121_;
	assign _01123_ = ~(_01122_ ^ _01053_);
	assign _01124_ = _01084_ ^ _01047_;
	assign _01125_ = (_01124_ ? _05810_ : _05809_);
	assign _01126_ = ~(_01125_ | _01123_);
	assign _01127_ = ~(_01112_ ^ _01084_);
	assign _01128_ = _01126_ & ~_01127_;
	assign _01129_ = ~(_01115_ ^ _01114_);
	assign _01130_ = _01128_ & ~_01129_;
	assign _01131_ = ~(_01116_ ^ _01108_);
	assign _01132_ = (_01124_ ? _05813_ : _05812_);
	assign _01133_ = (_01124_ ? _05815_ : _05816_);
	assign _01134_ = (_01127_ ? _01132_ : _01133_);
	assign _01135_ = (_01124_ ? _05820_ : _05819_);
	assign _01136_ = (_01124_ ? _05822_ : _05823_);
	assign _01137_ = (_01127_ ? _01135_ : _01136_);
	assign _01138_ = (_01129_ ? _01134_ : _01137_);
	assign _01139_ = ~(_01138_ | _01123_);
	assign _01140_ = (_01131_ ? _01130_ : _01139_);
	assign _01141_ = _01118_ ^ _01097_;
	assign _01142_ = _01140_ & ~_01141_;
	assign _01143_ = ~(_01118_ | _01097_);
	assign _01144_ = _01143_ | ~_01094_;
	assign _01145_ = _01144_ ^ _01077_;
	assign _01146_ = (_01124_ ? _05886_ : _05887_);
	assign _01147_ = (_01124_ ? _05889_ : _05890_);
	assign _01148_ = (_01127_ ? _01146_ : _01147_);
	assign _01149_ = (_01124_ ? _05893_ : _05894_);
	assign _01150_ = (_01124_ ? _05896_ : _05897_);
	assign _01151_ = (_01127_ ? _01149_ : _01150_);
	assign _01152_ = (_01129_ ? _01148_ : _01151_);
	assign _01153_ = (_01124_ ? _05901_ : _05902_);
	assign _01154_ = (_01124_ ? _05904_ : _05905_);
	assign _01155_ = (_01127_ ? _01153_ : _01154_);
	assign _01156_ = (_01124_ ? _05908_ : _05909_);
	assign _01157_ = (_01124_ ? _05911_ : _05912_);
	assign _01158_ = (_01127_ ? _01156_ : _01157_);
	assign _01159_ = (_01129_ ? _01155_ : _01158_);
	assign _01160_ = (_01131_ ? _01152_ : _01159_);
	assign _01161_ = (_01124_ ? _05778_ : _05779_);
	assign _01162_ = (_01124_ ? _05781_ : _05782_);
	assign _01163_ = (_01127_ ? _01161_ : _01162_);
	assign _01164_ = (_01124_ ? _05785_ : _05786_);
	assign _01165_ = (_01124_ ? _05788_ : _05789_);
	assign _01166_ = (_01127_ ? _01164_ : _01165_);
	assign _01167_ = (_01129_ ? _01163_ : _01166_);
	assign _01168_ = (_01124_ ? _05793_ : _05794_);
	assign _01169_ = (_01124_ ? _05796_ : _05797_);
	assign _01170_ = (_01127_ ? _01168_ : _01169_);
	assign _01171_ = (_01124_ ? _05800_ : _05801_);
	assign _01172_ = (_01124_ ? _05803_ : _05804_);
	assign _01173_ = (_01127_ ? _01171_ : _01172_);
	assign _01174_ = (_01129_ ? _01170_ : _01173_);
	assign _01175_ = (_01131_ ? _01167_ : _01174_);
	assign _01176_ = (_01141_ ? _01160_ : _01175_);
	assign _01177_ = ~(_01176_ | _01123_);
	assign _01178_ = (_01145_ ? _01142_ : _01177_);
	assign _01179_ = ~(_01120_ ^ _01062_);
	assign _01180_ = _01178_ & ~_01179_;
	assign _01181_ = (_01124_ ? _05748_ : _05742_);
	assign _01182_ = _01181_ | _01123_;
	assign _01183_ = _01182_ | _01127_;
	assign _01184_ = _01183_ | _01129_;
	assign _01185_ = (_01124_ ? _05764_ : _05763_);
	assign _01186_ = (_01124_ ? _05766_ : _05767_);
	assign _01187_ = (_01127_ ? _01185_ : _01186_);
	assign _01188_ = (_01124_ ? _05771_ : _05770_);
	assign _01189_ = (_01124_ ? _05773_ : _05774_);
	assign _01190_ = (_01127_ ? _01188_ : _01189_);
	assign _01191_ = (_01129_ ? _01187_ : _01190_);
	assign _01192_ = _01191_ | _01123_;
	assign _01193_ = (_01131_ ? _01184_ : _01192_);
	assign _01194_ = _01193_ | _01141_;
	assign _01195_ = (_01124_ ? _05833_ : _05834_);
	assign _01196_ = (_01124_ ? _05837_ : _05838_);
	assign _01197_ = (_01127_ ? _01195_ : _01196_);
	assign _01198_ = (_01124_ ? _05842_ : _05843_);
	assign _01199_ = (_01124_ ? _05845_ : _05846_);
	assign _01200_ = (_01127_ ? _01198_ : _01199_);
	assign _01201_ = (_01129_ ? _01197_ : _01200_);
	assign _01202_ = (_01124_ ? _05852_ : _05853_);
	assign _01203_ = (_01124_ ? _05855_ : _05856_);
	assign _01204_ = (_01127_ ? _01202_ : _01203_);
	assign _01205_ = (_01124_ ? _05859_ : _05860_);
	assign _01206_ = (_01124_ ? _05862_ : _05863_);
	assign _01207_ = (_01127_ ? _01205_ : _01206_);
	assign _01208_ = (_01129_ ? _01204_ : _01207_);
	assign _01209_ = (_01131_ ? _01201_ : _01208_);
	assign _01210_ = (_01124_ ? _05389_ : _05399_);
	assign _01211_ = (_01124_ ? _05453_ : _05464_);
	assign _01212_ = (_01127_ ? _01210_ : _01211_);
	assign _01213_ = (_01124_ ? _05505_ : _05516_);
	assign _01214_ = (_01124_ ? _05538_ : _05548_);
	assign _01215_ = (_01127_ ? _01213_ : _01214_);
	assign _01216_ = (_01129_ ? _01212_ : _01215_);
	assign _01217_ = (_01124_ ? _05613_ : _05623_);
	assign _01218_ = (_01124_ ? _05645_ : _05654_);
	assign _01219_ = (_01127_ ? _01217_ : _01218_);
	assign _01220_ = (_01124_ ? _05684_ : _05691_);
	assign _01221_ = (_01124_ ? _05705_ : _05712_);
	assign _01222_ = (_01127_ ? _01220_ : _01221_);
	assign _01223_ = (_01129_ ? _01219_ : _01222_);
	assign _01224_ = (_01131_ ? _01216_ : _01223_);
	assign _01225_ = (_01141_ ? _01209_ : _01224_);
	assign _01226_ = _01225_ | _01123_;
	assign _01227_ = (_01145_ ? _01194_ : _01226_);
	assign _01228_ = _01227_ | _01179_;
	assign _01229_ = ~(_01228_ & _01180_);
	assign _01230_ = _00905_ | ~_00857_;
	assign _01231_ = _01230_ | _00879_;
	assign _01232_ = _01231_ | _00964_;
	assign _01233_ = _00937_ & ~_01232_;
	assign _01234_ = _01233_ | _01229_;
	assign _01235_ = ~(_01228_ | _01180_);
	assign _01236_ = _01235_ & ~_01233_;
	assign _01237_ = _01234_ & ~_01236_;
	assign io_out[5] = _00688_ & ~_01237_;
	assign _01238_ = _01236_ | _01234_;
	assign io_out[7] = _00688_ & ~_01238_;
	assign _01239_ = _00202_ | _05836_;
	assign _01240_ = ~(_01239_ | _05260_);
	assign _01241_ = _00210_ | _00204_;
	assign _01242_ = _01240_ & ~_01241_;
	assign _01243_ = _00212_ | ~_01242_;
	assign _01244_ = _01241_ | _00212_;
	assign _01245_ = _01244_ | ~_01240_;
	assign _01246_ = \mchip.design.owner.fsm.currState  | ~\mchip.design.currStateConfirm [1];
	assign _01247_ = _01246_ | _01245_;
	assign _01248_ = _01247_ | _05260_;
	assign _01249_ = _05335_ | ~_05260_;
	assign _01250_ = ~(_01249_ & _05346_);
	assign _01251_ = _01250_ | _01248_;
	assign _01252_ = _00202_ ^ _05421_;
	assign _01253_ = _01252_ | _01251_;
	assign _01254_ = ~(_01240_ ^ _00204_);
	assign _01255_ = _01254_ | _01253_;
	assign _01256_ = _01240_ & ~_00204_;
	assign _01257_ = ~(_01256_ ^ _00210_);
	assign _01258_ = _01257_ | _01255_;
	assign _01259_ = _00212_ & ~_01242_;
	assign _01260_ = ~(_01258_ | _01243_);
	assign _01261_ = _01259_ | ~_01243_;
	assign _01262_ = _01245_ | _05260_;
	assign _01263_ = _01262_ | _01250_;
	assign _01264_ = _01263_ | _01252_;
	assign _01265_ = _01264_ | _01254_;
	assign _01266_ = _01265_ | _01257_;
	assign _01267_ = _01266_ | ~_01261_;
	assign _01268_ = ~(_01267_ | _01243_);
	assign _01269_ = \mchip.design.owner.tokens [0] & ~_01268_;
	assign _01270_ = _01269_ | _01260_;
	assign _01271_ = _05260_ & ~_05944_;
	assign _01272_ = _00140_ | _00137_;
	assign _01273_ = _01271_ & ~_01272_;
	assign _01274_ = _00134_ | ~_01273_;
	assign _01275_ = _01272_ | _00134_;
	assign _01276_ = _01275_ | ~_01271_;
	assign _01277_ = _01276_ | _01246_;
	assign _01278_ = _01277_ | ~_05260_;
	assign _01279_ = _01278_ | _06010_;
	assign _01280_ = _01279_ | ~_00202_;
	assign _01281_ = ~(_01271_ ^ _00137_);
	assign _01282_ = _01281_ | _01280_;
	assign _01283_ = _01271_ & ~_00137_;
	assign _01284_ = ~(_01283_ ^ _00140_);
	assign _01285_ = _01284_ | _01282_;
	assign _01286_ = _00134_ & ~_01273_;
	assign _01287_ = ~(_01285_ | _01274_);
	assign _01288_ = _01286_ | ~_01274_;
	assign _01289_ = _01276_ | ~_05260_;
	assign _01290_ = _01289_ | _06010_;
	assign _01291_ = _01290_ | ~_00202_;
	assign _01292_ = _01291_ | _01281_;
	assign _01293_ = _01292_ | _01284_;
	assign _01294_ = _01293_ | ~_01288_;
	assign _01295_ = ~(_01294_ | _01274_);
	assign _01296_ = \mchip.design.owner.tokens [0] & ~_01295_;
	assign _01297_ = _01296_ | _01287_;
	assign _01298_ = (_00199_ ? _01270_ : _01297_);
	assign _01299_ = _04767_ | _06010_;
	assign _01300_ = ~(_01299_ | _05260_);
	assign _01301_ = _06022_ | _01341_;
	assign _01302_ = _01300_ & ~_01301_;
	assign _01303_ = _06008_ | ~_01302_;
	assign _01304_ = _01301_ | _06008_;
	assign _01305_ = _01304_ | ~_01300_;
	assign _01306_ = _01305_ | _01246_;
	assign _01307_ = _01306_ | _05260_;
	assign _01308_ = _01307_ | ~_05442_;
	assign _01310_ = _01309_ | _01308_;
	assign _01311_ = ~(_01300_ ^ _01341_);
	assign _01312_ = _01311_ | _01310_;
	assign _01313_ = _01300_ & ~_01341_;
	assign _01314_ = ~(_01313_ ^ _06022_);
	assign _01315_ = _01314_ | _01312_;
	assign _01316_ = _06008_ & ~_01302_;
	assign _01317_ = ~(_01315_ | _01303_);
	assign _01318_ = _01316_ | ~_01303_;
	assign _01319_ = _01305_ | _05260_;
	assign _01320_ = _01319_ | ~_05442_;
	assign _01321_ = _01320_ | _01309_;
	assign _01322_ = _01321_ | _01311_;
	assign _01323_ = _01322_ | _01314_;
	assign _01324_ = _01323_ | ~_01318_;
	assign _01325_ = ~(_01324_ | _01303_);
	assign _01326_ = \mchip.design.owner.tokens [0] & ~_01325_;
	assign _01327_ = _01326_ | _01317_;
	assign _01328_ = (_00131_ ? _01298_ : _01327_);
	assign _01329_ = _01246_ | _05941_;
	assign _01330_ = _05260_ & ~_05943_;
	assign _01331_ = _05953_ | _05947_;
	assign _01332_ = _05955_ | _05941_;
	assign _01333_ = _01332_ | _01331_;
	assign _01334_ = _01330_ & ~_01333_;
	assign _01335_ = ~(_01334_ ^ _05941_);
	assign _01336_ = _01335_ | _01329_;
	assign _01337_ = _01336_ | ~_05260_;
	assign _01338_ = ~(_01337_ | _05836_);
	assign _01339_ = _01249_ ^ _05945_;
	assign _01340_ = _01338_ & ~_01339_;
	assign _01342_ = _01340_ & ~_01341_;
	assign _01344_ = _01342_ & ~_01343_;
	assign _01345_ = _01330_ & ~_01331_;
	assign _01346_ = _01345_ ^ _05955_;
	assign _01347_ = _01346_ & _01344_;
	assign _01348_ = _05955_ | ~_01345_;
	assign _01349_ = _01348_ ^ _05941_;
	assign _01350_ = _01347_ & ~_01349_;
	assign _01351_ = _05941_ | ~_01334_;
	assign _01352_ = _01351_ | ~_05260_;
	assign _01353_ = _01352_ | _05836_;
	assign _01354_ = _01353_ | _01339_;
	assign _01355_ = _01354_ | _01341_;
	assign _01356_ = _01355_ | _01343_;
	assign _01357_ = _01356_ | ~_01346_;
	assign _01358_ = ~(_01357_ | _01349_);
	assign _01359_ = \mchip.design.owner.tokens [0] & ~_01358_;
	assign _01360_ = _01359_ | _01350_;
	assign _01361_ = (_06005_ ? _01328_ : _01360_);
	assign _01362_ = _01246_ | _05832_;
	assign _01363_ = _05841_ | _05836_;
	assign _01364_ = ~(_01363_ | _05260_);
	assign _01365_ = _05868_ | _05851_;
	assign _01366_ = _01365_ | _05832_;
	assign _01367_ = _01364_ & ~_01366_;
	assign _01368_ = ~(_01367_ ^ _05832_);
	assign _01369_ = _01368_ | _01362_;
	assign _01370_ = _01369_ | _05260_;
	assign _01371_ = ~(_01370_ | _01250_);
	assign _01372_ = _05841_ ^ _05421_;
	assign _01373_ = _01371_ & ~_01372_;
	assign _01374_ = ~(_01364_ ^ _05851_);
	assign _01375_ = _01373_ & ~_01374_;
	assign _01376_ = _01364_ & ~_05851_;
	assign _01377_ = ~(_01376_ ^ _05868_);
	assign _01378_ = _01375_ & ~_01377_;
	assign _01379_ = _01364_ & ~_01365_;
	assign _01380_ = _01379_ ^ _05832_;
	assign _01381_ = _01380_ & _01378_;
	assign _01382_ = ~(_01379_ | _05832_);
	assign _01383_ = _01381_ & ~_01382_;
	assign _01384_ = _05832_ | ~_01367_;
	assign _01385_ = _01384_ | _05260_;
	assign _01386_ = _01385_ | _01250_;
	assign _01387_ = _01386_ | _01372_;
	assign _01388_ = _01387_ | _01374_;
	assign _01389_ = _01388_ | _01377_;
	assign _01390_ = _01389_ | ~_01380_;
	assign _01391_ = ~(_01390_ | _01382_);
	assign _01392_ = \mchip.design.owner.tokens [0] & ~_01391_;
	assign _01393_ = _01392_ | _01383_;
	assign _01394_ = (_05934_ ? _01361_ : _01393_);
	assign _01395_ = ~(_05602_ | _05378_);
	assign _01396_ = ~(_05938_ & _05260_);
	assign _01397_ = _01395_ & ~_01396_;
	assign _01398_ = _01397_ ^ _05378_;
	assign _01399_ = _01246_ | _05378_;
	assign _01400_ = _01399_ | ~_01398_;
	assign _01401_ = _01400_ | ~_05260_;
	assign _01402_ = _01401_ | _06010_;
	assign _01403_ = _01402_ | ~_05841_;
	assign _01404_ = _01396_ ^ _05602_;
	assign _01405_ = _01404_ | _01403_;
	assign _01406_ = ~(_01396_ | _05602_);
	assign _01407_ = ~(_01406_ ^ _05378_);
	assign _01408_ = _01407_ | _01405_;
	assign _01409_ = _01398_ & ~_01408_;
	assign _01410_ = ~(_01397_ | _05378_);
	assign _01411_ = _01409_ & ~_01410_;
	assign _01412_ = _05378_ | ~_01397_;
	assign _01413_ = _01412_ | ~_05260_;
	assign _01414_ = _01413_ | _06010_;
	assign _01415_ = _01414_ | ~_05841_;
	assign _01416_ = _01415_ | _01404_;
	assign _01417_ = _01416_ | _01407_;
	assign _01418_ = _01417_ | ~_01398_;
	assign _01419_ = ~(_01418_ | _01410_);
	assign _01420_ = \mchip.design.owner.tokens [0] & ~_01419_;
	assign _01421_ = _01420_ | _01411_;
	assign _00012_ = (_05827_ ? _01394_ : _01421_);
	assign _01422_ = ~(_00249_ & \mchip.design.owner.fsm.currState );
	assign _01423_ = _01422_ | _01245_;
	assign _01424_ = _01423_ | _05260_;
	assign _01425_ = _01424_ | _01250_;
	assign _01426_ = _01425_ | _01252_;
	assign _01427_ = _01426_ | _01254_;
	assign _01428_ = _01427_ | _01257_;
	assign _01429_ = _01428_ | ~_01261_;
	assign _01430_ = ~(_01429_ | _01243_);
	assign _01431_ = \mchip.design.owner.tokens [1] & ~_01268_;
	assign _01432_ = _01431_ | _01430_;
	assign _01433_ = _01422_ | _01276_;
	assign _01434_ = _01433_ | ~_05260_;
	assign _01435_ = _01434_ | _06010_;
	assign _01436_ = _01435_ | ~_00202_;
	assign _01437_ = _01436_ | _01281_;
	assign _01438_ = _01437_ | _01284_;
	assign _01439_ = _01438_ | ~_01288_;
	assign _01440_ = ~(_01439_ | _01274_);
	assign _01441_ = \mchip.design.owner.tokens [1] & ~_01295_;
	assign _01442_ = _01441_ | _01440_;
	assign _01443_ = (_00199_ ? _01432_ : _01442_);
	assign _01444_ = _01422_ | _01305_;
	assign _01445_ = _01444_ | _05260_;
	assign _01446_ = _01445_ | ~_05442_;
	assign _01447_ = _01446_ | _01309_;
	assign _01448_ = _01447_ | _01311_;
	assign _01449_ = _01448_ | _01314_;
	assign _01450_ = _01449_ | ~_01318_;
	assign _01451_ = ~(_01450_ | _01303_);
	assign _01452_ = \mchip.design.owner.tokens [1] & ~_01325_;
	assign _01453_ = _01452_ | _01451_;
	assign _01454_ = (_00131_ ? _01443_ : _01453_);
	assign _01455_ = _01422_ | _05941_;
	assign _01456_ = _01455_ | _01335_;
	assign _01457_ = _01456_ | ~_05260_;
	assign _01458_ = _01457_ | _05836_;
	assign _01459_ = _01458_ | _01339_;
	assign _01460_ = _01459_ | _01341_;
	assign _01461_ = _01460_ | _01343_;
	assign _01462_ = _01461_ | ~_01346_;
	assign _01463_ = ~(_01462_ | _01349_);
	assign _01464_ = \mchip.design.owner.tokens [1] & ~_01358_;
	assign _01465_ = _01464_ | _01463_;
	assign _01466_ = (_06005_ ? _01454_ : _01465_);
	assign _01467_ = _01422_ | _05832_;
	assign _01468_ = _01467_ | _01368_;
	assign _01469_ = _01468_ | _05260_;
	assign _01470_ = _01469_ | _01250_;
	assign _01471_ = _01470_ | _01372_;
	assign _01472_ = _01471_ | _01374_;
	assign _01473_ = _01472_ | _01377_;
	assign _01474_ = _01473_ | ~_01380_;
	assign _01475_ = ~(_01474_ | _01382_);
	assign _01476_ = \mchip.design.owner.tokens [1] & ~_01391_;
	assign _01477_ = _01476_ | _01475_;
	assign _01478_ = (_05934_ ? _01466_ : _01477_);
	assign _01479_ = _01422_ | _05378_;
	assign _01480_ = _01479_ | ~_01398_;
	assign _01481_ = _01480_ | ~_05260_;
	assign _01482_ = _01481_ | _06010_;
	assign _01483_ = _01482_ | ~_05841_;
	assign _01484_ = _01483_ | _01404_;
	assign _01485_ = _01484_ | _01407_;
	assign _01486_ = _01485_ | ~_01398_;
	assign _01487_ = ~(_01486_ | _01410_);
	assign _01488_ = \mchip.design.owner.tokens [1] & ~_01419_;
	assign _01489_ = _01488_ | _01487_;
	assign _00023_ = (_05827_ ? _01478_ : _01489_);
	assign _01490_ = ~_01257_;
	assign _01491_ = _01246_ | ~_01245_;
	assign _01492_ = _01491_ | ~_05260_;
	assign _01493_ = _01492_ | ~_01250_;
	assign _01494_ = _01493_ | ~_01252_;
	assign _01495_ = _01494_ | ~_01254_;
	assign _01496_ = _01495_ | _01490_;
	assign _01497_ = _01496_ | _01261_;
	assign _01498_ = _01243_ & ~_01497_;
	assign _01499_ = _01249_ | ~_01252_;
	assign _01500_ = _01499_ | ~_01254_;
	assign _01501_ = _01500_ | ~_01257_;
	assign _01502_ = _01501_ | _01261_;
	assign _01503_ = _01243_ & ~_01502_;
	assign _01504_ = \mchip.design.owner.tokens [2] & ~_01503_;
	assign _01505_ = _01504_ | _01498_;
	assign _01506_ = ~_01284_;
	assign _01507_ = _01246_ | ~_01276_;
	assign _01508_ = _01507_ | _05260_;
	assign _01509_ = _01508_ | ~_06010_;
	assign _01510_ = _01509_ | _00202_;
	assign _01511_ = _01510_ | ~_01281_;
	assign _01512_ = _01511_ | _01506_;
	assign _01513_ = _01512_ | _01288_;
	assign _01514_ = _01274_ & ~_01513_;
	assign _01515_ = _00202_ | _05421_;
	assign _01516_ = _01515_ | ~_01281_;
	assign _01517_ = _01516_ | ~_01284_;
	assign _01518_ = _01517_ | _01288_;
	assign _01519_ = _01274_ & ~_01518_;
	assign _01520_ = \mchip.design.owner.tokens [2] & ~_01519_;
	assign _01521_ = _01520_ | _01514_;
	assign _01522_ = (_00199_ ? _01505_ : _01521_);
	assign _01523_ = ~_01314_;
	assign _01524_ = _01246_ | ~_01305_;
	assign _01525_ = _01524_ | ~_05260_;
	assign _01526_ = _01525_ | _05442_;
	assign _01527_ = _01526_ | ~_01309_;
	assign _01528_ = _01527_ | ~_01311_;
	assign _01529_ = _01528_ | _01523_;
	assign _01530_ = _01529_ | _01318_;
	assign _01531_ = _01303_ & ~_01530_;
	assign _01532_ = _05431_ | ~_01309_;
	assign _01533_ = _01532_ | ~_01311_;
	assign _01534_ = _01533_ | ~_01314_;
	assign _01535_ = _01534_ | _01318_;
	assign _01536_ = _01303_ & ~_01535_;
	assign _01537_ = \mchip.design.owner.tokens [2] & ~_01536_;
	assign _01538_ = _01537_ | _01531_;
	assign _01539_ = (_00131_ ? _01522_ : _01538_);
	assign _01540_ = ~_01343_;
	assign _01541_ = _01334_ ^ _05941_;
	assign _01542_ = _01541_ | _01329_;
	assign _01543_ = _01542_ | _05260_;
	assign _01544_ = _01543_ | ~_05836_;
	assign _01545_ = _01544_ | ~_01339_;
	assign _01546_ = _01545_ | ~_01341_;
	assign _01547_ = _01546_ | _01540_;
	assign _01548_ = _01547_ | _01346_;
	assign _01549_ = _01349_ & ~_01548_;
	assign _01550_ = _05346_ | ~_01339_;
	assign _01551_ = _01550_ | ~_01341_;
	assign _01552_ = _01551_ | _01540_;
	assign _01553_ = _01552_ | _01346_;
	assign _01554_ = _01349_ & ~_01553_;
	assign _01555_ = \mchip.design.owner.tokens [2] & ~_01554_;
	assign _01556_ = _01555_ | _01549_;
	assign _01557_ = (_06005_ ? _01539_ : _01556_);
	assign _01558_ = _01367_ ^ _05832_;
	assign _01559_ = _01558_ | _01362_;
	assign _01560_ = _01559_ | ~_05260_;
	assign _01561_ = _01560_ | ~_01250_;
	assign _01562_ = _01561_ | ~_01372_;
	assign _01563_ = _01562_ | ~_01374_;
	assign _01564_ = _01563_ | ~_01377_;
	assign _01565_ = _01564_ | _01380_;
	assign _01566_ = _01382_ & ~_01565_;
	assign _01567_ = _01249_ | ~_01372_;
	assign _01568_ = _01567_ | ~_01374_;
	assign _01569_ = _01568_ | ~_01377_;
	assign _01570_ = _01569_ | _01380_;
	assign _01571_ = _01382_ & ~_01570_;
	assign _01572_ = \mchip.design.owner.tokens [2] & ~_01571_;
	assign _01573_ = _01572_ | _01566_;
	assign _01574_ = (_05934_ ? _01557_ : _01573_);
	assign _01575_ = ~_01407_;
	assign _01576_ = _01399_ | _01398_;
	assign _01577_ = _01576_ | _05260_;
	assign _01578_ = _01577_ | ~_06010_;
	assign _01579_ = _01578_ | _05841_;
	assign _01580_ = _01579_ | ~_01404_;
	assign _01581_ = _01580_ | _01575_;
	assign _01582_ = _01581_ | _01398_;
	assign _01583_ = _01410_ & ~_01582_;
	assign _01584_ = _05378_ | _05260_;
	assign _01585_ = _01584_ | ~_06010_;
	assign _01586_ = _01585_ | _05841_;
	assign _01587_ = _01586_ | ~_01404_;
	assign _01588_ = _01587_ | _01575_;
	assign _01589_ = _01588_ | _01398_;
	assign _01590_ = _01410_ & ~_01589_;
	assign _01591_ = \mchip.design.owner.tokens [2] & ~_01590_;
	assign _01592_ = _01591_ | _01583_;
	assign _00034_ = (_05827_ ? _01574_ : _01592_);
	assign _01593_ = _01422_ | ~_01245_;
	assign _01594_ = _01593_ | ~_05260_;
	assign _01595_ = _01594_ | ~_01250_;
	assign _01596_ = _01595_ | ~_01252_;
	assign _01597_ = _01596_ | ~_01254_;
	assign _01598_ = _01597_ | _01490_;
	assign _01599_ = _01598_ | _01261_;
	assign _01600_ = _01243_ & ~_01599_;
	assign _01601_ = \mchip.design.owner.tokens [3] & ~_01503_;
	assign _01602_ = _01601_ | _01600_;
	assign _01603_ = _01422_ | ~_01276_;
	assign _01604_ = _01603_ | _05260_;
	assign _01605_ = _01604_ | ~_06010_;
	assign _01606_ = _01605_ | _00202_;
	assign _01607_ = _01606_ | ~_01281_;
	assign _01608_ = _01607_ | _01506_;
	assign _01609_ = _01608_ | _01288_;
	assign _01610_ = _01274_ & ~_01609_;
	assign _01611_ = \mchip.design.owner.tokens [3] & ~_01519_;
	assign _01612_ = _01611_ | _01610_;
	assign _01613_ = (_00199_ ? _01602_ : _01612_);
	assign _01614_ = _01422_ | ~_01305_;
	assign _01615_ = _01614_ | ~_05260_;
	assign _01616_ = _01615_ | _05442_;
	assign _01617_ = _01616_ | ~_01309_;
	assign _01618_ = _01617_ | ~_01311_;
	assign _01619_ = _01618_ | _01523_;
	assign _01620_ = _01619_ | _01318_;
	assign _01621_ = _01303_ & ~_01620_;
	assign _01622_ = \mchip.design.owner.tokens [3] & ~_01536_;
	assign _01623_ = _01622_ | _01621_;
	assign _01624_ = (_00131_ ? _01613_ : _01623_);
	assign _01625_ = _01455_ | _01541_;
	assign _01626_ = _01625_ | _05260_;
	assign _01627_ = _01626_ | ~_05836_;
	assign _01628_ = _01627_ | ~_01339_;
	assign _01629_ = _01628_ | ~_01341_;
	assign _01630_ = _01629_ | _01540_;
	assign _01631_ = _01630_ | _01346_;
	assign _01632_ = _01349_ & ~_01631_;
	assign _01633_ = \mchip.design.owner.tokens [3] & ~_01554_;
	assign _01634_ = _01633_ | _01632_;
	assign _01635_ = (_06005_ ? _01624_ : _01634_);
	assign _01636_ = _01558_ | _01467_;
	assign _01637_ = _01636_ | ~_05260_;
	assign _01638_ = _01637_ | ~_01250_;
	assign _01639_ = _01638_ | ~_01372_;
	assign _01640_ = _01639_ | ~_01374_;
	assign _01641_ = _01640_ | ~_01377_;
	assign _01642_ = _01641_ | _01380_;
	assign _01643_ = _01382_ & ~_01642_;
	assign _01644_ = \mchip.design.owner.tokens [3] & ~_01571_;
	assign _01645_ = _01644_ | _01643_;
	assign _01646_ = (_05934_ ? _01635_ : _01645_);
	assign _01647_ = _01479_ | _01398_;
	assign _01648_ = _01647_ | _05260_;
	assign _01649_ = _01648_ | ~_06010_;
	assign _01650_ = _01649_ | _05841_;
	assign _01651_ = _01650_ | ~_01404_;
	assign _01652_ = _01651_ | _01575_;
	assign _01653_ = _01652_ | _01398_;
	assign _01654_ = _01410_ & ~_01653_;
	assign _01655_ = \mchip.design.owner.tokens [3] & ~_01590_;
	assign _01656_ = _01655_ | _01654_;
	assign _00045_ = (_05827_ ? _01646_ : _01656_);
	assign _01657_ = _01491_ | _05260_;
	assign _01658_ = _01657_ | ~_01250_;
	assign _01659_ = _01658_ | ~_01252_;
	assign _01660_ = _01659_ | ~_01254_;
	assign _01661_ = _01660_ | _01490_;
	assign _01662_ = _01661_ | _01261_;
	assign _01663_ = _01243_ & ~_01662_;
	assign _01664_ = _05346_ | ~_01252_;
	assign _01665_ = _01664_ | ~_01254_;
	assign _01666_ = _01665_ | ~_01257_;
	assign _01667_ = _01666_ | _01261_;
	assign _01668_ = _01243_ & ~_01667_;
	assign _01669_ = \mchip.design.owner.tokens [4] & ~_01668_;
	assign _01670_ = _01669_ | _01663_;
	assign _01671_ = _01507_ | ~_05260_;
	assign _01672_ = _01671_ | ~_06010_;
	assign _01673_ = _01672_ | _00202_;
	assign _01674_ = _01673_ | ~_01281_;
	assign _01675_ = _01674_ | _01506_;
	assign _01676_ = _01675_ | _01288_;
	assign _01677_ = _01274_ & ~_01676_;
	assign _01678_ = _01249_ | _00202_;
	assign _01679_ = _01678_ | ~_01281_;
	assign _01680_ = _01679_ | ~_01284_;
	assign _01681_ = _01680_ | _01288_;
	assign _01682_ = _01274_ & ~_01681_;
	assign _01683_ = \mchip.design.owner.tokens [4] & ~_01682_;
	assign _01684_ = _01683_ | _01677_;
	assign _01685_ = (_00199_ ? _01670_ : _01684_);
	assign _01686_ = _01524_ | _05260_;
	assign _01687_ = _01686_ | _05442_;
	assign _01688_ = _01687_ | ~_01309_;
	assign _01689_ = _01688_ | ~_01311_;
	assign _01690_ = _01689_ | _01523_;
	assign _01691_ = _01690_ | _01318_;
	assign _01692_ = _01303_ & ~_01691_;
	assign _01693_ = _05421_ | ~_01309_;
	assign _01694_ = _01693_ | ~_01311_;
	assign _01695_ = _01694_ | ~_01314_;
	assign _01696_ = _01695_ | _01318_;
	assign _01697_ = _01303_ & ~_01696_;
	assign _01698_ = \mchip.design.owner.tokens [4] & ~_01697_;
	assign _01699_ = _01698_ | _01692_;
	assign _01700_ = (_00131_ ? _01685_ : _01699_);
	assign _01701_ = _01542_ | ~_05260_;
	assign _01702_ = _01701_ | ~_05836_;
	assign _01703_ = _01702_ | ~_01339_;
	assign _01704_ = _01703_ | ~_01341_;
	assign _01705_ = _01704_ | _01540_;
	assign _01706_ = _01705_ | _01346_;
	assign _01707_ = _01349_ & ~_01706_;
	assign _01708_ = _05431_ | ~_01339_;
	assign _01709_ = _01708_ | ~_01341_;
	assign _01710_ = _01709_ | _01540_;
	assign _01711_ = _01710_ | _01346_;
	assign _01712_ = _01349_ & ~_01711_;
	assign _01713_ = \mchip.design.owner.tokens [4] & ~_01712_;
	assign _01714_ = _01713_ | _01707_;
	assign _01715_ = (_06005_ ? _01700_ : _01714_);
	assign _01716_ = _01559_ | _05260_;
	assign _01717_ = _01716_ | ~_01250_;
	assign _01718_ = _01717_ | ~_01372_;
	assign _01719_ = _01718_ | ~_01374_;
	assign _01720_ = _01719_ | ~_01377_;
	assign _01721_ = _01720_ | _01380_;
	assign _01722_ = _01382_ & ~_01721_;
	assign _01723_ = _01367_ | _05832_;
	assign _01724_ = _01723_ | _05260_;
	assign _01725_ = _01724_ | ~_01250_;
	assign _01726_ = _01725_ | ~_01372_;
	assign _01727_ = _01726_ | ~_01374_;
	assign _01728_ = _01727_ | ~_01377_;
	assign _01729_ = _01728_ | _01380_;
	assign _01730_ = _01382_ & ~_01729_;
	assign _01731_ = \mchip.design.owner.tokens [4] & ~_01730_;
	assign _01732_ = _01731_ | _01722_;
	assign _01733_ = (_05934_ ? _01715_ : _01732_);
	assign _01734_ = _01576_ | ~_05260_;
	assign _01735_ = _01734_ | ~_06010_;
	assign _01736_ = _01735_ | _05841_;
	assign _01737_ = _01736_ | ~_01404_;
	assign _01738_ = _01737_ | _01575_;
	assign _01739_ = _01738_ | _01398_;
	assign _01740_ = _01410_ & ~_01739_;
	assign _01741_ = ~(_01410_ & _05260_);
	assign _01742_ = _01741_ | ~_06010_;
	assign _01743_ = _01742_ | _05841_;
	assign _01744_ = _01743_ | ~_01404_;
	assign _01745_ = _01744_ | _01575_;
	assign _01746_ = _01745_ | _01398_;
	assign _01747_ = _01410_ & ~_01746_;
	assign _01748_ = \mchip.design.owner.tokens [4] & ~_01747_;
	assign _01749_ = _01748_ | _01740_;
	assign _00056_ = (_05827_ ? _01733_ : _01749_);
	assign _01750_ = _01593_ | _05260_;
	assign _01751_ = _01750_ | ~_01250_;
	assign _01752_ = _01751_ | ~_01252_;
	assign _01753_ = _01752_ | ~_01254_;
	assign _01754_ = _01753_ | _01490_;
	assign _01755_ = _01754_ | _01261_;
	assign _01756_ = _01243_ & ~_01755_;
	assign _01757_ = \mchip.design.owner.tokens [5] & ~_01668_;
	assign _01758_ = _01757_ | _01756_;
	assign _01759_ = _01603_ | ~_05260_;
	assign _01760_ = _01759_ | ~_06010_;
	assign _01761_ = _01760_ | _00202_;
	assign _01762_ = _01761_ | ~_01281_;
	assign _01763_ = _01762_ | _01506_;
	assign _01764_ = _01763_ | _01288_;
	assign _01765_ = _01274_ & ~_01764_;
	assign _01766_ = \mchip.design.owner.tokens [5] & ~_01682_;
	assign _01767_ = _01766_ | _01765_;
	assign _01768_ = (_00199_ ? _01758_ : _01767_);
	assign _01769_ = _01614_ | _05260_;
	assign _01770_ = _01769_ | _05442_;
	assign _01771_ = _01770_ | ~_01309_;
	assign _01772_ = _01771_ | ~_01311_;
	assign _01773_ = _01772_ | _01523_;
	assign _01774_ = _01773_ | _01318_;
	assign _01775_ = _01303_ & ~_01774_;
	assign _01776_ = \mchip.design.owner.tokens [5] & ~_01697_;
	assign _01777_ = _01776_ | _01775_;
	assign _01778_ = (_00131_ ? _01768_ : _01777_);
	assign _01779_ = _01625_ | ~_05260_;
	assign _01780_ = _01779_ | ~_05836_;
	assign _01781_ = _01780_ | ~_01339_;
	assign _01782_ = _01781_ | ~_01341_;
	assign _01783_ = _01782_ | _01540_;
	assign _01784_ = _01783_ | _01346_;
	assign _01785_ = _01349_ & ~_01784_;
	assign _01786_ = \mchip.design.owner.tokens [5] & ~_01712_;
	assign _01787_ = _01786_ | _01785_;
	assign _01788_ = (_06005_ ? _01778_ : _01787_);
	assign _01789_ = _01636_ | _05260_;
	assign _01790_ = _01789_ | ~_01250_;
	assign _01791_ = _01790_ | ~_01372_;
	assign _01792_ = _01791_ | ~_01374_;
	assign _01793_ = _01792_ | ~_01377_;
	assign _01794_ = _01793_ | _01380_;
	assign _01795_ = _01382_ & ~_01794_;
	assign _01796_ = \mchip.design.owner.tokens [5] & ~_01730_;
	assign _01797_ = _01796_ | _01795_;
	assign _01798_ = (_05934_ ? _01788_ : _01797_);
	assign _01799_ = _01647_ | ~_05260_;
	assign _01800_ = _01799_ | ~_06010_;
	assign _01801_ = _01800_ | _05841_;
	assign _01802_ = _01801_ | ~_01404_;
	assign _01803_ = _01802_ | _01575_;
	assign _01804_ = _01803_ | _01398_;
	assign _01805_ = _01410_ & ~_01804_;
	assign _01806_ = \mchip.design.owner.tokens [5] & ~_01747_;
	assign _01807_ = _01806_ | _01805_;
	assign _00067_ = (_05827_ ? _01798_ : _01807_);
	assign _01808_ = _01492_ | _01250_;
	assign _01809_ = _01808_ | ~_01252_;
	assign _01810_ = _01809_ | ~_01254_;
	assign _01811_ = _01810_ | _01490_;
	assign _01812_ = _01811_ | _01261_;
	assign _01813_ = _01243_ & ~_01812_;
	assign _01814_ = _05431_ | ~_01252_;
	assign _01815_ = _01814_ | ~_01254_;
	assign _01816_ = _01815_ | ~_01257_;
	assign _01817_ = _01816_ | _01261_;
	assign _01818_ = _01243_ & ~_01817_;
	assign _01819_ = \mchip.design.owner.tokens [6] & ~_01818_;
	assign _01820_ = _01819_ | _01813_;
	assign _01821_ = _01508_ | _06010_;
	assign _01822_ = _01821_ | _00202_;
	assign _01823_ = _01822_ | ~_01281_;
	assign _01824_ = _01823_ | _01506_;
	assign _01825_ = _01824_ | _01288_;
	assign _01826_ = _01274_ & ~_01825_;
	assign _01827_ = _00202_ | _05346_;
	assign _01828_ = _01827_ | ~_01281_;
	assign _01829_ = _01828_ | ~_01284_;
	assign _01830_ = _01829_ | _01288_;
	assign _01831_ = _01274_ & ~_01830_;
	assign _01832_ = \mchip.design.owner.tokens [6] & ~_01831_;
	assign _01833_ = _01832_ | _01826_;
	assign _01834_ = (_00199_ ? _01820_ : _01833_);
	assign _01835_ = _01525_ | ~_05442_;
	assign _01836_ = _01835_ | ~_01309_;
	assign _01837_ = _01836_ | ~_01311_;
	assign _01838_ = _01837_ | _01523_;
	assign _01839_ = _01838_ | _01318_;
	assign _01840_ = _01303_ & ~_01839_;
	assign _01841_ = _01249_ | ~_01309_;
	assign _01842_ = _01841_ | ~_01311_;
	assign _01843_ = _01842_ | ~_01314_;
	assign _01844_ = _01843_ | _01318_;
	assign _01845_ = _01303_ & ~_01844_;
	assign _01846_ = \mchip.design.owner.tokens [6] & ~_01845_;
	assign _01847_ = _01846_ | _01840_;
	assign _01848_ = (_00131_ ? _01834_ : _01847_);
	assign _01849_ = _01543_ | _05836_;
	assign _01850_ = _01849_ | ~_01339_;
	assign _01851_ = _01850_ | ~_01341_;
	assign _01852_ = _01851_ | _01540_;
	assign _01853_ = _01852_ | _01346_;
	assign _01854_ = _01349_ & ~_01853_;
	assign _01855_ = _05421_ | ~_01339_;
	assign _01856_ = _01855_ | ~_01341_;
	assign _01857_ = _01856_ | _01540_;
	assign _01858_ = _01857_ | _01346_;
	assign _01859_ = _01349_ & ~_01858_;
	assign _01860_ = \mchip.design.owner.tokens [6] & ~_01859_;
	assign _01861_ = _01860_ | _01854_;
	assign _01862_ = (_06005_ ? _01848_ : _01861_);
	assign _01863_ = _01560_ | _01250_;
	assign _01864_ = _01863_ | ~_01372_;
	assign _01865_ = _01864_ | ~_01374_;
	assign _01866_ = _01865_ | ~_01377_;
	assign _01867_ = _01866_ | _01380_;
	assign _01868_ = _01382_ & ~_01867_;
	assign _01869_ = _01723_ | _06012_;
	assign _01870_ = _01869_ | _01250_;
	assign _01871_ = _01870_ | ~_01372_;
	assign _01872_ = _01871_ | ~_01374_;
	assign _01873_ = _01872_ | ~_01377_;
	assign _01874_ = _01873_ | _01380_;
	assign _01875_ = _01382_ & ~_01874_;
	assign _01876_ = \mchip.design.owner.tokens [6] & ~_01875_;
	assign _01877_ = _01876_ | _01868_;
	assign _01878_ = (_05934_ ? _01862_ : _01877_);
	assign _01879_ = _01577_ | _06010_;
	assign _01880_ = _01879_ | _05841_;
	assign _01881_ = _01880_ | ~_01404_;
	assign _01882_ = _01881_ | _01575_;
	assign _01883_ = _01882_ | _01398_;
	assign _01884_ = _01410_ & ~_01883_;
	assign _01885_ = _01584_ | _06010_;
	assign _01886_ = _01885_ | _05841_;
	assign _01887_ = _01886_ | ~_01404_;
	assign _01888_ = _01887_ | _01575_;
	assign _01889_ = _01888_ | _01398_;
	assign _01890_ = _01410_ & ~_01889_;
	assign _01891_ = \mchip.design.owner.tokens [6] & ~_01890_;
	assign _01892_ = _01891_ | _01884_;
	assign _00078_ = (_05827_ ? _01878_ : _01892_);
	assign _01893_ = _01594_ | _01250_;
	assign _01894_ = _01893_ | ~_01252_;
	assign _01895_ = _01894_ | ~_01254_;
	assign _01896_ = _01895_ | _01490_;
	assign _01897_ = _01896_ | _01261_;
	assign _01898_ = _01243_ & ~_01897_;
	assign _01899_ = \mchip.design.owner.tokens [7] & ~_01818_;
	assign _01900_ = _01899_ | _01898_;
	assign _01901_ = _01604_ | _06010_;
	assign _01902_ = _01901_ | _00202_;
	assign _01903_ = _01902_ | ~_01281_;
	assign _01904_ = _01903_ | _01506_;
	assign _01905_ = _01904_ | _01288_;
	assign _01906_ = _01274_ & ~_01905_;
	assign _01907_ = \mchip.design.owner.tokens [7] & ~_01831_;
	assign _01908_ = _01907_ | _01906_;
	assign _01909_ = (_00199_ ? _01900_ : _01908_);
	assign _01910_ = _01615_ | ~_05442_;
	assign _01911_ = _01910_ | ~_01309_;
	assign _01912_ = _01911_ | ~_01311_;
	assign _01913_ = _01912_ | _01523_;
	assign _01914_ = _01913_ | _01318_;
	assign _01915_ = _01303_ & ~_01914_;
	assign _01916_ = \mchip.design.owner.tokens [7] & ~_01845_;
	assign _01917_ = _01916_ | _01915_;
	assign _01918_ = (_00131_ ? _01909_ : _01917_);
	assign _01919_ = _01626_ | _05836_;
	assign _01920_ = _01919_ | ~_01339_;
	assign _01921_ = _01920_ | ~_01341_;
	assign _01922_ = _01921_ | _01540_;
	assign _01923_ = _01922_ | _01346_;
	assign _01924_ = _01349_ & ~_01923_;
	assign _01925_ = \mchip.design.owner.tokens [7] & ~_01859_;
	assign _01926_ = _01925_ | _01924_;
	assign _01927_ = (_06005_ ? _01918_ : _01926_);
	assign _01928_ = _01637_ | _01250_;
	assign _01929_ = _01928_ | ~_01372_;
	assign _01930_ = _01929_ | ~_01374_;
	assign _01931_ = _01930_ | ~_01377_;
	assign _01932_ = _01931_ | _01380_;
	assign _01933_ = _01382_ & ~_01932_;
	assign _01934_ = \mchip.design.owner.tokens [7] & ~_01875_;
	assign _01935_ = _01934_ | _01933_;
	assign _01936_ = (_05934_ ? _01927_ : _01935_);
	assign _01937_ = _01648_ | _06010_;
	assign _01938_ = _01937_ | _05841_;
	assign _01939_ = _01938_ | ~_01404_;
	assign _01940_ = _01939_ | _01575_;
	assign _01941_ = _01940_ | _01398_;
	assign _01942_ = _01410_ & ~_01941_;
	assign _01943_ = \mchip.design.owner.tokens [7] & ~_01890_;
	assign _01944_ = _01943_ | _01942_;
	assign _00089_ = (_05827_ ? _01936_ : _01944_);
	assign _01945_ = _01657_ | _01250_;
	assign _01946_ = _01945_ | ~_01252_;
	assign _01947_ = _01946_ | ~_01254_;
	assign _01948_ = _01947_ | _01490_;
	assign _01949_ = _01948_ | _01261_;
	assign _01950_ = _01243_ & ~_01949_;
	assign _01951_ = _05421_ | ~_00202_;
	assign _01952_ = _01951_ | ~_01254_;
	assign _01953_ = _01952_ | ~_01257_;
	assign _01954_ = _01953_ | _01261_;
	assign _01955_ = _01243_ & ~_01954_;
	assign _01956_ = \mchip.design.owner.tokens [8] & ~_01955_;
	assign _01957_ = _01956_ | _01950_;
	assign _01958_ = _01671_ | _06010_;
	assign _01959_ = _01958_ | _00202_;
	assign _01960_ = _01959_ | ~_01281_;
	assign _01961_ = _01960_ | _01506_;
	assign _01962_ = _01961_ | _01288_;
	assign _01963_ = _01274_ & ~_01962_;
	assign _01964_ = _01309_ | _05431_;
	assign _01965_ = _01964_ | ~_01281_;
	assign _01966_ = _01965_ | ~_01284_;
	assign _01967_ = _01966_ | _01288_;
	assign _01968_ = _01274_ & ~_01967_;
	assign _01969_ = \mchip.design.owner.tokens [8] & ~_01968_;
	assign _01970_ = _01969_ | _01963_;
	assign _01971_ = (_00199_ ? _01957_ : _01970_);
	assign _01972_ = _01686_ | ~_05442_;
	assign _01973_ = _01972_ | ~_01309_;
	assign _01974_ = _01973_ | ~_01311_;
	assign _01975_ = _01974_ | _01523_;
	assign _01976_ = _01975_ | _01318_;
	assign _01977_ = _01303_ & ~_01976_;
	assign _01978_ = _05346_ | ~_04767_;
	assign _01979_ = _01978_ | ~_01311_;
	assign _01980_ = _01979_ | ~_01314_;
	assign _01981_ = _01980_ | _01318_;
	assign _01982_ = _01303_ & ~_01981_;
	assign _01983_ = \mchip.design.owner.tokens [8] & ~_01982_;
	assign _01984_ = _01983_ | _01977_;
	assign _01985_ = (_00131_ ? _01971_ : _01984_);
	assign _01986_ = _01701_ | _05836_;
	assign _01987_ = _01986_ | ~_01339_;
	assign _01988_ = _01987_ | ~_01341_;
	assign _01989_ = _01988_ | _01540_;
	assign _01990_ = _01989_ | _01346_;
	assign _01991_ = _01349_ & ~_01990_;
	assign _01992_ = _01249_ | ~_05945_;
	assign _01993_ = _01992_ | ~_01341_;
	assign _01994_ = _01993_ | _01540_;
	assign _01995_ = _01994_ | _01346_;
	assign _01996_ = _01349_ & ~_01995_;
	assign _01997_ = \mchip.design.owner.tokens [8] & ~_01996_;
	assign _01998_ = _01997_ | _01991_;
	assign _01999_ = (_06005_ ? _01985_ : _01998_);
	assign _02000_ = _01716_ | _01250_;
	assign _02001_ = _02000_ | ~_01372_;
	assign _02002_ = _02001_ | ~_01374_;
	assign _02003_ = _02002_ | ~_01377_;
	assign _02004_ = _02003_ | _01380_;
	assign _02005_ = _01382_ & ~_02004_;
	assign _02006_ = _01724_ | _01250_;
	assign _02007_ = _02006_ | ~_01372_;
	assign _02008_ = _02007_ | ~_01374_;
	assign _02009_ = _02008_ | ~_01377_;
	assign _02010_ = _02009_ | _01380_;
	assign _02011_ = _01382_ & ~_02010_;
	assign _02012_ = \mchip.design.owner.tokens [8] & ~_02011_;
	assign _02013_ = _02012_ | _02005_;
	assign _02014_ = (_05934_ ? _01999_ : _02013_);
	assign _02015_ = _01734_ | _06010_;
	assign _02016_ = _02015_ | _05841_;
	assign _02017_ = _02016_ | ~_01404_;
	assign _02018_ = _02017_ | _01575_;
	assign _02019_ = _02018_ | _01398_;
	assign _02020_ = _01410_ & ~_02019_;
	assign _02021_ = _01741_ | _06010_;
	assign _02022_ = _02021_ | _05841_;
	assign _02023_ = _02022_ | ~_01404_;
	assign _02024_ = _02023_ | _01575_;
	assign _02025_ = _02024_ | _01398_;
	assign _02026_ = _01410_ & ~_02025_;
	assign _02027_ = \mchip.design.owner.tokens [8] & ~_02026_;
	assign _02028_ = _02027_ | _02020_;
	assign _00094_ = (_05827_ ? _02014_ : _02028_);
	assign _02029_ = _01750_ | _01250_;
	assign _02030_ = _02029_ | ~_01252_;
	assign _02031_ = _02030_ | ~_01254_;
	assign _02032_ = _02031_ | _01490_;
	assign _02033_ = _02032_ | _01261_;
	assign _02034_ = _01243_ & ~_02033_;
	assign _02035_ = \mchip.design.owner.tokens [9] & ~_01955_;
	assign _02036_ = _02035_ | _02034_;
	assign _02037_ = _01759_ | _06010_;
	assign _02038_ = _02037_ | _00202_;
	assign _02039_ = _02038_ | ~_01281_;
	assign _02040_ = _02039_ | _01506_;
	assign _02041_ = _02040_ | _01288_;
	assign _02042_ = _01274_ & ~_02041_;
	assign _02043_ = \mchip.design.owner.tokens [9] & ~_01968_;
	assign _02044_ = _02043_ | _02042_;
	assign _02045_ = (_00199_ ? _02036_ : _02044_);
	assign _02046_ = _01769_ | ~_05442_;
	assign _02047_ = _02046_ | ~_01309_;
	assign _02048_ = _02047_ | ~_01311_;
	assign _02049_ = _02048_ | _01523_;
	assign _02050_ = _02049_ | _01318_;
	assign _02051_ = _01303_ & ~_02050_;
	assign _02052_ = \mchip.design.owner.tokens [9] & ~_01982_;
	assign _02053_ = _02052_ | _02051_;
	assign _02054_ = (_00131_ ? _02045_ : _02053_);
	assign _02055_ = _01779_ | _05836_;
	assign _02056_ = _02055_ | ~_01339_;
	assign _02057_ = _02056_ | ~_01341_;
	assign _02058_ = _02057_ | _01540_;
	assign _02059_ = _02058_ | _01346_;
	assign _02060_ = _01349_ & ~_02059_;
	assign _02061_ = \mchip.design.owner.tokens [9] & ~_01996_;
	assign _02062_ = _02061_ | _02060_;
	assign _02063_ = (_06005_ ? _02054_ : _02062_);
	assign _02064_ = _01789_ | _01250_;
	assign _02065_ = _02064_ | ~_01372_;
	assign _02066_ = _02065_ | ~_01374_;
	assign _02067_ = _02066_ | ~_01377_;
	assign _02068_ = _02067_ | _01380_;
	assign _02069_ = _01382_ & ~_02068_;
	assign _02070_ = \mchip.design.owner.tokens [9] & ~_02011_;
	assign _02071_ = _02070_ | _02069_;
	assign _02072_ = (_05934_ ? _02063_ : _02071_);
	assign _02073_ = _01799_ | _06010_;
	assign _02074_ = _02073_ | _05841_;
	assign _02075_ = _02074_ | ~_01404_;
	assign _02076_ = _02075_ | _01575_;
	assign _02077_ = _02076_ | _01398_;
	assign _02078_ = _01410_ & ~_02077_;
	assign _02079_ = \mchip.design.owner.tokens [9] & ~_02026_;
	assign _02080_ = _02079_ | _02078_;
	assign _00095_ = (_05827_ ? _02072_ : _02080_);
	assign _02081_ = _01493_ | _01252_;
	assign _02082_ = _02081_ | ~_01254_;
	assign _02083_ = _02082_ | _01490_;
	assign _02084_ = _02083_ | _01261_;
	assign _02085_ = _01243_ & ~_02084_;
	assign _02086_ = _01252_ | _01249_;
	assign _02087_ = _02086_ | ~_01254_;
	assign _02088_ = _02087_ | ~_01257_;
	assign _02089_ = _02088_ | _01261_;
	assign _02090_ = _01243_ & ~_02089_;
	assign _02091_ = \mchip.design.owner.tokens [10] & ~_02090_;
	assign _02092_ = _02091_ | _02085_;
	assign _02093_ = _01509_ | ~_00202_;
	assign _02094_ = _02093_ | ~_01281_;
	assign _02095_ = _02094_ | _01506_;
	assign _02096_ = _02095_ | _01288_;
	assign _02097_ = _01274_ & ~_02096_;
	assign _02098_ = _01951_ | ~_01281_;
	assign _02099_ = _02098_ | ~_01284_;
	assign _02100_ = _02099_ | _01288_;
	assign _02101_ = _01274_ & ~_02100_;
	assign _02102_ = \mchip.design.owner.tokens [10] & ~_02101_;
	assign _02103_ = _02102_ | _02097_;
	assign _02104_ = (_00199_ ? _02092_ : _02103_);
	assign _02105_ = _01526_ | _01309_;
	assign _02106_ = _02105_ | ~_01311_;
	assign _02107_ = _02106_ | _01523_;
	assign _02108_ = _02107_ | _01318_;
	assign _02109_ = _01303_ & ~_02108_;
	assign _02110_ = _01964_ | ~_01311_;
	assign _02111_ = _02110_ | ~_01314_;
	assign _02112_ = _02111_ | _01318_;
	assign _02113_ = _01303_ & ~_02112_;
	assign _02114_ = \mchip.design.owner.tokens [10] & ~_02113_;
	assign _02115_ = _02114_ | _02109_;
	assign _02116_ = (_00131_ ? _02104_ : _02115_);
	assign _02117_ = _01544_ | _01339_;
	assign _02118_ = _02117_ | ~_01341_;
	assign _02119_ = _02118_ | _01540_;
	assign _02120_ = _02119_ | _01346_;
	assign _02121_ = _01349_ & ~_02120_;
	assign _02122_ = _01339_ | _05346_;
	assign _02123_ = _02122_ | ~_01341_;
	assign _02124_ = _02123_ | _01540_;
	assign _02125_ = _02124_ | _01346_;
	assign _02126_ = _01349_ & ~_02125_;
	assign _02127_ = \mchip.design.owner.tokens [10] & ~_02126_;
	assign _02128_ = _02127_ | _02121_;
	assign _02129_ = (_06005_ ? _02116_ : _02128_);
	assign _02130_ = _01561_ | _01372_;
	assign _02131_ = _02130_ | ~_01374_;
	assign _02132_ = _02131_ | ~_01377_;
	assign _02133_ = _02132_ | _01380_;
	assign _02134_ = _01382_ & ~_02133_;
	assign _02135_ = _01372_ | _01249_;
	assign _02136_ = _02135_ | ~_01374_;
	assign _02137_ = _02136_ | ~_01377_;
	assign _02138_ = _02137_ | _01380_;
	assign _02139_ = _01382_ & ~_02138_;
	assign _02140_ = \mchip.design.owner.tokens [10] & ~_02139_;
	assign _02141_ = _02140_ | _02134_;
	assign _02142_ = (_05934_ ? _02129_ : _02141_);
	assign _02143_ = _01578_ | ~_05841_;
	assign _02144_ = _02143_ | ~_01404_;
	assign _02145_ = _02144_ | _01575_;
	assign _02146_ = _02145_ | _01398_;
	assign _02147_ = _01410_ & ~_02146_;
	assign _02148_ = _01585_ | ~_05841_;
	assign _02149_ = _02148_ | ~_01404_;
	assign _02150_ = _02149_ | _01575_;
	assign _02151_ = _02150_ | _01398_;
	assign _02152_ = _01410_ & ~_02151_;
	assign _02153_ = \mchip.design.owner.tokens [10] & ~_02152_;
	assign _02154_ = _02153_ | _02147_;
	assign _00013_ = (_05827_ ? _02142_ : _02154_);
	assign _02155_ = _01595_ | _01252_;
	assign _02156_ = _02155_ | ~_01254_;
	assign _02157_ = _02156_ | _01490_;
	assign _02158_ = _02157_ | _01261_;
	assign _02159_ = _01243_ & ~_02158_;
	assign _02160_ = \mchip.design.owner.tokens [11] & ~_02090_;
	assign _02161_ = _02160_ | _02159_;
	assign _02162_ = _01605_ | ~_00202_;
	assign _02163_ = _02162_ | ~_01281_;
	assign _02164_ = _02163_ | _01506_;
	assign _02165_ = _02164_ | _01288_;
	assign _02166_ = _01274_ & ~_02165_;
	assign _02167_ = \mchip.design.owner.tokens [11] & ~_02101_;
	assign _02168_ = _02167_ | _02166_;
	assign _02169_ = (_00199_ ? _02161_ : _02168_);
	assign _02170_ = _01616_ | _01309_;
	assign _02171_ = _02170_ | ~_01311_;
	assign _02172_ = _02171_ | _01523_;
	assign _02173_ = _02172_ | _01318_;
	assign _02174_ = _01303_ & ~_02173_;
	assign _02175_ = \mchip.design.owner.tokens [11] & ~_02113_;
	assign _02176_ = _02175_ | _02174_;
	assign _02177_ = (_00131_ ? _02169_ : _02176_);
	assign _02178_ = _01627_ | _01339_;
	assign _02179_ = _02178_ | ~_01341_;
	assign _02180_ = _02179_ | _01540_;
	assign _02181_ = _02180_ | _01346_;
	assign _02182_ = _01349_ & ~_02181_;
	assign _02183_ = \mchip.design.owner.tokens [11] & ~_02126_;
	assign _02184_ = _02183_ | _02182_;
	assign _02185_ = (_06005_ ? _02177_ : _02184_);
	assign _02186_ = _01638_ | _01372_;
	assign _02187_ = _02186_ | ~_01374_;
	assign _02188_ = _02187_ | ~_01377_;
	assign _02189_ = _02188_ | _01380_;
	assign _02190_ = _01382_ & ~_02189_;
	assign _02191_ = \mchip.design.owner.tokens [11] & ~_02139_;
	assign _02192_ = _02191_ | _02190_;
	assign _02193_ = (_05934_ ? _02185_ : _02192_);
	assign _02194_ = _01649_ | ~_05841_;
	assign _02195_ = _02194_ | ~_01404_;
	assign _02196_ = _02195_ | _01575_;
	assign _02197_ = _02196_ | _01398_;
	assign _02198_ = _01410_ & ~_02197_;
	assign _02199_ = \mchip.design.owner.tokens [11] & ~_02152_;
	assign _02200_ = _02199_ | _02198_;
	assign _00014_ = (_05827_ ? _02193_ : _02200_);
	assign _02201_ = _01658_ | _01252_;
	assign _02202_ = _02201_ | ~_01254_;
	assign _02203_ = _02202_ | _01490_;
	assign _02204_ = _02203_ | _01261_;
	assign _02205_ = _01243_ & ~_02204_;
	assign _02206_ = _01252_ | _05346_;
	assign _02207_ = _02206_ | ~_01254_;
	assign _02208_ = _02207_ | ~_01257_;
	assign _02209_ = _02208_ | _01261_;
	assign _02210_ = _01243_ & ~_02209_;
	assign _02211_ = \mchip.design.owner.tokens [12] & ~_02210_;
	assign _02212_ = _02211_ | _02205_;
	assign _02213_ = _01672_ | ~_00202_;
	assign _02214_ = _02213_ | ~_01281_;
	assign _02215_ = _02214_ | _01506_;
	assign _02216_ = _02215_ | _01288_;
	assign _02217_ = _01274_ & ~_02216_;
	assign _02218_ = _01249_ | ~_00202_;
	assign _02219_ = _02218_ | ~_01281_;
	assign _02220_ = _02219_ | ~_01284_;
	assign _02221_ = _02220_ | _01288_;
	assign _02222_ = _01274_ & ~_02221_;
	assign _02223_ = \mchip.design.owner.tokens [12] & ~_02222_;
	assign _02224_ = _02223_ | _02217_;
	assign _02225_ = (_00199_ ? _02212_ : _02224_);
	assign _02226_ = _01687_ | _01309_;
	assign _02227_ = _02226_ | ~_01311_;
	assign _02228_ = _02227_ | _01523_;
	assign _02229_ = _02228_ | _01318_;
	assign _02230_ = _01303_ & ~_02229_;
	assign _02231_ = _01309_ | _05421_;
	assign _02232_ = _02231_ | ~_01311_;
	assign _02233_ = _02232_ | ~_01314_;
	assign _02234_ = _02233_ | _01318_;
	assign _02235_ = _01303_ & ~_02234_;
	assign _02236_ = \mchip.design.owner.tokens [12] & ~_02235_;
	assign _02237_ = _02236_ | _02230_;
	assign _02238_ = (_00131_ ? _02225_ : _02237_);
	assign _02239_ = _01702_ | _01339_;
	assign _02240_ = _02239_ | ~_01341_;
	assign _02241_ = _02240_ | _01540_;
	assign _02242_ = _02241_ | _01346_;
	assign _02243_ = _01349_ & ~_02242_;
	assign _02244_ = _01339_ | _05431_;
	assign _02245_ = _02244_ | ~_01341_;
	assign _02246_ = _02245_ | _01540_;
	assign _02247_ = _02246_ | _01346_;
	assign _02248_ = _01349_ & ~_02247_;
	assign _02249_ = \mchip.design.owner.tokens [12] & ~_02248_;
	assign _02250_ = _02249_ | _02243_;
	assign _02251_ = (_06005_ ? _02238_ : _02250_);
	assign _02252_ = _01717_ | _01372_;
	assign _02253_ = _02252_ | ~_01374_;
	assign _02254_ = _02253_ | ~_01377_;
	assign _02255_ = _02254_ | _01380_;
	assign _02256_ = _01382_ & ~_02255_;
	assign _02257_ = _01725_ | _01372_;
	assign _02258_ = _02257_ | ~_01374_;
	assign _02259_ = _02258_ | ~_01377_;
	assign _02260_ = _02259_ | _01380_;
	assign _02261_ = _01382_ & ~_02260_;
	assign _02262_ = \mchip.design.owner.tokens [12] & ~_02261_;
	assign _02263_ = _02262_ | _02256_;
	assign _02264_ = (_05934_ ? _02251_ : _02263_);
	assign _02265_ = _01735_ | ~_05841_;
	assign _02266_ = _02265_ | ~_01404_;
	assign _02267_ = _02266_ | _01575_;
	assign _02268_ = _02267_ | _01398_;
	assign _02269_ = _01410_ & ~_02268_;
	assign _02270_ = _01742_ | ~_05841_;
	assign _02271_ = _02270_ | ~_01404_;
	assign _02272_ = _02271_ | _01575_;
	assign _02273_ = _02272_ | _01398_;
	assign _02274_ = _01410_ & ~_02273_;
	assign _02275_ = \mchip.design.owner.tokens [12] & ~_02274_;
	assign _02276_ = _02275_ | _02269_;
	assign _00015_ = (_05827_ ? _02264_ : _02276_);
	assign _02277_ = _01751_ | _01252_;
	assign _02278_ = _02277_ | ~_01254_;
	assign _02279_ = _02278_ | _01490_;
	assign _02280_ = _02279_ | _01261_;
	assign _02281_ = _01243_ & ~_02280_;
	assign _02282_ = \mchip.design.owner.tokens [13] & ~_02210_;
	assign _02283_ = _02282_ | _02281_;
	assign _02284_ = _01760_ | ~_00202_;
	assign _02285_ = _02284_ | ~_01281_;
	assign _02286_ = _02285_ | _01506_;
	assign _02287_ = _02286_ | _01288_;
	assign _02288_ = _01274_ & ~_02287_;
	assign _02289_ = \mchip.design.owner.tokens [13] & ~_02222_;
	assign _02290_ = _02289_ | _02288_;
	assign _02291_ = (_00199_ ? _02283_ : _02290_);
	assign _02292_ = _01770_ | _01309_;
	assign _02293_ = _02292_ | ~_01311_;
	assign _02294_ = _02293_ | _01523_;
	assign _02295_ = _02294_ | _01318_;
	assign _02296_ = _01303_ & ~_02295_;
	assign _02297_ = \mchip.design.owner.tokens [13] & ~_02235_;
	assign _02298_ = _02297_ | _02296_;
	assign _02299_ = (_00131_ ? _02291_ : _02298_);
	assign _02300_ = _01780_ | _01339_;
	assign _02301_ = _02300_ | ~_01341_;
	assign _02302_ = _02301_ | _01540_;
	assign _02303_ = _02302_ | _01346_;
	assign _02304_ = _01349_ & ~_02303_;
	assign _02305_ = \mchip.design.owner.tokens [13] & ~_02248_;
	assign _02306_ = _02305_ | _02304_;
	assign _02307_ = (_06005_ ? _02299_ : _02306_);
	assign _02308_ = _01790_ | _01372_;
	assign _02309_ = _02308_ | ~_01374_;
	assign _02310_ = _02309_ | ~_01377_;
	assign _02311_ = _02310_ | _01380_;
	assign _02312_ = _01382_ & ~_02311_;
	assign _02313_ = \mchip.design.owner.tokens [13] & ~_02261_;
	assign _02314_ = _02313_ | _02312_;
	assign _02315_ = (_05934_ ? _02307_ : _02314_);
	assign _02316_ = _01800_ | ~_05841_;
	assign _02317_ = _02316_ | ~_01404_;
	assign _02318_ = _02317_ | _01575_;
	assign _02319_ = _02318_ | _01398_;
	assign _02320_ = _01410_ & ~_02319_;
	assign _02321_ = \mchip.design.owner.tokens [13] & ~_02274_;
	assign _02322_ = _02321_ | _02320_;
	assign _00016_ = (_05827_ ? _02315_ : _02322_);
	assign _02323_ = _01808_ | _01252_;
	assign _02324_ = _02323_ | ~_01254_;
	assign _02325_ = _02324_ | _01490_;
	assign _02326_ = _02325_ | _01261_;
	assign _02327_ = _01243_ & ~_02326_;
	assign _02328_ = _01252_ | _05431_;
	assign _02329_ = _02328_ | ~_01254_;
	assign _02330_ = _02329_ | ~_01257_;
	assign _02331_ = _02330_ | _01261_;
	assign _02332_ = _01243_ & ~_02331_;
	assign _02333_ = \mchip.design.owner.tokens [14] & ~_02332_;
	assign _02334_ = _02333_ | _02327_;
	assign _02335_ = _01821_ | ~_00202_;
	assign _02336_ = _02335_ | ~_01281_;
	assign _02337_ = _02336_ | _01506_;
	assign _02338_ = _02337_ | _01288_;
	assign _02339_ = _01274_ & ~_02338_;
	assign _02340_ = _05346_ | ~_00202_;
	assign _02341_ = _02340_ | ~_01281_;
	assign _02342_ = _02341_ | ~_01284_;
	assign _02343_ = _02342_ | _01288_;
	assign _02344_ = _01274_ & ~_02343_;
	assign _02345_ = \mchip.design.owner.tokens [14] & ~_02344_;
	assign _02346_ = _02345_ | _02339_;
	assign _02347_ = (_00199_ ? _02334_ : _02346_);
	assign _02348_ = _01835_ | _01309_;
	assign _02349_ = _02348_ | ~_01311_;
	assign _02350_ = _02349_ | _01523_;
	assign _02351_ = _02350_ | _01318_;
	assign _02352_ = _01303_ & ~_02351_;
	assign _02353_ = _01309_ | _01249_;
	assign _02354_ = _02353_ | ~_01311_;
	assign _02355_ = _02354_ | ~_01314_;
	assign _02356_ = _02355_ | _01318_;
	assign _02357_ = _01303_ & ~_02356_;
	assign _02358_ = \mchip.design.owner.tokens [14] & ~_02357_;
	assign _02359_ = _02358_ | _02352_;
	assign _02360_ = (_00131_ ? _02347_ : _02359_);
	assign _02361_ = _01849_ | _01339_;
	assign _02362_ = _02361_ | ~_01341_;
	assign _02363_ = _02362_ | _01540_;
	assign _02364_ = _02363_ | _01346_;
	assign _02365_ = _01349_ & ~_02364_;
	assign _02366_ = _01339_ | _05421_;
	assign _02367_ = _02366_ | ~_01341_;
	assign _02368_ = _02367_ | _01540_;
	assign _02369_ = _02368_ | _01346_;
	assign _02370_ = _01349_ & ~_02369_;
	assign _02371_ = \mchip.design.owner.tokens [14] & ~_02370_;
	assign _02372_ = _02371_ | _02365_;
	assign _02373_ = (_06005_ ? _02360_ : _02372_);
	assign _02374_ = _01863_ | _01372_;
	assign _02375_ = _02374_ | ~_01374_;
	assign _02376_ = _02375_ | ~_01377_;
	assign _02377_ = _02376_ | _01380_;
	assign _02378_ = _01382_ & ~_02377_;
	assign _02379_ = _01870_ | _01372_;
	assign _02380_ = _02379_ | ~_01374_;
	assign _02381_ = _02380_ | ~_01377_;
	assign _02382_ = _02381_ | _01380_;
	assign _02383_ = _01382_ & ~_02382_;
	assign _02384_ = \mchip.design.owner.tokens [14] & ~_02383_;
	assign _02385_ = _02384_ | _02378_;
	assign _02386_ = (_05934_ ? _02373_ : _02385_);
	assign _02387_ = _01879_ | ~_05841_;
	assign _02388_ = _02387_ | ~_01404_;
	assign _02389_ = _02388_ | _01575_;
	assign _02390_ = _02389_ | _01398_;
	assign _02391_ = _01410_ & ~_02390_;
	assign _02392_ = _01885_ | ~_05841_;
	assign _02393_ = _02392_ | ~_01404_;
	assign _02394_ = _02393_ | _01575_;
	assign _02395_ = _02394_ | _01398_;
	assign _02396_ = _01410_ & ~_02395_;
	assign _02397_ = \mchip.design.owner.tokens [14] & ~_02396_;
	assign _02398_ = _02397_ | _02391_;
	assign _00017_ = (_05827_ ? _02386_ : _02398_);
	assign _02399_ = _01893_ | _01252_;
	assign _02400_ = _02399_ | ~_01254_;
	assign _02401_ = _02400_ | _01490_;
	assign _02402_ = _02401_ | _01261_;
	assign _02403_ = _01243_ & ~_02402_;
	assign _02404_ = \mchip.design.owner.tokens [15] & ~_02332_;
	assign _02405_ = _02404_ | _02403_;
	assign _02406_ = _01901_ | ~_00202_;
	assign _02407_ = _02406_ | ~_01281_;
	assign _02408_ = _02407_ | _01506_;
	assign _02409_ = _02408_ | _01288_;
	assign _02410_ = _01274_ & ~_02409_;
	assign _02411_ = \mchip.design.owner.tokens [15] & ~_02344_;
	assign _02412_ = _02411_ | _02410_;
	assign _02413_ = (_00199_ ? _02405_ : _02412_);
	assign _02414_ = _01910_ | _01309_;
	assign _02415_ = _02414_ | ~_01311_;
	assign _02416_ = _02415_ | _01523_;
	assign _02417_ = _02416_ | _01318_;
	assign _02418_ = _01303_ & ~_02417_;
	assign _02419_ = \mchip.design.owner.tokens [15] & ~_02357_;
	assign _02420_ = _02419_ | _02418_;
	assign _02421_ = (_00131_ ? _02413_ : _02420_);
	assign _02422_ = _01919_ | _01339_;
	assign _02423_ = _02422_ | ~_01341_;
	assign _02424_ = _02423_ | _01540_;
	assign _02425_ = _02424_ | _01346_;
	assign _02426_ = _01349_ & ~_02425_;
	assign _02427_ = \mchip.design.owner.tokens [15] & ~_02370_;
	assign _02428_ = _02427_ | _02426_;
	assign _02429_ = (_06005_ ? _02421_ : _02428_);
	assign _02430_ = _01928_ | _01372_;
	assign _02431_ = _02430_ | ~_01374_;
	assign _02432_ = _02431_ | ~_01377_;
	assign _02433_ = _02432_ | _01380_;
	assign _02434_ = _01382_ & ~_02433_;
	assign _02435_ = \mchip.design.owner.tokens [15] & ~_02383_;
	assign _02436_ = _02435_ | _02434_;
	assign _02437_ = (_05934_ ? _02429_ : _02436_);
	assign _02438_ = _01937_ | ~_05841_;
	assign _02439_ = _02438_ | ~_01404_;
	assign _02440_ = _02439_ | _01575_;
	assign _02441_ = _02440_ | _01398_;
	assign _02442_ = _01410_ & ~_02441_;
	assign _02443_ = \mchip.design.owner.tokens [15] & ~_02396_;
	assign _02444_ = _02443_ | _02442_;
	assign _00018_ = (_05827_ ? _02437_ : _02444_);
	assign _02445_ = _01945_ | _01252_;
	assign _02446_ = _02445_ | ~_01254_;
	assign _02447_ = _02446_ | _01490_;
	assign _02448_ = _02447_ | _01261_;
	assign _02449_ = _01243_ & ~_02448_;
	assign _02450_ = _01515_ | ~_01254_;
	assign _02451_ = _02450_ | ~_01257_;
	assign _02452_ = _02451_ | _01261_;
	assign _02453_ = _01243_ & ~_02452_;
	assign _02454_ = \mchip.design.owner.tokens [16] & ~_02453_;
	assign _02455_ = _02454_ | _02449_;
	assign _02456_ = _01958_ | ~_00202_;
	assign _02457_ = _02456_ | ~_01281_;
	assign _02458_ = _02457_ | _01506_;
	assign _02459_ = _02458_ | _01288_;
	assign _02460_ = _01274_ & ~_02459_;
	assign _02461_ = _01532_ | ~_01281_;
	assign _02462_ = _02461_ | ~_01284_;
	assign _02463_ = _02462_ | _01288_;
	assign _02464_ = _01274_ & ~_02463_;
	assign _02465_ = \mchip.design.owner.tokens [16] & ~_02464_;
	assign _02466_ = _02465_ | _02460_;
	assign _02467_ = (_00199_ ? _02455_ : _02466_);
	assign _02468_ = _01972_ | _01309_;
	assign _02469_ = _02468_ | ~_01311_;
	assign _02470_ = _02469_ | _01523_;
	assign _02471_ = _02470_ | _01318_;
	assign _02472_ = _01303_ & ~_02471_;
	assign _02473_ = _04767_ | _05346_;
	assign _02474_ = _02473_ | ~_01311_;
	assign _02475_ = _02474_ | ~_01314_;
	assign _02476_ = _02475_ | _01318_;
	assign _02477_ = _01303_ & ~_02476_;
	assign _02478_ = \mchip.design.owner.tokens [16] & ~_02477_;
	assign _02479_ = _02478_ | _02472_;
	assign _02480_ = (_00131_ ? _02467_ : _02479_);
	assign _02481_ = _01986_ | _01339_;
	assign _02482_ = _02481_ | ~_01341_;
	assign _02483_ = _02482_ | _01540_;
	assign _02484_ = _02483_ | _01346_;
	assign _02485_ = _01349_ & ~_02484_;
	assign _02486_ = _01249_ | _05945_;
	assign _02487_ = _02486_ | ~_01341_;
	assign _02488_ = _02487_ | _01540_;
	assign _02489_ = _02488_ | _01346_;
	assign _02490_ = _01349_ & ~_02489_;
	assign _02491_ = \mchip.design.owner.tokens [16] & ~_02490_;
	assign _02492_ = _02491_ | _02485_;
	assign _02493_ = (_06005_ ? _02480_ : _02492_);
	assign _02494_ = _02000_ | _01372_;
	assign _02495_ = _02494_ | ~_01374_;
	assign _02496_ = _02495_ | ~_01377_;
	assign _02497_ = _02496_ | _01380_;
	assign _02498_ = _01382_ & ~_02497_;
	assign _02499_ = _02006_ | _01372_;
	assign _02500_ = _02499_ | ~_01374_;
	assign _02501_ = _02500_ | ~_01377_;
	assign _02502_ = _02501_ | _01380_;
	assign _02503_ = _01382_ & ~_02502_;
	assign _02504_ = \mchip.design.owner.tokens [16] & ~_02503_;
	assign _02505_ = _02504_ | _02498_;
	assign _02506_ = (_05934_ ? _02493_ : _02505_);
	assign _02507_ = _02015_ | ~_05841_;
	assign _02508_ = _02507_ | ~_01404_;
	assign _02509_ = _02508_ | _01575_;
	assign _02510_ = _02509_ | _01398_;
	assign _02511_ = _01410_ & ~_02510_;
	assign _02512_ = _02021_ | ~_05841_;
	assign _02513_ = _02512_ | ~_01404_;
	assign _02514_ = _02513_ | _01575_;
	assign _02515_ = _02514_ | _01398_;
	assign _02516_ = _01410_ & ~_02515_;
	assign _02517_ = \mchip.design.owner.tokens [16] & ~_02516_;
	assign _02518_ = _02517_ | _02511_;
	assign _00019_ = (_05827_ ? _02506_ : _02518_);
	assign _02519_ = _02029_ | _01252_;
	assign _02520_ = _02519_ | ~_01254_;
	assign _02521_ = _02520_ | _01490_;
	assign _02522_ = _02521_ | _01261_;
	assign _02523_ = _01243_ & ~_02522_;
	assign _02524_ = \mchip.design.owner.tokens [17] & ~_02453_;
	assign _02525_ = _02524_ | _02523_;
	assign _02526_ = _02037_ | ~_00202_;
	assign _02527_ = _02526_ | ~_01281_;
	assign _02528_ = _02527_ | _01506_;
	assign _02529_ = _02528_ | _01288_;
	assign _02530_ = _01274_ & ~_02529_;
	assign _02531_ = \mchip.design.owner.tokens [17] & ~_02464_;
	assign _02532_ = _02531_ | _02530_;
	assign _02533_ = (_00199_ ? _02525_ : _02532_);
	assign _02534_ = _02046_ | _01309_;
	assign _02535_ = _02534_ | ~_01311_;
	assign _02536_ = _02535_ | _01523_;
	assign _02537_ = _02536_ | _01318_;
	assign _02538_ = _01303_ & ~_02537_;
	assign _02539_ = \mchip.design.owner.tokens [17] & ~_02477_;
	assign _02540_ = _02539_ | _02538_;
	assign _02541_ = (_00131_ ? _02533_ : _02540_);
	assign _02542_ = _02055_ | _01339_;
	assign _02543_ = _02542_ | ~_01341_;
	assign _02544_ = _02543_ | _01540_;
	assign _02545_ = _02544_ | _01346_;
	assign _02546_ = _01349_ & ~_02545_;
	assign _02547_ = \mchip.design.owner.tokens [17] & ~_02490_;
	assign _02548_ = _02547_ | _02546_;
	assign _02549_ = (_06005_ ? _02541_ : _02548_);
	assign _02550_ = _02064_ | _01372_;
	assign _02551_ = _02550_ | ~_01374_;
	assign _02552_ = _02551_ | ~_01377_;
	assign _02553_ = _02552_ | _01380_;
	assign _02554_ = _01382_ & ~_02553_;
	assign _02555_ = \mchip.design.owner.tokens [17] & ~_02503_;
	assign _02556_ = _02555_ | _02554_;
	assign _02557_ = (_05934_ ? _02549_ : _02556_);
	assign _02558_ = _02073_ | ~_05841_;
	assign _02559_ = _02558_ | ~_01404_;
	assign _02560_ = _02559_ | _01575_;
	assign _02561_ = _02560_ | _01398_;
	assign _02562_ = _01410_ & ~_02561_;
	assign _02563_ = \mchip.design.owner.tokens [17] & ~_02516_;
	assign _02564_ = _02563_ | _02562_;
	assign _00020_ = (_05827_ ? _02557_ : _02564_);
	assign _02565_ = _01494_ | _01254_;
	assign _02566_ = _02565_ | _01490_;
	assign _02567_ = _02566_ | _01261_;
	assign _02568_ = _01243_ & ~_02567_;
	assign _02569_ = _01499_ | _01254_;
	assign _02570_ = _02569_ | ~_01257_;
	assign _02571_ = _02570_ | _01261_;
	assign _02572_ = _01243_ & ~_02571_;
	assign _02573_ = \mchip.design.owner.tokens [18] & ~_02572_;
	assign _02574_ = _02573_ | _02568_;
	assign _02575_ = _01510_ | _01281_;
	assign _02576_ = _02575_ | _01506_;
	assign _02577_ = _02576_ | _01288_;
	assign _02578_ = _01274_ & ~_02577_;
	assign _02579_ = _01515_ | _01281_;
	assign _02580_ = _02579_ | ~_01284_;
	assign _02581_ = _02580_ | _01288_;
	assign _02582_ = _01274_ & ~_02581_;
	assign _02583_ = \mchip.design.owner.tokens [18] & ~_02582_;
	assign _02584_ = _02583_ | _02578_;
	assign _02585_ = (_00199_ ? _02574_ : _02584_);
	assign _02586_ = _01527_ | _01311_;
	assign _02587_ = _02586_ | _01523_;
	assign _02588_ = _02587_ | _01318_;
	assign _02589_ = _01303_ & ~_02588_;
	assign _02590_ = _01532_ | _01311_;
	assign _02591_ = _02590_ | ~_01314_;
	assign _02592_ = _02591_ | _01318_;
	assign _02593_ = _01303_ & ~_02592_;
	assign _02594_ = \mchip.design.owner.tokens [18] & ~_02593_;
	assign _02595_ = _02594_ | _02589_;
	assign _02596_ = (_00131_ ? _02585_ : _02595_);
	assign _02597_ = _01545_ | _01341_;
	assign _02598_ = _02597_ | _01540_;
	assign _02599_ = _02598_ | _01346_;
	assign _02600_ = _01349_ & ~_02599_;
	assign _02601_ = _01550_ | _01341_;
	assign _02602_ = _02601_ | _01540_;
	assign _02603_ = _02602_ | _01346_;
	assign _02604_ = _01349_ & ~_02603_;
	assign _02605_ = \mchip.design.owner.tokens [18] & ~_02604_;
	assign _02606_ = _02605_ | _02600_;
	assign _02607_ = (_06005_ ? _02596_ : _02606_);
	assign _02608_ = _01562_ | _01374_;
	assign _02609_ = _02608_ | ~_01377_;
	assign _02610_ = _02609_ | _01380_;
	assign _02611_ = _01382_ & ~_02610_;
	assign _02612_ = _01567_ | _01374_;
	assign _02613_ = _02612_ | ~_01377_;
	assign _02614_ = _02613_ | _01380_;
	assign _02615_ = _01382_ & ~_02614_;
	assign _02616_ = \mchip.design.owner.tokens [18] & ~_02615_;
	assign _02617_ = _02616_ | _02611_;
	assign _02618_ = (_05934_ ? _02607_ : _02617_);
	assign _02619_ = _01579_ | _01404_;
	assign _02620_ = _02619_ | _01575_;
	assign _02621_ = _02620_ | _01398_;
	assign _02622_ = _01410_ & ~_02621_;
	assign _02623_ = _01586_ | _01404_;
	assign _02624_ = _02623_ | _01575_;
	assign _02625_ = _02624_ | _01398_;
	assign _02626_ = _01410_ & ~_02625_;
	assign _02627_ = \mchip.design.owner.tokens [18] & ~_02626_;
	assign _02628_ = _02627_ | _02622_;
	assign _00021_ = (_05827_ ? _02618_ : _02628_);
	assign _02629_ = _01596_ | _01254_;
	assign _02630_ = _02629_ | _01490_;
	assign _02631_ = _02630_ | _01261_;
	assign _02632_ = _01243_ & ~_02631_;
	assign _02633_ = \mchip.design.owner.tokens [19] & ~_02572_;
	assign _02634_ = _02633_ | _02632_;
	assign _02635_ = _01606_ | _01281_;
	assign _02636_ = _02635_ | _01506_;
	assign _02637_ = _02636_ | _01288_;
	assign _02638_ = _01274_ & ~_02637_;
	assign _02639_ = \mchip.design.owner.tokens [19] & ~_02582_;
	assign _02640_ = _02639_ | _02638_;
	assign _02641_ = (_00199_ ? _02634_ : _02640_);
	assign _02642_ = _01617_ | _01311_;
	assign _02643_ = _02642_ | _01523_;
	assign _02644_ = _02643_ | _01318_;
	assign _02645_ = _01303_ & ~_02644_;
	assign _02646_ = \mchip.design.owner.tokens [19] & ~_02593_;
	assign _02647_ = _02646_ | _02645_;
	assign _02648_ = (_00131_ ? _02641_ : _02647_);
	assign _02649_ = _01628_ | _01341_;
	assign _02650_ = _02649_ | _01540_;
	assign _02651_ = _02650_ | _01346_;
	assign _02652_ = _01349_ & ~_02651_;
	assign _02653_ = \mchip.design.owner.tokens [19] & ~_02604_;
	assign _02654_ = _02653_ | _02652_;
	assign _02655_ = (_06005_ ? _02648_ : _02654_);
	assign _02656_ = _01639_ | _01374_;
	assign _02657_ = _02656_ | ~_01377_;
	assign _02658_ = _02657_ | _01380_;
	assign _02659_ = _01382_ & ~_02658_;
	assign _02660_ = \mchip.design.owner.tokens [19] & ~_02615_;
	assign _02662_ = _02660_ | _02659_;
	assign _02663_ = (_05934_ ? _02655_ : _02662_);
	assign _02664_ = _01650_ | _01404_;
	assign _02665_ = _02664_ | _01575_;
	assign _02666_ = _02665_ | _01398_;
	assign _02667_ = _01410_ & ~_02666_;
	assign _02668_ = \mchip.design.owner.tokens [19] & ~_02626_;
	assign _02669_ = _02668_ | _02667_;
	assign _00022_ = (_05827_ ? _02663_ : _02669_);
	assign _02670_ = _01659_ | _01254_;
	assign _02672_ = _02670_ | _01490_;
	assign _02673_ = _02672_ | _01261_;
	assign _02674_ = _01243_ & ~_02673_;
	assign _02675_ = _01664_ | _01254_;
	assign _02676_ = _02675_ | ~_01257_;
	assign _02677_ = _02676_ | _01261_;
	assign _02678_ = _01243_ & ~_02677_;
	assign _02679_ = \mchip.design.owner.tokens [20] & ~_02678_;
	assign _02680_ = _02679_ | _02674_;
	assign _02681_ = _01673_ | _01281_;
	assign _02683_ = _02681_ | _01506_;
	assign _02684_ = _02683_ | _01288_;
	assign _02685_ = _01274_ & ~_02684_;
	assign _02686_ = _01678_ | _01281_;
	assign _02687_ = _02686_ | ~_01284_;
	assign _02688_ = _02687_ | _01288_;
	assign _02689_ = _01274_ & ~_02688_;
	assign _02690_ = \mchip.design.owner.tokens [20] & ~_02689_;
	assign _02691_ = _02690_ | _02685_;
	assign _02692_ = (_00199_ ? _02680_ : _02691_);
	assign _02694_ = _01688_ | _01311_;
	assign _02695_ = _02694_ | _01523_;
	assign _02696_ = _02695_ | _01318_;
	assign _02697_ = _01303_ & ~_02696_;
	assign _02698_ = _01693_ | _01311_;
	assign _02699_ = _02698_ | ~_01314_;
	assign _02700_ = _02699_ | _01318_;
	assign _02701_ = _01303_ & ~_02700_;
	assign _02702_ = \mchip.design.owner.tokens [20] & ~_02701_;
	assign _02703_ = _02702_ | _02697_;
	assign _02705_ = (_00131_ ? _02692_ : _02703_);
	assign _02706_ = _01703_ | _01341_;
	assign _02707_ = _02706_ | _01540_;
	assign _02708_ = _02707_ | _01346_;
	assign _02709_ = _01349_ & ~_02708_;
	assign _02710_ = _01708_ | _01341_;
	assign _02711_ = _02710_ | _01540_;
	assign _02712_ = _02711_ | _01346_;
	assign _02713_ = _01349_ & ~_02712_;
	assign _02714_ = \mchip.design.owner.tokens [20] & ~_02713_;
	assign _02716_ = _02714_ | _02709_;
	assign _02717_ = (_06005_ ? _02705_ : _02716_);
	assign _02718_ = _01718_ | _01374_;
	assign _02719_ = _02718_ | ~_01377_;
	assign _02720_ = _02719_ | _01380_;
	assign _02721_ = _01382_ & ~_02720_;
	assign _02722_ = _01726_ | _01374_;
	assign _02723_ = _02722_ | ~_01377_;
	assign _02724_ = _02723_ | _01380_;
	assign _02725_ = _01382_ & ~_02724_;
	assign _02727_ = \mchip.design.owner.tokens [20] & ~_02725_;
	assign _02728_ = _02727_ | _02721_;
	assign _02729_ = (_05934_ ? _02717_ : _02728_);
	assign _02730_ = _01736_ | _01404_;
	assign _02731_ = _02730_ | _01575_;
	assign _02732_ = _02731_ | _01398_;
	assign _02733_ = _01410_ & ~_02732_;
	assign _02734_ = _01743_ | _01404_;
	assign _02735_ = _02734_ | _01575_;
	assign _02736_ = _02735_ | _01398_;
	assign _02738_ = _01410_ & ~_02736_;
	assign _02739_ = \mchip.design.owner.tokens [20] & ~_02738_;
	assign _02740_ = _02739_ | _02733_;
	assign _00024_ = (_05827_ ? _02729_ : _02740_);
	assign _02741_ = _01752_ | _01254_;
	assign _02742_ = _02741_ | _01490_;
	assign _02743_ = _02742_ | _01261_;
	assign _02744_ = _01243_ & ~_02743_;
	assign _02745_ = \mchip.design.owner.tokens [21] & ~_02678_;
	assign _02746_ = _02745_ | _02744_;
	assign _02748_ = _01761_ | _01281_;
	assign _02749_ = _02748_ | _01506_;
	assign _02750_ = _02749_ | _01288_;
	assign _02751_ = _01274_ & ~_02750_;
	assign _02752_ = \mchip.design.owner.tokens [21] & ~_02689_;
	assign _02753_ = _02752_ | _02751_;
	assign _02754_ = (_00199_ ? _02746_ : _02753_);
	assign _02755_ = _01771_ | _01311_;
	assign _02756_ = _02755_ | _01523_;
	assign _02757_ = _02756_ | _01318_;
	assign _02759_ = _01303_ & ~_02757_;
	assign _02760_ = \mchip.design.owner.tokens [21] & ~_02701_;
	assign _02761_ = _02760_ | _02759_;
	assign _02762_ = (_00131_ ? _02754_ : _02761_);
	assign _02763_ = _01781_ | _01341_;
	assign _02764_ = _02763_ | _01540_;
	assign _02765_ = _02764_ | _01346_;
	assign _02766_ = _01349_ & ~_02765_;
	assign _02767_ = \mchip.design.owner.tokens [21] & ~_02713_;
	assign _02768_ = _02767_ | _02766_;
	assign _02770_ = (_06005_ ? _02762_ : _02768_);
	assign _02771_ = _01791_ | _01374_;
	assign _02772_ = _02771_ | ~_01377_;
	assign _02773_ = _02772_ | _01380_;
	assign _02774_ = _01382_ & ~_02773_;
	assign _02775_ = \mchip.design.owner.tokens [21] & ~_02725_;
	assign _02776_ = _02775_ | _02774_;
	assign _02777_ = (_05934_ ? _02770_ : _02776_);
	assign _02778_ = _01801_ | _01404_;
	assign _02779_ = _02778_ | _01575_;
	assign _02781_ = _02779_ | _01398_;
	assign _02782_ = _01410_ & ~_02781_;
	assign _02783_ = \mchip.design.owner.tokens [21] & ~_02738_;
	assign _02784_ = _02783_ | _02782_;
	assign _00025_ = (_05827_ ? _02777_ : _02784_);
	assign _02785_ = _01809_ | _01254_;
	assign _02786_ = _02785_ | _01490_;
	assign _02787_ = _02786_ | _01261_;
	assign _02788_ = _01243_ & ~_02787_;
	assign _02789_ = _01814_ | _01254_;
	assign _02791_ = _02789_ | ~_01257_;
	assign _02792_ = _02791_ | _01261_;
	assign _02793_ = _01243_ & ~_02792_;
	assign _02794_ = \mchip.design.owner.tokens [22] & ~_02793_;
	assign _02795_ = _02794_ | _02788_;
	assign _02796_ = _01822_ | _01281_;
	assign _02797_ = _02796_ | _01506_;
	assign _02798_ = _02797_ | _01288_;
	assign _02799_ = _01274_ & ~_02798_;
	assign _02800_ = _01827_ | _01281_;
	assign _02802_ = _02800_ | ~_01284_;
	assign _02803_ = _02802_ | _01288_;
	assign _02804_ = _01274_ & ~_02803_;
	assign _02805_ = \mchip.design.owner.tokens [22] & ~_02804_;
	assign _02806_ = _02805_ | _02799_;
	assign _02807_ = (_00199_ ? _02795_ : _02806_);
	assign _02808_ = _01836_ | _01311_;
	assign _02809_ = _02808_ | _01523_;
	assign _02810_ = _02809_ | _01318_;
	assign _02811_ = _01303_ & ~_02810_;
	assign _02813_ = _01841_ | _01311_;
	assign _02814_ = _02813_ | ~_01314_;
	assign _02815_ = _02814_ | _01318_;
	assign _02816_ = _01303_ & ~_02815_;
	assign _02817_ = \mchip.design.owner.tokens [22] & ~_02816_;
	assign _02818_ = _02817_ | _02811_;
	assign _02819_ = (_00131_ ? _02807_ : _02818_);
	assign _02820_ = _01850_ | _01341_;
	assign _02821_ = _02820_ | _01540_;
	assign _02822_ = _02821_ | _01346_;
	assign _02824_ = _01349_ & ~_02822_;
	assign _02825_ = _01855_ | _01341_;
	assign _02826_ = _02825_ | _01540_;
	assign _02827_ = _02826_ | _01346_;
	assign _02828_ = _01349_ & ~_02827_;
	assign _02829_ = \mchip.design.owner.tokens [22] & ~_02828_;
	assign _02830_ = _02829_ | _02824_;
	assign _02831_ = (_06005_ ? _02819_ : _02830_);
	assign _02832_ = _01864_ | _01374_;
	assign _02833_ = _02832_ | ~_01377_;
	assign _02835_ = _02833_ | _01380_;
	assign _02836_ = _01382_ & ~_02835_;
	assign _02837_ = _01871_ | _01374_;
	assign _02838_ = _02837_ | ~_01377_;
	assign _02839_ = _02838_ | _01380_;
	assign _02840_ = _01382_ & ~_02839_;
	assign _02841_ = \mchip.design.owner.tokens [22] & ~_02840_;
	assign _02842_ = _02841_ | _02836_;
	assign _02843_ = (_05934_ ? _02831_ : _02842_);
	assign _02844_ = _01880_ | _01404_;
	assign _02846_ = _02844_ | _01575_;
	assign _02847_ = _02846_ | _01398_;
	assign _02848_ = _01410_ & ~_02847_;
	assign _02849_ = _01886_ | _01404_;
	assign _02850_ = _02849_ | _01575_;
	assign _02851_ = _02850_ | _01398_;
	assign _02852_ = _01410_ & ~_02851_;
	assign _02853_ = \mchip.design.owner.tokens [22] & ~_02852_;
	assign _02854_ = _02853_ | _02848_;
	assign _00026_ = (_05827_ ? _02843_ : _02854_);
	assign _02856_ = _01894_ | _01254_;
	assign _02857_ = _02856_ | _01490_;
	assign _02858_ = _02857_ | _01261_;
	assign _02859_ = _01243_ & ~_02858_;
	assign _02860_ = \mchip.design.owner.tokens [23] & ~_02793_;
	assign _02861_ = _02860_ | _02859_;
	assign _02862_ = _01902_ | _01281_;
	assign _02863_ = _02862_ | _01506_;
	assign _02864_ = _02863_ | _01288_;
	assign _02865_ = _01274_ & ~_02864_;
	assign _02867_ = \mchip.design.owner.tokens [23] & ~_02804_;
	assign _02868_ = _02867_ | _02865_;
	assign _02869_ = (_00199_ ? _02861_ : _02868_);
	assign _02870_ = _01911_ | _01311_;
	assign _02871_ = _02870_ | _01523_;
	assign _02872_ = _02871_ | _01318_;
	assign _02873_ = _01303_ & ~_02872_;
	assign _02874_ = \mchip.design.owner.tokens [23] & ~_02816_;
	assign _02875_ = _02874_ | _02873_;
	assign _02876_ = (_00131_ ? _02869_ : _02875_);
	assign _02878_ = _01920_ | _01341_;
	assign _02879_ = _02878_ | _01540_;
	assign _02880_ = _02879_ | _01346_;
	assign _02881_ = _01349_ & ~_02880_;
	assign _02882_ = \mchip.design.owner.tokens [23] & ~_02828_;
	assign _02883_ = _02882_ | _02881_;
	assign _02884_ = (_06005_ ? _02876_ : _02883_);
	assign _02885_ = _01929_ | _01374_;
	assign _02886_ = _02885_ | ~_01377_;
	assign _02887_ = _02886_ | _01380_;
	assign _02889_ = _01382_ & ~_02887_;
	assign _02890_ = \mchip.design.owner.tokens [23] & ~_02840_;
	assign _02891_ = _02890_ | _02889_;
	assign _02892_ = (_05934_ ? _02884_ : _02891_);
	assign _02893_ = _01938_ | _01404_;
	assign _02894_ = _02893_ | _01575_;
	assign _02895_ = _02894_ | _01398_;
	assign _02896_ = _01410_ & ~_02895_;
	assign _02897_ = \mchip.design.owner.tokens [23] & ~_02852_;
	assign _02898_ = _02897_ | _02896_;
	assign _00027_ = (_05827_ ? _02892_ : _02898_);
	assign _02900_ = _01946_ | _01254_;
	assign _02901_ = _02900_ | _01490_;
	assign _02902_ = _02901_ | _01261_;
	assign _02903_ = _01243_ & ~_02902_;
	assign _02904_ = _01951_ | _01254_;
	assign _02905_ = _02904_ | ~_01257_;
	assign _02906_ = _02905_ | _01261_;
	assign _02907_ = _01243_ & ~_02906_;
	assign _02908_ = \mchip.design.owner.tokens [24] & ~_02907_;
	assign _02910_ = _02908_ | _02903_;
	assign _02911_ = _01959_ | _01281_;
	assign _02912_ = _02911_ | _01506_;
	assign _02913_ = _02912_ | _01288_;
	assign _02914_ = _01274_ & ~_02913_;
	assign _02915_ = _01964_ | _01281_;
	assign _02916_ = _02915_ | ~_01284_;
	assign _02917_ = _02916_ | _01288_;
	assign _02918_ = _01274_ & ~_02917_;
	assign _02919_ = \mchip.design.owner.tokens [24] & ~_02918_;
	assign _02921_ = _02919_ | _02914_;
	assign _02922_ = (_00199_ ? _02910_ : _02921_);
	assign _02923_ = _01973_ | _01311_;
	assign _02924_ = _02923_ | _01523_;
	assign _02925_ = _02924_ | _01318_;
	assign _02926_ = _01303_ & ~_02925_;
	assign _02927_ = _01978_ | _01311_;
	assign _02928_ = _02927_ | ~_01314_;
	assign _02929_ = _02928_ | _01318_;
	assign _02930_ = _01303_ & ~_02929_;
	assign _02932_ = \mchip.design.owner.tokens [24] & ~_02930_;
	assign _02933_ = _02932_ | _02926_;
	assign _02934_ = (_00131_ ? _02922_ : _02933_);
	assign _02935_ = _01987_ | _01341_;
	assign _02936_ = _02935_ | _01540_;
	assign _02937_ = _02936_ | _01346_;
	assign _02938_ = _01349_ & ~_02937_;
	assign _02939_ = _01992_ | _01341_;
	assign _02940_ = _02939_ | _01540_;
	assign _02941_ = _02940_ | _01346_;
	assign _02943_ = _01349_ & ~_02941_;
	assign _02944_ = \mchip.design.owner.tokens [24] & ~_02943_;
	assign _02945_ = _02944_ | _02938_;
	assign _02946_ = (_06005_ ? _02934_ : _02945_);
	assign _02947_ = _02001_ | _01374_;
	assign _02948_ = _02947_ | ~_01377_;
	assign _02949_ = _02948_ | _01380_;
	assign _02950_ = _01382_ & ~_02949_;
	assign _02951_ = _02007_ | _01374_;
	assign _02952_ = _02951_ | ~_01377_;
	assign _02954_ = _02952_ | _01380_;
	assign _02955_ = _01382_ & ~_02954_;
	assign _02956_ = \mchip.design.owner.tokens [24] & ~_02955_;
	assign _02957_ = _02956_ | _02950_;
	assign _02958_ = (_05934_ ? _02946_ : _02957_);
	assign _02959_ = _02016_ | _01404_;
	assign _02960_ = _02959_ | _01575_;
	assign _02961_ = _02960_ | _01398_;
	assign _02962_ = _01410_ & ~_02961_;
	assign _02963_ = _02022_ | _01404_;
	assign _02965_ = _02963_ | _01575_;
	assign _02966_ = _02965_ | _01398_;
	assign _02967_ = _01410_ & ~_02966_;
	assign _02968_ = \mchip.design.owner.tokens [24] & ~_02967_;
	assign _02969_ = _02968_ | _02962_;
	assign _00028_ = (_05827_ ? _02958_ : _02969_);
	assign _02970_ = _02030_ | _01254_;
	assign _02971_ = _02970_ | _01490_;
	assign _02972_ = _02971_ | _01261_;
	assign _02973_ = _01243_ & ~_02972_;
	assign _02975_ = \mchip.design.owner.tokens [25] & ~_02907_;
	assign _02976_ = _02975_ | _02973_;
	assign _02977_ = _02038_ | _01281_;
	assign _02978_ = _02977_ | _01506_;
	assign _02979_ = _02978_ | _01288_;
	assign _02980_ = _01274_ & ~_02979_;
	assign _02981_ = \mchip.design.owner.tokens [25] & ~_02918_;
	assign _02982_ = _02981_ | _02980_;
	assign _02983_ = (_00199_ ? _02976_ : _02982_);
	assign _02984_ = _02047_ | _01311_;
	assign _02986_ = _02984_ | _01523_;
	assign _02987_ = _02986_ | _01318_;
	assign _02988_ = _01303_ & ~_02987_;
	assign _02989_ = \mchip.design.owner.tokens [25] & ~_02930_;
	assign _02990_ = _02989_ | _02988_;
	assign _02991_ = (_00131_ ? _02983_ : _02990_);
	assign _02992_ = _02056_ | _01341_;
	assign _02993_ = _02992_ | _01540_;
	assign _02994_ = _02993_ | _01346_;
	assign _02995_ = _01349_ & ~_02994_;
	assign _02997_ = \mchip.design.owner.tokens [25] & ~_02943_;
	assign _02998_ = _02997_ | _02995_;
	assign _02999_ = (_06005_ ? _02991_ : _02998_);
	assign _03000_ = _02065_ | _01374_;
	assign _03001_ = _03000_ | ~_01377_;
	assign _03002_ = _03001_ | _01380_;
	assign _03003_ = _01382_ & ~_03002_;
	assign _03004_ = \mchip.design.owner.tokens [25] & ~_02955_;
	assign _03005_ = _03004_ | _03003_;
	assign _03006_ = (_05934_ ? _02999_ : _03005_);
	assign _03008_ = _02074_ | _01404_;
	assign _03009_ = _03008_ | _01575_;
	assign _03010_ = _03009_ | _01398_;
	assign _03011_ = _01410_ & ~_03010_;
	assign _03012_ = \mchip.design.owner.tokens [25] & ~_02967_;
	assign _03013_ = _03012_ | _03011_;
	assign _00029_ = (_05827_ ? _03006_ : _03013_);
	assign _03014_ = _02081_ | _01254_;
	assign _03015_ = _03014_ | _01490_;
	assign _03016_ = _03015_ | _01261_;
	assign _03018_ = _01243_ & ~_03016_;
	assign _03019_ = _02086_ | _01254_;
	assign _03020_ = _03019_ | ~_01257_;
	assign _03021_ = _03020_ | _01261_;
	assign _03022_ = _01243_ & ~_03021_;
	assign _03023_ = \mchip.design.owner.tokens [26] & ~_03022_;
	assign _03024_ = _03023_ | _03018_;
	assign _03025_ = _02093_ | _01281_;
	assign _03026_ = _03025_ | _01506_;
	assign _03027_ = _03026_ | _01288_;
	assign _03029_ = _01274_ & ~_03027_;
	assign _03030_ = _01281_ | _01951_;
	assign _03031_ = _03030_ | ~_01284_;
	assign _03032_ = _03031_ | _01288_;
	assign _03033_ = _01274_ & ~_03032_;
	assign _03034_ = \mchip.design.owner.tokens [26] & ~_03033_;
	assign _03035_ = _03034_ | _03029_;
	assign _03036_ = (_00199_ ? _03024_ : _03035_);
	assign _03037_ = _02105_ | _01311_;
	assign _03038_ = _03037_ | _01523_;
	assign _03040_ = _03038_ | _01318_;
	assign _03041_ = _01303_ & ~_03040_;
	assign _03042_ = _01964_ | _01311_;
	assign _03043_ = _03042_ | ~_01314_;
	assign _03044_ = _03043_ | _01318_;
	assign _03045_ = _01303_ & ~_03044_;
	assign _03046_ = \mchip.design.owner.tokens [26] & ~_03045_;
	assign _03047_ = _03046_ | _03041_;
	assign _03048_ = (_00131_ ? _03036_ : _03047_);
	assign _03049_ = _02117_ | _01341_;
	assign _03051_ = _03049_ | _01540_;
	assign _03052_ = _03051_ | _01346_;
	assign _03053_ = _01349_ & ~_03052_;
	assign _03054_ = _02122_ | _01341_;
	assign _03055_ = _03054_ | _01540_;
	assign _03056_ = _03055_ | _01346_;
	assign _03057_ = _01349_ & ~_03056_;
	assign _03058_ = \mchip.design.owner.tokens [26] & ~_03057_;
	assign _03059_ = _03058_ | _03053_;
	assign _03060_ = (_06005_ ? _03048_ : _03059_);
	assign _03062_ = _02130_ | _01374_;
	assign _03063_ = _03062_ | ~_01377_;
	assign _03064_ = _03063_ | _01380_;
	assign _03065_ = _01382_ & ~_03064_;
	assign _03066_ = _02135_ | _01374_;
	assign _03067_ = _03066_ | ~_01377_;
	assign _03068_ = _03067_ | _01380_;
	assign _03069_ = _01382_ & ~_03068_;
	assign _03070_ = \mchip.design.owner.tokens [26] & ~_03069_;
	assign _03071_ = _03070_ | _03065_;
	assign _03073_ = (_05934_ ? _03060_ : _03071_);
	assign _03074_ = _02143_ | _01404_;
	assign _03075_ = _03074_ | _01575_;
	assign _03076_ = _03075_ | _01398_;
	assign _03077_ = _01410_ & ~_03076_;
	assign _03078_ = _02148_ | _01404_;
	assign _03079_ = _03078_ | _01575_;
	assign _03080_ = _03079_ | _01398_;
	assign _03081_ = _01410_ & ~_03080_;
	assign _03082_ = \mchip.design.owner.tokens [26] & ~_03081_;
	assign _03084_ = _03082_ | _03077_;
	assign _00030_ = (_05827_ ? _03073_ : _03084_);
	assign _03085_ = _02155_ | _01254_;
	assign _03086_ = _03085_ | _01490_;
	assign _03087_ = _03086_ | _01261_;
	assign _03088_ = _01243_ & ~_03087_;
	assign _03089_ = \mchip.design.owner.tokens [27] & ~_03022_;
	assign _03090_ = _03089_ | _03088_;
	assign _03091_ = _02162_ | _01281_;
	assign _03092_ = _03091_ | _01506_;
	assign _03094_ = _03092_ | _01288_;
	assign _03095_ = _01274_ & ~_03094_;
	assign _03096_ = \mchip.design.owner.tokens [27] & ~_03033_;
	assign _03097_ = _03096_ | _03095_;
	assign _03098_ = (_00199_ ? _03090_ : _03097_);
	assign _03099_ = _02170_ | _01311_;
	assign _03100_ = _03099_ | _01523_;
	assign _03101_ = _03100_ | _01318_;
	assign _03102_ = _01303_ & ~_03101_;
	assign _03103_ = \mchip.design.owner.tokens [27] & ~_03045_;
	assign _03105_ = _03103_ | _03102_;
	assign _03106_ = (_00131_ ? _03098_ : _03105_);
	assign _03107_ = _02178_ | _01341_;
	assign _03108_ = _03107_ | _01540_;
	assign _03109_ = _03108_ | _01346_;
	assign _03110_ = _01349_ & ~_03109_;
	assign _03111_ = \mchip.design.owner.tokens [27] & ~_03057_;
	assign _03112_ = _03111_ | _03110_;
	assign _03113_ = (_06005_ ? _03106_ : _03112_);
	assign _03114_ = _02186_ | _01374_;
	assign _03116_ = _03114_ | ~_01377_;
	assign _03117_ = _03116_ | _01380_;
	assign _03118_ = _01382_ & ~_03117_;
	assign _03119_ = \mchip.design.owner.tokens [27] & ~_03069_;
	assign _03120_ = _03119_ | _03118_;
	assign _03121_ = (_05934_ ? _03113_ : _03120_);
	assign _03122_ = _02194_ | _01404_;
	assign _03123_ = _03122_ | _01575_;
	assign _03124_ = _03123_ | _01398_;
	assign _03125_ = _01410_ & ~_03124_;
	assign _03126_ = \mchip.design.owner.tokens [27] & ~_03081_;
	assign _03127_ = _03126_ | _03125_;
	assign _00031_ = (_05827_ ? _03121_ : _03127_);
	assign _03128_ = _02201_ | _01254_;
	assign _03129_ = _03128_ | _01490_;
	assign _03130_ = _03129_ | _01261_;
	assign _03131_ = _01243_ & ~_03130_;
	assign _03132_ = _02206_ | _01254_;
	assign _03133_ = _03132_ | ~_01257_;
	assign _03134_ = _03133_ | _01261_;
	assign _03136_ = _01243_ & ~_03134_;
	assign _03137_ = \mchip.design.owner.tokens [28] & ~_03136_;
	assign _03138_ = _03137_ | _03131_;
	assign _03139_ = _02213_ | _01281_;
	assign _03140_ = _03139_ | _01506_;
	assign _03141_ = _03140_ | _01288_;
	assign _03142_ = _01274_ & ~_03141_;
	assign _03143_ = _02218_ | _01281_;
	assign _03144_ = _03143_ | ~_01284_;
	assign _03145_ = _03144_ | _01288_;
	assign _03147_ = _01274_ & ~_03145_;
	assign _03148_ = \mchip.design.owner.tokens [28] & ~_03147_;
	assign _03149_ = _03148_ | _03142_;
	assign _03150_ = (_00199_ ? _03138_ : _03149_);
	assign _03151_ = _02226_ | _01311_;
	assign _03152_ = _03151_ | _01523_;
	assign _03153_ = _03152_ | _01318_;
	assign _03154_ = _01303_ & ~_03153_;
	assign _03155_ = _02231_ | _01311_;
	assign _03156_ = _03155_ | ~_01314_;
	assign _03158_ = _03156_ | _01318_;
	assign _03159_ = _01303_ & ~_03158_;
	assign _03160_ = \mchip.design.owner.tokens [28] & ~_03159_;
	assign _03161_ = _03160_ | _03154_;
	assign _03162_ = (_00131_ ? _03150_ : _03161_);
	assign _03163_ = _02239_ | _01341_;
	assign _03164_ = _03163_ | _01540_;
	assign _03165_ = _03164_ | _01346_;
	assign _03166_ = _01349_ & ~_03165_;
	assign _03167_ = _02244_ | _01341_;
	assign _03169_ = _03167_ | _01540_;
	assign _03170_ = _03169_ | _01346_;
	assign _03171_ = _01349_ & ~_03170_;
	assign _03172_ = \mchip.design.owner.tokens [28] & ~_03171_;
	assign _03173_ = _03172_ | _03166_;
	assign _03174_ = (_06005_ ? _03162_ : _03173_);
	assign _03175_ = _02252_ | _01374_;
	assign _03176_ = _03175_ | ~_01377_;
	assign _03177_ = _03176_ | _01380_;
	assign _03178_ = _01382_ & ~_03177_;
	assign _03180_ = _02257_ | _01374_;
	assign _03181_ = _03180_ | ~_01377_;
	assign _03182_ = _03181_ | _01380_;
	assign _03183_ = _01382_ & ~_03182_;
	assign _03184_ = \mchip.design.owner.tokens [28] & ~_03183_;
	assign _03185_ = _03184_ | _03178_;
	assign _03186_ = (_05934_ ? _03174_ : _03185_);
	assign _03187_ = _02265_ | _01404_;
	assign _03188_ = _03187_ | _01575_;
	assign _03189_ = _03188_ | _01398_;
	assign _03191_ = _01410_ & ~_03189_;
	assign _03192_ = _02270_ | _01404_;
	assign _03193_ = _03192_ | _01575_;
	assign _03194_ = _03193_ | _01398_;
	assign _03195_ = _01410_ & ~_03194_;
	assign _03196_ = \mchip.design.owner.tokens [28] & ~_03195_;
	assign _03197_ = _03196_ | _03191_;
	assign _00032_ = (_05827_ ? _03186_ : _03197_);
	assign _03198_ = _02277_ | _01254_;
	assign _03199_ = _03198_ | _01490_;
	assign _03201_ = _03199_ | _01261_;
	assign _03202_ = _01243_ & ~_03201_;
	assign _03203_ = \mchip.design.owner.tokens [29] & ~_03136_;
	assign _03204_ = _03203_ | _03202_;
	assign _03205_ = _02284_ | _01281_;
	assign _03206_ = _03205_ | _01506_;
	assign _03207_ = _03206_ | _01288_;
	assign _03208_ = _01274_ & ~_03207_;
	assign _03209_ = \mchip.design.owner.tokens [29] & ~_03147_;
	assign _03210_ = _03209_ | _03208_;
	assign _03212_ = (_00199_ ? _03204_ : _03210_);
	assign _03213_ = _02292_ | _01311_;
	assign _03214_ = _03213_ | _01523_;
	assign _03215_ = _03214_ | _01318_;
	assign _03216_ = _01303_ & ~_03215_;
	assign _03217_ = \mchip.design.owner.tokens [29] & ~_03159_;
	assign _03218_ = _03217_ | _03216_;
	assign _03219_ = (_00131_ ? _03212_ : _03218_);
	assign _03220_ = _02300_ | _01341_;
	assign _03221_ = _03220_ | _01540_;
	assign _03223_ = _03221_ | _01346_;
	assign _03224_ = _01349_ & ~_03223_;
	assign _03225_ = \mchip.design.owner.tokens [29] & ~_03171_;
	assign _03226_ = _03225_ | _03224_;
	assign _03227_ = (_06005_ ? _03219_ : _03226_);
	assign _03228_ = _02308_ | _01374_;
	assign _03229_ = _03228_ | ~_01377_;
	assign _03230_ = _03229_ | _01380_;
	assign _03231_ = _01382_ & ~_03230_;
	assign _03232_ = \mchip.design.owner.tokens [29] & ~_03183_;
	assign _03234_ = _03232_ | _03231_;
	assign _03235_ = (_05934_ ? _03227_ : _03234_);
	assign _03236_ = _02316_ | _01404_;
	assign _03237_ = _03236_ | _01575_;
	assign _03238_ = _03237_ | _01398_;
	assign _03239_ = _01410_ & ~_03238_;
	assign _03240_ = \mchip.design.owner.tokens [29] & ~_03195_;
	assign _03241_ = _03240_ | _03239_;
	assign _00033_ = (_05827_ ? _03235_ : _03241_);
	assign _03242_ = _02323_ | _01254_;
	assign _03244_ = _03242_ | _01490_;
	assign _03245_ = _03244_ | _01261_;
	assign _03246_ = _01243_ & ~_03245_;
	assign _03247_ = _02328_ | _01254_;
	assign _03248_ = _03247_ | ~_01257_;
	assign _03249_ = _03248_ | _01261_;
	assign _03250_ = _01243_ & ~_03249_;
	assign _03251_ = \mchip.design.owner.tokens [30] & ~_03250_;
	assign _03252_ = _03251_ | _03246_;
	assign _03253_ = _02335_ | _01281_;
	assign _03255_ = _03253_ | _01506_;
	assign _03256_ = _03255_ | _01288_;
	assign _03257_ = _01274_ & ~_03256_;
	assign _03258_ = _02340_ | _01281_;
	assign _03259_ = _03258_ | ~_01284_;
	assign _03260_ = _03259_ | _01288_;
	assign _03261_ = _01274_ & ~_03260_;
	assign _03262_ = \mchip.design.owner.tokens [30] & ~_03261_;
	assign _03263_ = _03262_ | _03257_;
	assign _03264_ = (_00199_ ? _03252_ : _03263_);
	assign _03266_ = _02348_ | _01311_;
	assign _03267_ = _03266_ | _01523_;
	assign _03268_ = _03267_ | _01318_;
	assign _03269_ = _01303_ & ~_03268_;
	assign _03270_ = _02353_ | _01311_;
	assign _03271_ = _03270_ | ~_01314_;
	assign _03272_ = _03271_ | _01318_;
	assign _03273_ = _01303_ & ~_03272_;
	assign _03274_ = \mchip.design.owner.tokens [30] & ~_03273_;
	assign _03275_ = _03274_ | _03269_;
	assign _03277_ = (_00131_ ? _03264_ : _03275_);
	assign _03278_ = _02361_ | _01341_;
	assign _03279_ = _03278_ | _01540_;
	assign _03280_ = _03279_ | _01346_;
	assign _03281_ = _01349_ & ~_03280_;
	assign _03282_ = _02366_ | _01341_;
	assign _03283_ = _03282_ | _01540_;
	assign _03284_ = _03283_ | _01346_;
	assign _03285_ = _01349_ & ~_03284_;
	assign _03286_ = \mchip.design.owner.tokens [30] & ~_03285_;
	assign _03288_ = _03286_ | _03281_;
	assign _03289_ = (_06005_ ? _03277_ : _03288_);
	assign _03290_ = _02374_ | _01374_;
	assign _03291_ = _03290_ | ~_01377_;
	assign _03292_ = _03291_ | _01380_;
	assign _03293_ = _01382_ & ~_03292_;
	assign _03294_ = _02379_ | _01374_;
	assign _03295_ = _03294_ | ~_01377_;
	assign _03296_ = _03295_ | _01380_;
	assign _03297_ = _01382_ & ~_03296_;
	assign _03299_ = \mchip.design.owner.tokens [30] & ~_03297_;
	assign _03300_ = _03299_ | _03293_;
	assign _03301_ = (_05934_ ? _03289_ : _03300_);
	assign _03302_ = _02387_ | _01404_;
	assign _03303_ = _03302_ | _01575_;
	assign _03304_ = _03303_ | _01398_;
	assign _03305_ = _01410_ & ~_03304_;
	assign _03306_ = _02392_ | _01404_;
	assign _03307_ = _03306_ | _01575_;
	assign _03308_ = _03307_ | _01398_;
	assign _03310_ = _01410_ & ~_03308_;
	assign _03311_ = \mchip.design.owner.tokens [30] & ~_03310_;
	assign _03312_ = _03311_ | _03305_;
	assign _00035_ = (_05827_ ? _03301_ : _03312_);
	assign _03313_ = _02399_ | _01254_;
	assign _03314_ = _03313_ | _01490_;
	assign _03315_ = _03314_ | _01261_;
	assign _03316_ = _01243_ & ~_03315_;
	assign _03317_ = \mchip.design.owner.tokens [31] & ~_03250_;
	assign _03318_ = _03317_ | _03316_;
	assign _03320_ = _02406_ | _01281_;
	assign _03321_ = _03320_ | _01506_;
	assign _03322_ = _03321_ | _01288_;
	assign _03323_ = _01274_ & ~_03322_;
	assign _03324_ = \mchip.design.owner.tokens [31] & ~_03261_;
	assign _03325_ = _03324_ | _03323_;
	assign _03326_ = (_00199_ ? _03318_ : _03325_);
	assign _03327_ = _02414_ | _01311_;
	assign _03328_ = _03327_ | _01523_;
	assign _03329_ = _03328_ | _01318_;
	assign _03331_ = _01303_ & ~_03329_;
	assign _03332_ = \mchip.design.owner.tokens [31] & ~_03273_;
	assign _03333_ = _03332_ | _03331_;
	assign _03334_ = (_00131_ ? _03326_ : _03333_);
	assign _03335_ = _02422_ | _01341_;
	assign _03336_ = _03335_ | _01540_;
	assign _03337_ = _03336_ | _01346_;
	assign _03338_ = _01349_ & ~_03337_;
	assign _03339_ = \mchip.design.owner.tokens [31] & ~_03285_;
	assign _03340_ = _03339_ | _03338_;
	assign _03342_ = (_06005_ ? _03334_ : _03340_);
	assign _03343_ = _02430_ | _01374_;
	assign _03344_ = _03343_ | ~_01377_;
	assign _03345_ = _03344_ | _01380_;
	assign _03346_ = _01382_ & ~_03345_;
	assign _03347_ = \mchip.design.owner.tokens [31] & ~_03297_;
	assign _03348_ = _03347_ | _03346_;
	assign _03349_ = (_05934_ ? _03342_ : _03348_);
	assign _03350_ = _02438_ | _01404_;
	assign _03351_ = _03350_ | _01575_;
	assign _03353_ = _03351_ | _01398_;
	assign _03354_ = _01410_ & ~_03353_;
	assign _03355_ = \mchip.design.owner.tokens [31] & ~_03310_;
	assign _03356_ = _03355_ | _03354_;
	assign _00036_ = (_05827_ ? _03349_ : _03356_);
	assign _03357_ = _02445_ | _01254_;
	assign _03358_ = _03357_ | _01490_;
	assign _03359_ = _03358_ | _01261_;
	assign _03360_ = _01243_ & ~_03359_;
	assign _03361_ = _01515_ | _01254_;
	assign _03363_ = _03361_ | ~_01257_;
	assign _03364_ = _03363_ | _01261_;
	assign _03365_ = _01243_ & ~_03364_;
	assign _03366_ = \mchip.design.owner.tokens [32] & ~_03365_;
	assign _03367_ = _03366_ | _03360_;
	assign _03368_ = _02456_ | _01281_;
	assign _03369_ = _03368_ | _01506_;
	assign _03370_ = _03369_ | _01288_;
	assign _03371_ = _01274_ & ~_03370_;
	assign _03372_ = _01532_ | _01281_;
	assign _03374_ = _03372_ | ~_01284_;
	assign _03375_ = _03374_ | _01288_;
	assign _03376_ = _01274_ & ~_03375_;
	assign _03377_ = \mchip.design.owner.tokens [32] & ~_03376_;
	assign _03378_ = _03377_ | _03371_;
	assign _03379_ = (_00199_ ? _03367_ : _03378_);
	assign _03380_ = _02468_ | _01311_;
	assign _03381_ = _03380_ | _01523_;
	assign _03382_ = _03381_ | _01318_;
	assign _03383_ = _01303_ & ~_03382_;
	assign _03385_ = _02473_ | _01311_;
	assign _03386_ = _03385_ | ~_01314_;
	assign _03387_ = _03386_ | _01318_;
	assign _03388_ = _01303_ & ~_03387_;
	assign _03389_ = \mchip.design.owner.tokens [32] & ~_03388_;
	assign _03390_ = _03389_ | _03383_;
	assign _03391_ = (_00131_ ? _03379_ : _03390_);
	assign _03392_ = _02481_ | _01341_;
	assign _03393_ = _03392_ | _01540_;
	assign _03394_ = _03393_ | _01346_;
	assign _03396_ = _01349_ & ~_03394_;
	assign _03397_ = _02486_ | _01341_;
	assign _03398_ = _03397_ | _01540_;
	assign _03399_ = _03398_ | _01346_;
	assign _03400_ = _01349_ & ~_03399_;
	assign _03401_ = \mchip.design.owner.tokens [32] & ~_03400_;
	assign _03402_ = _03401_ | _03396_;
	assign _03403_ = (_06005_ ? _03391_ : _03402_);
	assign _03404_ = _02494_ | _01374_;
	assign _03405_ = _03404_ | ~_01377_;
	assign _03407_ = _03405_ | _01380_;
	assign _03408_ = _01382_ & ~_03407_;
	assign _03409_ = _02499_ | _01374_;
	assign _03410_ = _03409_ | ~_01377_;
	assign _03411_ = _03410_ | _01380_;
	assign _03412_ = _01382_ & ~_03411_;
	assign _03413_ = \mchip.design.owner.tokens [32] & ~_03412_;
	assign _03414_ = _03413_ | _03408_;
	assign _03415_ = (_05934_ ? _03403_ : _03414_);
	assign _03416_ = _02507_ | _01404_;
	assign _03418_ = _03416_ | _01575_;
	assign _03419_ = _03418_ | _01398_;
	assign _03420_ = _01410_ & ~_03419_;
	assign _03421_ = _02512_ | _01404_;
	assign _03422_ = _03421_ | _01575_;
	assign _03423_ = _03422_ | _01398_;
	assign _03424_ = _01410_ & ~_03423_;
	assign _03425_ = \mchip.design.owner.tokens [32] & ~_03424_;
	assign _03426_ = _03425_ | _03420_;
	assign _00037_ = (_05827_ ? _03415_ : _03426_);
	assign _03428_ = _02519_ | _01254_;
	assign _03429_ = _03428_ | _01490_;
	assign _03430_ = _03429_ | _01261_;
	assign _03431_ = _01243_ & ~_03430_;
	assign _03432_ = \mchip.design.owner.tokens [33] & ~_03365_;
	assign _03433_ = _03432_ | _03431_;
	assign _03434_ = _02526_ | _01281_;
	assign _03435_ = _03434_ | _01506_;
	assign _03436_ = _03435_ | _01288_;
	assign _03437_ = _01274_ & ~_03436_;
	assign _03439_ = \mchip.design.owner.tokens [33] & ~_03376_;
	assign _03440_ = _03439_ | _03437_;
	assign _03441_ = (_00199_ ? _03433_ : _03440_);
	assign _03442_ = _02534_ | _01311_;
	assign _03443_ = _03442_ | _01523_;
	assign _03444_ = _03443_ | _01318_;
	assign _03445_ = _01303_ & ~_03444_;
	assign _03446_ = \mchip.design.owner.tokens [33] & ~_03388_;
	assign _03447_ = _03446_ | _03445_;
	assign _03448_ = (_00131_ ? _03441_ : _03447_);
	assign _03450_ = _02542_ | _01341_;
	assign _03451_ = _03450_ | _01540_;
	assign _03452_ = _03451_ | _01346_;
	assign _03453_ = _01349_ & ~_03452_;
	assign _03454_ = \mchip.design.owner.tokens [33] & ~_03400_;
	assign _03455_ = _03454_ | _03453_;
	assign _03456_ = (_06005_ ? _03448_ : _03455_);
	assign _03457_ = _02550_ | _01374_;
	assign _03458_ = _03457_ | ~_01377_;
	assign _03459_ = _03458_ | _01380_;
	assign _03461_ = _01382_ & ~_03459_;
	assign _03462_ = \mchip.design.owner.tokens [33] & ~_03412_;
	assign _03463_ = _03462_ | _03461_;
	assign _03464_ = (_05934_ ? _03456_ : _03463_);
	assign _03465_ = _02558_ | _01404_;
	assign _03466_ = _03465_ | _01575_;
	assign _03467_ = _03466_ | _01398_;
	assign _03468_ = _01410_ & ~_03467_;
	assign _03469_ = \mchip.design.owner.tokens [33] & ~_03424_;
	assign _03470_ = _03469_ | _03468_;
	assign _00038_ = (_05827_ ? _03464_ : _03470_);
	assign _03472_ = _01495_ | _01257_;
	assign _03473_ = _03472_ | _01261_;
	assign _03474_ = _01243_ & ~_03473_;
	assign _03475_ = _01500_ | _01257_;
	assign _03476_ = _03475_ | _01261_;
	assign _03477_ = _01243_ & ~_03476_;
	assign _03478_ = \mchip.design.owner.tokens [34] & ~_03477_;
	assign _03479_ = _03478_ | _03474_;
	assign _03480_ = _01511_ | _01284_;
	assign _03482_ = _03480_ | _01288_;
	assign _03483_ = _01274_ & ~_03482_;
	assign _03484_ = _01516_ | _01284_;
	assign _03485_ = _03484_ | _01288_;
	assign _03486_ = _01274_ & ~_03485_;
	assign _03487_ = \mchip.design.owner.tokens [34] & ~_03486_;
	assign _03488_ = _03487_ | _03483_;
	assign _03489_ = (_00199_ ? _03479_ : _03488_);
	assign _03490_ = _01528_ | _01314_;
	assign _03491_ = _03490_ | _01318_;
	assign _03493_ = _01303_ & ~_03491_;
	assign _03494_ = _01533_ | _01314_;
	assign _03495_ = _03494_ | _01318_;
	assign _03496_ = _01303_ & ~_03495_;
	assign _03497_ = \mchip.design.owner.tokens [34] & ~_03496_;
	assign _03498_ = _03497_ | _03493_;
	assign _03499_ = (_00131_ ? _03489_ : _03498_);
	assign _03500_ = _01546_ | _01343_;
	assign _03501_ = _03500_ | _01346_;
	assign _03502_ = _01349_ & ~_03501_;
	assign _03504_ = _01551_ | _01343_;
	assign _03505_ = _03504_ | _01346_;
	assign _03506_ = _01349_ & ~_03505_;
	assign _03507_ = \mchip.design.owner.tokens [34] & ~_03506_;
	assign _03508_ = _03507_ | _03502_;
	assign _03509_ = (_06005_ ? _03499_ : _03508_);
	assign _03510_ = _01563_ | _01377_;
	assign _03511_ = _03510_ | _01380_;
	assign _03512_ = _01382_ & ~_03511_;
	assign _03513_ = _01568_ | _01377_;
	assign _03515_ = _03513_ | _01380_;
	assign _03516_ = _01382_ & ~_03515_;
	assign _03517_ = \mchip.design.owner.tokens [34] & ~_03516_;
	assign _03518_ = _03517_ | _03512_;
	assign _03519_ = (_05934_ ? _03509_ : _03518_);
	assign _03520_ = _01580_ | _01407_;
	assign _03521_ = _03520_ | _01398_;
	assign _03522_ = _01410_ & ~_03521_;
	assign _03523_ = _01587_ | _01407_;
	assign _03524_ = _03523_ | _01398_;
	assign _03526_ = _01410_ & ~_03524_;
	assign _03527_ = \mchip.design.owner.tokens [34] & ~_03526_;
	assign _03528_ = _03527_ | _03522_;
	assign _00039_ = (_05827_ ? _03519_ : _03528_);
	assign _03529_ = _01597_ | _01257_;
	assign _03530_ = _03529_ | _01261_;
	assign _03531_ = _01243_ & ~_03530_;
	assign _03532_ = \mchip.design.owner.tokens [35] & ~_03477_;
	assign _03533_ = _03532_ | _03531_;
	assign _03534_ = _01607_ | _01284_;
	assign _03536_ = _03534_ | _01288_;
	assign _03537_ = _01274_ & ~_03536_;
	assign _03538_ = \mchip.design.owner.tokens [35] & ~_03486_;
	assign _03539_ = _03538_ | _03537_;
	assign _03540_ = (_00199_ ? _03533_ : _03539_);
	assign _03541_ = _01618_ | _01314_;
	assign _03542_ = _03541_ | _01318_;
	assign _03543_ = _01303_ & ~_03542_;
	assign _03544_ = \mchip.design.owner.tokens [35] & ~_03496_;
	assign _03545_ = _03544_ | _03543_;
	assign _03547_ = (_00131_ ? _03540_ : _03545_);
	assign _03548_ = _01629_ | _01343_;
	assign _03549_ = _03548_ | _01346_;
	assign _03550_ = _01349_ & ~_03549_;
	assign _03551_ = \mchip.design.owner.tokens [35] & ~_03506_;
	assign _03552_ = _03551_ | _03550_;
	assign _03553_ = (_06005_ ? _03547_ : _03552_);
	assign _03554_ = _01640_ | _01377_;
	assign _03555_ = _03554_ | _01380_;
	assign _03556_ = _01382_ & ~_03555_;
	assign _03558_ = \mchip.design.owner.tokens [35] & ~_03516_;
	assign _03559_ = _03558_ | _03556_;
	assign _03560_ = (_05934_ ? _03553_ : _03559_);
	assign _03561_ = _01651_ | _01407_;
	assign _03562_ = _03561_ | _01398_;
	assign _03563_ = _01410_ & ~_03562_;
	assign _03564_ = \mchip.design.owner.tokens [35] & ~_03526_;
	assign _03565_ = _03564_ | _03563_;
	assign _00040_ = (_05827_ ? _03560_ : _03565_);
	assign _03566_ = _01660_ | _01257_;
	assign _03568_ = _03566_ | _01261_;
	assign _03569_ = _01243_ & ~_03568_;
	assign _03570_ = _01665_ | _01257_;
	assign _03571_ = _03570_ | _01261_;
	assign _03572_ = _01243_ & ~_03571_;
	assign _03573_ = \mchip.design.owner.tokens [36] & ~_03572_;
	assign _03574_ = _03573_ | _03569_;
	assign _03575_ = _01674_ | _01284_;
	assign _03576_ = _03575_ | _01288_;
	assign _03577_ = _01274_ & ~_03576_;
	assign _03579_ = _01679_ | _01284_;
	assign _03580_ = _03579_ | _01288_;
	assign _03581_ = _01274_ & ~_03580_;
	assign _03582_ = \mchip.design.owner.tokens [36] & ~_03581_;
	assign _03583_ = _03582_ | _03577_;
	assign _03584_ = (_00199_ ? _03574_ : _03583_);
	assign _03585_ = _01689_ | _01314_;
	assign _03586_ = _03585_ | _01318_;
	assign _03587_ = _01303_ & ~_03586_;
	assign _03588_ = _01694_ | _01314_;
	assign _03590_ = _03588_ | _01318_;
	assign _03591_ = _01303_ & ~_03590_;
	assign _03592_ = \mchip.design.owner.tokens [36] & ~_03591_;
	assign _03593_ = _03592_ | _03587_;
	assign _03594_ = (_00131_ ? _03584_ : _03593_);
	assign _03595_ = _01704_ | _01343_;
	assign _03596_ = _03595_ | _01346_;
	assign _03597_ = _01349_ & ~_03596_;
	assign _03598_ = _01709_ | _01343_;
	assign _03599_ = _03598_ | _01346_;
	assign _03601_ = _01349_ & ~_03599_;
	assign _03602_ = \mchip.design.owner.tokens [36] & ~_03601_;
	assign _03603_ = _03602_ | _03597_;
	assign _03604_ = (_06005_ ? _03594_ : _03603_);
	assign _03605_ = _01719_ | _01377_;
	assign _03606_ = _03605_ | _01380_;
	assign _03607_ = _01382_ & ~_03606_;
	assign _03608_ = _01727_ | _01377_;
	assign _03609_ = _03608_ | _01380_;
	assign _03610_ = _01382_ & ~_03609_;
	assign _03612_ = \mchip.design.owner.tokens [36] & ~_03610_;
	assign _03613_ = _03612_ | _03607_;
	assign _03614_ = (_05934_ ? _03604_ : _03613_);
	assign _03615_ = _01737_ | _01407_;
	assign _03616_ = _03615_ | _01398_;
	assign _03617_ = _01410_ & ~_03616_;
	assign _03618_ = _01744_ | _01407_;
	assign _03619_ = _03618_ | _01398_;
	assign _03620_ = _01410_ & ~_03619_;
	assign _03621_ = \mchip.design.owner.tokens [36] & ~_03620_;
	assign _03623_ = _03621_ | _03617_;
	assign _00041_ = (_05827_ ? _03614_ : _03623_);
	assign _03624_ = _01753_ | _01257_;
	assign _03625_ = _03624_ | _01261_;
	assign _03626_ = _01243_ & ~_03625_;
	assign _03627_ = \mchip.design.owner.tokens [37] & ~_03572_;
	assign _03628_ = _03627_ | _03626_;
	assign _03629_ = _01762_ | _01284_;
	assign _03630_ = _03629_ | _01288_;
	assign _03631_ = _01274_ & ~_03630_;
	assign _03633_ = \mchip.design.owner.tokens [37] & ~_03581_;
	assign _03634_ = _03633_ | _03631_;
	assign _03635_ = (_00199_ ? _03628_ : _03634_);
	assign _03636_ = _01772_ | _01314_;
	assign _03637_ = _03636_ | _01318_;
	assign _03638_ = _01303_ & ~_03637_;
	assign _03639_ = \mchip.design.owner.tokens [37] & ~_03591_;
	assign _03640_ = _03639_ | _03638_;
	assign _03641_ = (_00131_ ? _03635_ : _03640_);
	assign _03642_ = _01782_ | _01343_;
	assign _03644_ = _03642_ | _01346_;
	assign _03645_ = _01349_ & ~_03644_;
	assign _03646_ = \mchip.design.owner.tokens [37] & ~_03601_;
	assign _03647_ = _03646_ | _03645_;
	assign _03648_ = (_06005_ ? _03641_ : _03647_);
	assign _03649_ = _01792_ | _01377_;
	assign _03650_ = _03649_ | _01380_;
	assign _03651_ = _01382_ & ~_03650_;
	assign _03652_ = \mchip.design.owner.tokens [37] & ~_03610_;
	assign _03653_ = _03652_ | _03651_;
	assign _03655_ = (_05934_ ? _03648_ : _03653_);
	assign _03656_ = _01802_ | _01407_;
	assign _03657_ = _03656_ | _01398_;
	assign _03658_ = _01410_ & ~_03657_;
	assign _03659_ = \mchip.design.owner.tokens [37] & ~_03620_;
	assign _03660_ = _03659_ | _03658_;
	assign _00042_ = (_05827_ ? _03655_ : _03660_);
	assign _03661_ = _01810_ | _01257_;
	assign _03662_ = _03661_ | _01261_;
	assign _03663_ = _01243_ & ~_03662_;
	assign _03665_ = _01815_ | _01257_;
	assign _03666_ = _03665_ | _01261_;
	assign _03667_ = _01243_ & ~_03666_;
	assign _03668_ = \mchip.design.owner.tokens [38] & ~_03667_;
	assign _03669_ = _03668_ | _03663_;
	assign _03670_ = _01823_ | _01284_;
	assign _03671_ = _03670_ | _01288_;
	assign _03672_ = _01274_ & ~_03671_;
	assign _03673_ = _01828_ | _01284_;
	assign _03674_ = _03673_ | _01288_;
	assign _03676_ = _01274_ & ~_03674_;
	assign _03677_ = \mchip.design.owner.tokens [38] & ~_03676_;
	assign _03678_ = _03677_ | _03672_;
	assign _03679_ = (_00199_ ? _03669_ : _03678_);
	assign _03680_ = _01837_ | _01314_;
	assign _03681_ = _03680_ | _01318_;
	assign _03682_ = _01303_ & ~_03681_;
	assign _03683_ = _01842_ | _01314_;
	assign _03684_ = _03683_ | _01318_;
	assign _03685_ = _01303_ & ~_03684_;
	assign _03687_ = \mchip.design.owner.tokens [38] & ~_03685_;
	assign _03688_ = _03687_ | _03682_;
	assign _03689_ = (_00131_ ? _03679_ : _03688_);
	assign _03690_ = _01851_ | _01343_;
	assign _03691_ = _03690_ | _01346_;
	assign _03692_ = _01349_ & ~_03691_;
	assign _03693_ = _01856_ | _01343_;
	assign _03694_ = _03693_ | _01346_;
	assign _03695_ = _01349_ & ~_03694_;
	assign _03696_ = \mchip.design.owner.tokens [38] & ~_03695_;
	assign _03698_ = _03696_ | _03692_;
	assign _03699_ = (_06005_ ? _03689_ : _03698_);
	assign _03700_ = _01865_ | _01377_;
	assign _03701_ = _03700_ | _01380_;
	assign _03702_ = _01382_ & ~_03701_;
	assign _03703_ = _01872_ | _01377_;
	assign _03704_ = _03703_ | _01380_;
	assign _03705_ = _01382_ & ~_03704_;
	assign _03706_ = \mchip.design.owner.tokens [38] & ~_03705_;
	assign _03707_ = _03706_ | _03702_;
	assign _03709_ = (_05934_ ? _03699_ : _03707_);
	assign _03710_ = _01881_ | _01407_;
	assign _03711_ = _03710_ | _01398_;
	assign _03712_ = _01410_ & ~_03711_;
	assign _03713_ = _01887_ | _01407_;
	assign _03714_ = _03713_ | _01398_;
	assign _03715_ = _01410_ & ~_03714_;
	assign _03716_ = \mchip.design.owner.tokens [38] & ~_03715_;
	assign _03717_ = _03716_ | _03712_;
	assign _00043_ = (_05827_ ? _03709_ : _03717_);
	assign _03719_ = _01895_ | _01257_;
	assign _03720_ = _03719_ | _01261_;
	assign _03721_ = _01243_ & ~_03720_;
	assign _03722_ = \mchip.design.owner.tokens [39] & ~_03667_;
	assign _03723_ = _03722_ | _03721_;
	assign _03724_ = _01903_ | _01284_;
	assign _03725_ = _03724_ | _01288_;
	assign _03726_ = _01274_ & ~_03725_;
	assign _03727_ = \mchip.design.owner.tokens [39] & ~_03676_;
	assign _03728_ = _03727_ | _03726_;
	assign _03730_ = (_00199_ ? _03723_ : _03728_);
	assign _03731_ = _01912_ | _01314_;
	assign _03732_ = _03731_ | _01318_;
	assign _03733_ = _01303_ & ~_03732_;
	assign _03734_ = \mchip.design.owner.tokens [39] & ~_03685_;
	assign _03735_ = _03734_ | _03733_;
	assign _03736_ = (_00131_ ? _03730_ : _03735_);
	assign _03737_ = _01921_ | _01343_;
	assign _03738_ = _03737_ | _01346_;
	assign _03739_ = _01349_ & ~_03738_;
	assign _03740_ = \mchip.design.owner.tokens [39] & ~_03695_;
	assign _03741_ = _03740_ | _03739_;
	assign _03742_ = (_06005_ ? _03736_ : _03741_);
	assign _03743_ = _01930_ | _01377_;
	assign _03744_ = _03743_ | _01380_;
	assign _03745_ = _01382_ & ~_03744_;
	assign _03746_ = \mchip.design.owner.tokens [39] & ~_03705_;
	assign _03747_ = _03746_ | _03745_;
	assign _03748_ = (_05934_ ? _03742_ : _03747_);
	assign _03749_ = _01939_ | _01407_;
	assign _03751_ = _03749_ | _01398_;
	assign _03752_ = _01410_ & ~_03751_;
	assign _03753_ = \mchip.design.owner.tokens [39] & ~_03715_;
	assign _03754_ = _03753_ | _03752_;
	assign _00044_ = (_05827_ ? _03748_ : _03754_);
	assign _03755_ = _01947_ | _01257_;
	assign _03756_ = _03755_ | _01261_;
	assign _03757_ = _01243_ & ~_03756_;
	assign _03758_ = _01952_ | _01257_;
	assign _03759_ = _03758_ | _01261_;
	assign _03761_ = _01243_ & ~_03759_;
	assign _03762_ = \mchip.design.owner.tokens [40] & ~_03761_;
	assign _03763_ = _03762_ | _03757_;
	assign _03764_ = _01960_ | _01284_;
	assign _03765_ = _03764_ | _01288_;
	assign _03766_ = _01274_ & ~_03765_;
	assign _03767_ = _01965_ | _01284_;
	assign _03768_ = _03767_ | _01288_;
	assign _03769_ = _01274_ & ~_03768_;
	assign _03770_ = \mchip.design.owner.tokens [40] & ~_03769_;
	assign _03772_ = _03770_ | _03766_;
	assign _03773_ = (_00199_ ? _03763_ : _03772_);
	assign _03774_ = _01974_ | _01314_;
	assign _03775_ = _03774_ | _01318_;
	assign _03776_ = _01303_ & ~_03775_;
	assign _03777_ = _01979_ | _01314_;
	assign _03778_ = _03777_ | _01318_;
	assign _03779_ = _01303_ & ~_03778_;
	assign _03780_ = \mchip.design.owner.tokens [40] & ~_03779_;
	assign _03781_ = _03780_ | _03776_;
	assign _03783_ = (_00131_ ? _03773_ : _03781_);
	assign _03784_ = _01988_ | _01343_;
	assign _03785_ = _03784_ | _01346_;
	assign _03786_ = _01349_ & ~_03785_;
	assign _03787_ = _01993_ | _01343_;
	assign _03788_ = _03787_ | _01346_;
	assign _03789_ = _01349_ & ~_03788_;
	assign _03790_ = \mchip.design.owner.tokens [40] & ~_03789_;
	assign _03791_ = _03790_ | _03786_;
	assign _03792_ = (_06005_ ? _03783_ : _03791_);
	assign _03794_ = _02002_ | _01377_;
	assign _03795_ = _03794_ | _01380_;
	assign _03796_ = _01382_ & ~_03795_;
	assign _03797_ = _02008_ | _01377_;
	assign _03798_ = _03797_ | _01380_;
	assign _03799_ = _01382_ & ~_03798_;
	assign _03800_ = \mchip.design.owner.tokens [40] & ~_03799_;
	assign _03801_ = _03800_ | _03796_;
	assign _03802_ = (_05934_ ? _03792_ : _03801_);
	assign _03803_ = _02017_ | _01407_;
	assign _03805_ = _03803_ | _01398_;
	assign _03806_ = _01410_ & ~_03805_;
	assign _03807_ = _02023_ | _01407_;
	assign _03808_ = _03807_ | _01398_;
	assign _03809_ = _01410_ & ~_03808_;
	assign _03810_ = \mchip.design.owner.tokens [40] & ~_03809_;
	assign _03811_ = _03810_ | _03806_;
	assign _00046_ = (_05827_ ? _03802_ : _03811_);
	assign _03812_ = _02031_ | _01257_;
	assign _03813_ = _03812_ | _01261_;
	assign _03815_ = _01243_ & ~_03813_;
	assign _03816_ = \mchip.design.owner.tokens [41] & ~_03761_;
	assign _03817_ = _03816_ | _03815_;
	assign _03818_ = _02039_ | _01284_;
	assign _03819_ = _03818_ | _01288_;
	assign _03820_ = _01274_ & ~_03819_;
	assign _03821_ = \mchip.design.owner.tokens [41] & ~_03769_;
	assign _03822_ = _03821_ | _03820_;
	assign _03823_ = (_00199_ ? _03817_ : _03822_);
	assign _03824_ = _02048_ | _01314_;
	assign _03826_ = _03824_ | _01318_;
	assign _03827_ = _01303_ & ~_03826_;
	assign _03828_ = \mchip.design.owner.tokens [41] & ~_03779_;
	assign _03829_ = _03828_ | _03827_;
	assign _03830_ = (_00131_ ? _03823_ : _03829_);
	assign _03831_ = _02057_ | _01343_;
	assign _03832_ = _03831_ | _01346_;
	assign _03833_ = _01349_ & ~_03832_;
	assign _03834_ = \mchip.design.owner.tokens [41] & ~_03789_;
	assign _03835_ = _03834_ | _03833_;
	assign _03837_ = (_06005_ ? _03830_ : _03835_);
	assign _03838_ = _02066_ | _01377_;
	assign _03839_ = _03838_ | _01380_;
	assign _03840_ = _01382_ & ~_03839_;
	assign _03841_ = \mchip.design.owner.tokens [41] & ~_03799_;
	assign _03842_ = _03841_ | _03840_;
	assign _03843_ = (_05934_ ? _03837_ : _03842_);
	assign _03844_ = _02075_ | _01407_;
	assign _03845_ = _03844_ | _01398_;
	assign _03846_ = _01410_ & ~_03845_;
	assign _03848_ = \mchip.design.owner.tokens [41] & ~_03809_;
	assign _03849_ = _03848_ | _03846_;
	assign _00047_ = (_05827_ ? _03843_ : _03849_);
	assign _03850_ = _02082_ | _01257_;
	assign _03851_ = _03850_ | _01261_;
	assign _03852_ = _01243_ & ~_03851_;
	assign _03853_ = _02087_ | _01257_;
	assign _03854_ = _03853_ | _01261_;
	assign _03855_ = _01243_ & ~_03854_;
	assign _03856_ = \mchip.design.owner.tokens [42] & ~_03855_;
	assign _03858_ = _03856_ | _03852_;
	assign _03859_ = _02094_ | _01284_;
	assign _03860_ = _03859_ | _01288_;
	assign _03861_ = _01274_ & ~_03860_;
	assign _03862_ = _02098_ | _01284_;
	assign _03863_ = _03862_ | _01288_;
	assign _03864_ = _01274_ & ~_03863_;
	assign _03865_ = \mchip.design.owner.tokens [42] & ~_03864_;
	assign _03866_ = _03865_ | _03861_;
	assign _03867_ = (_00199_ ? _03858_ : _03866_);
	assign _03869_ = _02106_ | _01314_;
	assign _03870_ = _03869_ | _01318_;
	assign _03871_ = _01303_ & ~_03870_;
	assign _03872_ = _02110_ | _01314_;
	assign _03873_ = _03872_ | _01318_;
	assign _03874_ = _01303_ & ~_03873_;
	assign _03875_ = \mchip.design.owner.tokens [42] & ~_03874_;
	assign _03876_ = _03875_ | _03871_;
	assign _03877_ = (_00131_ ? _03867_ : _03876_);
	assign _03878_ = _02118_ | _01343_;
	assign _03880_ = _03878_ | _01346_;
	assign _03881_ = _01349_ & ~_03880_;
	assign _03882_ = _02123_ | _01343_;
	assign _03883_ = _03882_ | _01346_;
	assign _03884_ = _01349_ & ~_03883_;
	assign _03885_ = \mchip.design.owner.tokens [42] & ~_03884_;
	assign _03886_ = _03885_ | _03881_;
	assign _03887_ = (_06005_ ? _03877_ : _03886_);
	assign _03888_ = _02131_ | _01377_;
	assign _03889_ = _03888_ | _01380_;
	assign _03891_ = _01382_ & ~_03889_;
	assign _03892_ = _02136_ | _01377_;
	assign _03893_ = _03892_ | _01380_;
	assign _03894_ = _01382_ & ~_03893_;
	assign _03895_ = \mchip.design.owner.tokens [42] & ~_03894_;
	assign _03896_ = _03895_ | _03891_;
	assign _03897_ = (_05934_ ? _03887_ : _03896_);
	assign _03898_ = _02144_ | _01407_;
	assign _03899_ = _03898_ | _01398_;
	assign _03900_ = _01410_ & ~_03899_;
	assign _03902_ = _02149_ | _01407_;
	assign _03903_ = _03902_ | _01398_;
	assign _03904_ = _01410_ & ~_03903_;
	assign _03905_ = \mchip.design.owner.tokens [42] & ~_03904_;
	assign _03906_ = _03905_ | _03900_;
	assign _00048_ = (_05827_ ? _03897_ : _03906_);
	assign _03907_ = _02156_ | _01257_;
	assign _03908_ = _03907_ | _01261_;
	assign _03909_ = _01243_ & ~_03908_;
	assign _03910_ = \mchip.design.owner.tokens [43] & ~_03855_;
	assign _03912_ = _03910_ | _03909_;
	assign _03913_ = _02163_ | _01284_;
	assign _03914_ = _03913_ | _01288_;
	assign _03915_ = _01274_ & ~_03914_;
	assign _03916_ = \mchip.design.owner.tokens [43] & ~_03864_;
	assign _03917_ = _03916_ | _03915_;
	assign _03918_ = (_00199_ ? _03912_ : _03917_);
	assign _03919_ = _02171_ | _01314_;
	assign _03920_ = _03919_ | _01318_;
	assign _03921_ = _01303_ & ~_03920_;
	assign _03923_ = \mchip.design.owner.tokens [43] & ~_03874_;
	assign _03924_ = _03923_ | _03921_;
	assign _03925_ = (_00131_ ? _03918_ : _03924_);
	assign _03926_ = _02179_ | _01343_;
	assign _03927_ = _03926_ | _01346_;
	assign _03928_ = _01349_ & ~_03927_;
	assign _03929_ = \mchip.design.owner.tokens [43] & ~_03884_;
	assign _03930_ = _03929_ | _03928_;
	assign _03931_ = (_06005_ ? _03925_ : _03930_);
	assign _03932_ = _02187_ | _01377_;
	assign _03933_ = _03932_ | _01380_;
	assign _03934_ = _01382_ & ~_03933_;
	assign _03935_ = \mchip.design.owner.tokens [43] & ~_03894_;
	assign _03936_ = _03935_ | _03934_;
	assign _03937_ = (_05934_ ? _03931_ : _03936_);
	assign _03938_ = _02195_ | _01407_;
	assign _03939_ = _03938_ | _01398_;
	assign _03940_ = _01410_ & ~_03939_;
	assign _03941_ = \mchip.design.owner.tokens [43] & ~_03904_;
	assign _03942_ = _03941_ | _03940_;
	assign _00049_ = (_05827_ ? _03937_ : _03942_);
	assign _03943_ = _02202_ | _01257_;
	assign _03944_ = _03943_ | _01261_;
	assign _03945_ = _01243_ & ~_03944_;
	assign _03946_ = _02207_ | _01257_;
	assign _03947_ = _03946_ | _01261_;
	assign _03948_ = _01243_ & ~_03947_;
	assign _03949_ = \mchip.design.owner.tokens [44] & ~_03948_;
	assign _03950_ = _03949_ | _03945_;
	assign _03951_ = _02214_ | _01284_;
	assign _03952_ = _03951_ | _01288_;
	assign _03953_ = _01274_ & ~_03952_;
	assign _03954_ = _02219_ | _01284_;
	assign _03955_ = _03954_ | _01288_;
	assign _03956_ = _01274_ & ~_03955_;
	assign _03957_ = \mchip.design.owner.tokens [44] & ~_03956_;
	assign _03958_ = _03957_ | _03953_;
	assign _03959_ = (_00199_ ? _03950_ : _03958_);
	assign _03960_ = _02227_ | _01314_;
	assign _03961_ = _03960_ | _01318_;
	assign _03962_ = _01303_ & ~_03961_;
	assign _03963_ = _02232_ | _01314_;
	assign _03964_ = _03963_ | _01318_;
	assign _03965_ = _01303_ & ~_03964_;
	assign _03966_ = \mchip.design.owner.tokens [44] & ~_03965_;
	assign _03967_ = _03966_ | _03962_;
	assign _03968_ = (_00131_ ? _03959_ : _03967_);
	assign _03969_ = _02240_ | _01343_;
	assign _03970_ = _03969_ | _01346_;
	assign _03971_ = _01349_ & ~_03970_;
	assign _03972_ = _02245_ | _01343_;
	assign _03973_ = _03972_ | _01346_;
	assign _03974_ = _01349_ & ~_03973_;
	assign _03975_ = \mchip.design.owner.tokens [44] & ~_03974_;
	assign _03976_ = _03975_ | _03971_;
	assign _03977_ = (_06005_ ? _03968_ : _03976_);
	assign _03978_ = _02253_ | _01377_;
	assign _03979_ = _03978_ | _01380_;
	assign _03980_ = _01382_ & ~_03979_;
	assign _03981_ = _02258_ | _01377_;
	assign _03982_ = _03981_ | _01380_;
	assign _03983_ = _01382_ & ~_03982_;
	assign _03984_ = \mchip.design.owner.tokens [44] & ~_03983_;
	assign _03985_ = _03984_ | _03980_;
	assign _03986_ = (_05934_ ? _03977_ : _03985_);
	assign _03987_ = _02266_ | _01407_;
	assign _03988_ = _03987_ | _01398_;
	assign _03989_ = _01410_ & ~_03988_;
	assign _03990_ = _02271_ | _01407_;
	assign _03991_ = _03990_ | _01398_;
	assign _03993_ = _01410_ & ~_03991_;
	assign _03994_ = \mchip.design.owner.tokens [44] & ~_03993_;
	assign _03995_ = _03994_ | _03989_;
	assign _00050_ = (_05827_ ? _03986_ : _03995_);
	assign _03996_ = _02278_ | _01257_;
	assign _03997_ = _03996_ | _01261_;
	assign _03998_ = _01243_ & ~_03997_;
	assign _03999_ = \mchip.design.owner.tokens [45] & ~_03948_;
	assign _04000_ = _03999_ | _03998_;
	assign _04001_ = _02285_ | _01284_;
	assign _04003_ = _04001_ | _01288_;
	assign _04004_ = _01274_ & ~_04003_;
	assign _04005_ = \mchip.design.owner.tokens [45] & ~_03956_;
	assign _04006_ = _04005_ | _04004_;
	assign _04007_ = (_00199_ ? _04000_ : _04006_);
	assign _04008_ = _02293_ | _01314_;
	assign _04009_ = _04008_ | _01318_;
	assign _04010_ = _01303_ & ~_04009_;
	assign _04011_ = \mchip.design.owner.tokens [45] & ~_03965_;
	assign _04012_ = _04011_ | _04010_;
	assign _04014_ = (_00131_ ? _04007_ : _04012_);
	assign _04015_ = _02301_ | _01343_;
	assign _04016_ = _04015_ | _01346_;
	assign _04017_ = _01349_ & ~_04016_;
	assign _04018_ = \mchip.design.owner.tokens [45] & ~_03974_;
	assign _04019_ = _04018_ | _04017_;
	assign _04020_ = (_06005_ ? _04014_ : _04019_);
	assign _04021_ = _02309_ | _01377_;
	assign _04022_ = _04021_ | _01380_;
	assign _04023_ = _01382_ & ~_04022_;
	assign _04025_ = \mchip.design.owner.tokens [45] & ~_03983_;
	assign _04026_ = _04025_ | _04023_;
	assign _04027_ = (_05934_ ? _04020_ : _04026_);
	assign _04028_ = _02317_ | _01407_;
	assign _04029_ = _04028_ | _01398_;
	assign _04030_ = _01410_ & ~_04029_;
	assign _04031_ = \mchip.design.owner.tokens [45] & ~_03993_;
	assign _04032_ = _04031_ | _04030_;
	assign _00051_ = (_05827_ ? _04027_ : _04032_);
	assign _04033_ = _02324_ | _01257_;
	assign _04035_ = _04033_ | _01261_;
	assign _04036_ = _01243_ & ~_04035_;
	assign _04037_ = _02329_ | _01257_;
	assign _04038_ = _04037_ | _01261_;
	assign _04039_ = _01243_ & ~_04038_;
	assign _04040_ = \mchip.design.owner.tokens [46] & ~_04039_;
	assign _04041_ = _04040_ | _04036_;
	assign _04042_ = _02336_ | _01284_;
	assign _04043_ = _04042_ | _01288_;
	assign _04044_ = _01274_ & ~_04043_;
	assign _04046_ = _02341_ | _01284_;
	assign _04047_ = _04046_ | _01288_;
	assign _04048_ = _01274_ & ~_04047_;
	assign _04049_ = \mchip.design.owner.tokens [46] & ~_04048_;
	assign _04050_ = _04049_ | _04044_;
	assign _04051_ = (_00199_ ? _04041_ : _04050_);
	assign _04052_ = _02349_ | _01314_;
	assign _04053_ = _04052_ | _01318_;
	assign _04054_ = _01303_ & ~_04053_;
	assign _04055_ = _02354_ | _01314_;
	assign _04057_ = _04055_ | _01318_;
	assign _04058_ = _01303_ & ~_04057_;
	assign _04059_ = \mchip.design.owner.tokens [46] & ~_04058_;
	assign _04060_ = _04059_ | _04054_;
	assign _04061_ = (_00131_ ? _04051_ : _04060_);
	assign _04062_ = _02362_ | _01343_;
	assign _04063_ = _04062_ | _01346_;
	assign _04064_ = _01349_ & ~_04063_;
	assign _04065_ = _02367_ | _01343_;
	assign _04066_ = _04065_ | _01346_;
	assign _04068_ = _01349_ & ~_04066_;
	assign _04069_ = \mchip.design.owner.tokens [46] & ~_04068_;
	assign _04070_ = _04069_ | _04064_;
	assign _04071_ = (_06005_ ? _04061_ : _04070_);
	assign _04072_ = _02375_ | _01377_;
	assign _04073_ = _04072_ | _01380_;
	assign _04074_ = _01382_ & ~_04073_;
	assign _04075_ = _02380_ | _01377_;
	assign _04076_ = _04075_ | _01380_;
	assign _04077_ = _01382_ & ~_04076_;
	assign _04079_ = \mchip.design.owner.tokens [46] & ~_04077_;
	assign _04080_ = _04079_ | _04074_;
	assign _04081_ = (_05934_ ? _04071_ : _04080_);
	assign _04082_ = _02388_ | _01407_;
	assign _04083_ = _04082_ | _01398_;
	assign _04084_ = _01410_ & ~_04083_;
	assign _04085_ = _02393_ | _01407_;
	assign _04086_ = _04085_ | _01398_;
	assign _04087_ = _01410_ & ~_04086_;
	assign _04088_ = \mchip.design.owner.tokens [46] & ~_04087_;
	assign _04090_ = _04088_ | _04084_;
	assign _00052_ = (_05827_ ? _04081_ : _04090_);
	assign _04091_ = _02400_ | _01257_;
	assign _04092_ = _04091_ | _01261_;
	assign _04093_ = _01243_ & ~_04092_;
	assign _04094_ = \mchip.design.owner.tokens [47] & ~_04039_;
	assign _04095_ = _04094_ | _04093_;
	assign _04096_ = _02407_ | _01284_;
	assign _04097_ = _04096_ | _01288_;
	assign _04098_ = _01274_ & ~_04097_;
	assign _04100_ = \mchip.design.owner.tokens [47] & ~_04048_;
	assign _04101_ = _04100_ | _04098_;
	assign _04102_ = (_00199_ ? _04095_ : _04101_);
	assign _04103_ = _02415_ | _01314_;
	assign _04104_ = _04103_ | _01318_;
	assign _04105_ = _01303_ & ~_04104_;
	assign _04106_ = \mchip.design.owner.tokens [47] & ~_04058_;
	assign _04107_ = _04106_ | _04105_;
	assign _04108_ = (_00131_ ? _04102_ : _04107_);
	assign _04109_ = _02423_ | _01343_;
	assign _04111_ = _04109_ | _01346_;
	assign _04112_ = _01349_ & ~_04111_;
	assign _04113_ = \mchip.design.owner.tokens [47] & ~_04068_;
	assign _04114_ = _04113_ | _04112_;
	assign _04115_ = (_06005_ ? _04108_ : _04114_);
	assign _04116_ = _02431_ | _01377_;
	assign _04117_ = _04116_ | _01380_;
	assign _04118_ = _01382_ & ~_04117_;
	assign _04119_ = \mchip.design.owner.tokens [47] & ~_04077_;
	assign _04120_ = _04119_ | _04118_;
	assign _04122_ = (_05934_ ? _04115_ : _04120_);
	assign _04123_ = _02439_ | _01407_;
	assign _04124_ = _04123_ | _01398_;
	assign _04125_ = _01410_ & ~_04124_;
	assign _04126_ = \mchip.design.owner.tokens [47] & ~_04087_;
	assign _04127_ = _04126_ | _04125_;
	assign _00053_ = (_05827_ ? _04122_ : _04127_);
	assign _04128_ = _02446_ | _01257_;
	assign _04129_ = _04128_ | _01261_;
	assign _04130_ = _01243_ & ~_04129_;
	assign _04132_ = _02450_ | _01257_;
	assign _04133_ = _04132_ | _01261_;
	assign _04134_ = _01243_ & ~_04133_;
	assign _04135_ = \mchip.design.owner.tokens [48] & ~_04134_;
	assign _04136_ = _04135_ | _04130_;
	assign _04137_ = _02457_ | _01284_;
	assign _04138_ = _04137_ | _01288_;
	assign _04139_ = _01274_ & ~_04138_;
	assign _04140_ = _02461_ | _01284_;
	assign _04141_ = _04140_ | _01288_;
	assign _04143_ = _01274_ & ~_04141_;
	assign _04144_ = \mchip.design.owner.tokens [48] & ~_04143_;
	assign _04145_ = _04144_ | _04139_;
	assign _04146_ = (_00199_ ? _04136_ : _04145_);
	assign _04147_ = _02469_ | _01314_;
	assign _04148_ = _04147_ | _01318_;
	assign _04149_ = _01303_ & ~_04148_;
	assign _04150_ = _02474_ | _01314_;
	assign _04151_ = _04150_ | _01318_;
	assign _04152_ = _01303_ & ~_04151_;
	assign _04154_ = \mchip.design.owner.tokens [48] & ~_04152_;
	assign _04155_ = _04154_ | _04149_;
	assign _04156_ = (_00131_ ? _04146_ : _04155_);
	assign _04157_ = _02482_ | _01343_;
	assign _04158_ = _04157_ | _01346_;
	assign _04159_ = _01349_ & ~_04158_;
	assign _04160_ = _02487_ | _01343_;
	assign _04161_ = _04160_ | _01346_;
	assign _04162_ = _01349_ & ~_04161_;
	assign _04163_ = \mchip.design.owner.tokens [48] & ~_04162_;
	assign _04165_ = _04163_ | _04159_;
	assign _04166_ = (_06005_ ? _04156_ : _04165_);
	assign _04167_ = _02495_ | _01377_;
	assign _04168_ = _04167_ | _01380_;
	assign _04169_ = _01382_ & ~_04168_;
	assign _04170_ = _02500_ | _01377_;
	assign _04171_ = _04170_ | _01380_;
	assign _04172_ = _01382_ & ~_04171_;
	assign _04173_ = \mchip.design.owner.tokens [48] & ~_04172_;
	assign _04174_ = _04173_ | _04169_;
	assign _04176_ = (_05934_ ? _04166_ : _04174_);
	assign _04177_ = _02508_ | _01407_;
	assign _04178_ = _04177_ | _01398_;
	assign _04179_ = _01410_ & ~_04178_;
	assign _04180_ = _02513_ | _01407_;
	assign _04181_ = _04180_ | _01398_;
	assign _04182_ = _01410_ & ~_04181_;
	assign _04183_ = \mchip.design.owner.tokens [48] & ~_04182_;
	assign _04184_ = _04183_ | _04179_;
	assign _00054_ = (_05827_ ? _04176_ : _04184_);
	assign _04186_ = _02520_ | _01257_;
	assign _04187_ = _04186_ | _01261_;
	assign _04188_ = _01243_ & ~_04187_;
	assign _04189_ = \mchip.design.owner.tokens [49] & ~_04134_;
	assign _04190_ = _04189_ | _04188_;
	assign _04191_ = _02527_ | _01284_;
	assign _04192_ = _04191_ | _01288_;
	assign _04193_ = _01274_ & ~_04192_;
	assign _04194_ = \mchip.design.owner.tokens [49] & ~_04143_;
	assign _04195_ = _04194_ | _04193_;
	assign _04197_ = (_00199_ ? _04190_ : _04195_);
	assign _04198_ = _02535_ | _01314_;
	assign _04199_ = _04198_ | _01318_;
	assign _04200_ = _01303_ & ~_04199_;
	assign _04201_ = \mchip.design.owner.tokens [49] & ~_04152_;
	assign _04202_ = _04201_ | _04200_;
	assign _04203_ = (_00131_ ? _04197_ : _04202_);
	assign _04204_ = _02543_ | _01343_;
	assign _04205_ = _04204_ | _01346_;
	assign _04206_ = _01349_ & ~_04205_;
	assign _04208_ = \mchip.design.owner.tokens [49] & ~_04162_;
	assign _04209_ = _04208_ | _04206_;
	assign _04210_ = (_06005_ ? _04203_ : _04209_);
	assign _04211_ = _02551_ | _01377_;
	assign _04212_ = _04211_ | _01380_;
	assign _04213_ = _01382_ & ~_04212_;
	assign _04214_ = \mchip.design.owner.tokens [49] & ~_04172_;
	assign _04215_ = _04214_ | _04213_;
	assign _04216_ = (_05934_ ? _04210_ : _04215_);
	assign _04217_ = _02559_ | _01407_;
	assign _04219_ = _04217_ | _01398_;
	assign _04220_ = _01410_ & ~_04219_;
	assign _04221_ = \mchip.design.owner.tokens [49] & ~_04182_;
	assign _04222_ = _04221_ | _04220_;
	assign _00055_ = (_05827_ ? _04216_ : _04222_);
	assign _04223_ = _02565_ | _01257_;
	assign _04224_ = _04223_ | _01261_;
	assign _04225_ = _01243_ & ~_04224_;
	assign _04226_ = _02569_ | _01257_;
	assign _04227_ = _04226_ | _01261_;
	assign _04229_ = _01243_ & ~_04227_;
	assign _04230_ = \mchip.design.owner.tokens [50] & ~_04229_;
	assign _04231_ = _04230_ | _04225_;
	assign _04232_ = _02575_ | _01284_;
	assign _04233_ = _04232_ | _01288_;
	assign _04234_ = _01274_ & ~_04233_;
	assign _04235_ = _02579_ | _01284_;
	assign _04236_ = _04235_ | _01288_;
	assign _04237_ = _01274_ & ~_04236_;
	assign _04238_ = \mchip.design.owner.tokens [50] & ~_04237_;
	assign _04240_ = _04238_ | _04234_;
	assign _04241_ = (_00199_ ? _04231_ : _04240_);
	assign _04242_ = _02586_ | _01314_;
	assign _04243_ = _04242_ | _01318_;
	assign _04244_ = _01303_ & ~_04243_;
	assign _04245_ = _02590_ | _01314_;
	assign _04246_ = _04245_ | _01318_;
	assign _04247_ = _01303_ & ~_04246_;
	assign _04248_ = \mchip.design.owner.tokens [50] & ~_04247_;
	assign _04249_ = _04248_ | _04244_;
	assign _04251_ = (_00131_ ? _04241_ : _04249_);
	assign _04252_ = _02597_ | _01343_;
	assign _04253_ = _04252_ | _01346_;
	assign _04254_ = _01349_ & ~_04253_;
	assign _04255_ = _02601_ | _01343_;
	assign _04256_ = _04255_ | _01346_;
	assign _04257_ = _01349_ & ~_04256_;
	assign _04258_ = \mchip.design.owner.tokens [50] & ~_04257_;
	assign _04259_ = _04258_ | _04254_;
	assign _04260_ = (_06005_ ? _04251_ : _04259_);
	assign _04262_ = _02608_ | _01377_;
	assign _04263_ = _04262_ | _01380_;
	assign _04264_ = _01382_ & ~_04263_;
	assign _04265_ = _02612_ | _01377_;
	assign _04266_ = _04265_ | _01380_;
	assign _04267_ = _01382_ & ~_04266_;
	assign _04268_ = \mchip.design.owner.tokens [50] & ~_04267_;
	assign _04269_ = _04268_ | _04264_;
	assign _04270_ = (_05934_ ? _04260_ : _04269_);
	assign _04271_ = _02619_ | _01407_;
	assign _04273_ = _04271_ | _01398_;
	assign _04274_ = _01410_ & ~_04273_;
	assign _04275_ = _02623_ | _01407_;
	assign _04276_ = _04275_ | _01398_;
	assign _04277_ = _01410_ & ~_04276_;
	assign _04278_ = \mchip.design.owner.tokens [50] & ~_04277_;
	assign _04279_ = _04278_ | _04274_;
	assign _00057_ = (_05827_ ? _04270_ : _04279_);
	assign _04280_ = _02629_ | _01257_;
	assign _04281_ = _04280_ | _01261_;
	assign _04283_ = _01243_ & ~_04281_;
	assign _04284_ = \mchip.design.owner.tokens [51] & ~_04229_;
	assign _04285_ = _04284_ | _04283_;
	assign _04286_ = _02635_ | _01284_;
	assign _04287_ = _04286_ | _01288_;
	assign _04288_ = _01274_ & ~_04287_;
	assign _04289_ = \mchip.design.owner.tokens [51] & ~_04237_;
	assign _04290_ = _04289_ | _04288_;
	assign _04291_ = (_00199_ ? _04285_ : _04290_);
	assign _04292_ = _02642_ | _01314_;
	assign _04294_ = _04292_ | _01318_;
	assign _04295_ = _01303_ & ~_04294_;
	assign _04296_ = \mchip.design.owner.tokens [51] & ~_04247_;
	assign _04297_ = _04296_ | _04295_;
	assign _04298_ = (_00131_ ? _04291_ : _04297_);
	assign _04299_ = _02649_ | _01343_;
	assign _04300_ = _04299_ | _01346_;
	assign _04301_ = _01349_ & ~_04300_;
	assign _04302_ = \mchip.design.owner.tokens [51] & ~_04257_;
	assign _04303_ = _04302_ | _04301_;
	assign _04305_ = (_06005_ ? _04298_ : _04303_);
	assign _04306_ = _02656_ | _01377_;
	assign _04307_ = _04306_ | _01380_;
	assign _04308_ = _01382_ & ~_04307_;
	assign _04309_ = \mchip.design.owner.tokens [51] & ~_04267_;
	assign _04310_ = _04309_ | _04308_;
	assign _04311_ = (_05934_ ? _04305_ : _04310_);
	assign _04312_ = _02664_ | _01407_;
	assign _04313_ = _04312_ | _01398_;
	assign _04314_ = _01410_ & ~_04313_;
	assign _04316_ = \mchip.design.owner.tokens [51] & ~_04277_;
	assign _04317_ = _04316_ | _04314_;
	assign _00058_ = (_05827_ ? _04311_ : _04317_);
	assign _04318_ = _02670_ | _01257_;
	assign _04319_ = _04318_ | _01261_;
	assign _04320_ = _01243_ & ~_04319_;
	assign _04321_ = _02675_ | _01257_;
	assign _04322_ = _04321_ | _01261_;
	assign _04323_ = _01243_ & ~_04322_;
	assign _04324_ = \mchip.design.owner.tokens [52] & ~_04323_;
	assign _04326_ = _04324_ | _04320_;
	assign _04327_ = _02681_ | _01284_;
	assign _04328_ = _04327_ | _01288_;
	assign _04329_ = _01274_ & ~_04328_;
	assign _04330_ = _02686_ | _01284_;
	assign _04331_ = _04330_ | _01288_;
	assign _04332_ = _01274_ & ~_04331_;
	assign _04333_ = \mchip.design.owner.tokens [52] & ~_04332_;
	assign _04334_ = _04333_ | _04329_;
	assign _04335_ = (_00199_ ? _04326_ : _04334_);
	assign _04337_ = _02694_ | _01314_;
	assign _04338_ = _04337_ | _01318_;
	assign _04339_ = _01303_ & ~_04338_;
	assign _04340_ = _02698_ | _01314_;
	assign _04341_ = _04340_ | _01318_;
	assign _04342_ = _01303_ & ~_04341_;
	assign _04343_ = \mchip.design.owner.tokens [52] & ~_04342_;
	assign _04344_ = _04343_ | _04339_;
	assign _04345_ = (_00131_ ? _04335_ : _04344_);
	assign _04346_ = _02706_ | _01343_;
	assign _04348_ = _04346_ | _01346_;
	assign _04349_ = _01349_ & ~_04348_;
	assign _04350_ = _02710_ | _01343_;
	assign _04351_ = _04350_ | _01346_;
	assign _04352_ = _01349_ & ~_04351_;
	assign _04353_ = \mchip.design.owner.tokens [52] & ~_04352_;
	assign _04354_ = _04353_ | _04349_;
	assign _04355_ = (_06005_ ? _04345_ : _04354_);
	assign _04356_ = _02718_ | _01377_;
	assign _04357_ = _04356_ | _01380_;
	assign _04359_ = _01382_ & ~_04357_;
	assign _04360_ = _02722_ | _01377_;
	assign _04361_ = _04360_ | _01380_;
	assign _04362_ = _01382_ & ~_04361_;
	assign _04363_ = \mchip.design.owner.tokens [52] & ~_04362_;
	assign _04364_ = _04363_ | _04359_;
	assign _04365_ = (_05934_ ? _04355_ : _04364_);
	assign _04366_ = _02730_ | _01407_;
	assign _04367_ = _04366_ | _01398_;
	assign _04368_ = _01410_ & ~_04367_;
	assign _04370_ = _02734_ | _01407_;
	assign _04371_ = _04370_ | _01398_;
	assign _04372_ = _01410_ & ~_04371_;
	assign _04373_ = \mchip.design.owner.tokens [52] & ~_04372_;
	assign _04374_ = _04373_ | _04368_;
	assign _00059_ = (_05827_ ? _04365_ : _04374_);
	assign _04375_ = _02741_ | _01257_;
	assign _04376_ = _04375_ | _01261_;
	assign _04377_ = _01243_ & ~_04376_;
	assign _04378_ = \mchip.design.owner.tokens [53] & ~_04323_;
	assign _04380_ = _04378_ | _04377_;
	assign _04381_ = _02748_ | _01284_;
	assign _04382_ = _04381_ | _01288_;
	assign _04383_ = _01274_ & ~_04382_;
	assign _04384_ = \mchip.design.owner.tokens [53] & ~_04332_;
	assign _04385_ = _04384_ | _04383_;
	assign _04386_ = (_00199_ ? _04380_ : _04385_);
	assign _04387_ = _02755_ | _01314_;
	assign _04388_ = _04387_ | _01318_;
	assign _04389_ = _01303_ & ~_04388_;
	assign _04391_ = \mchip.design.owner.tokens [53] & ~_04342_;
	assign _04392_ = _04391_ | _04389_;
	assign _04393_ = (_00131_ ? _04386_ : _04392_);
	assign _04394_ = _02763_ | _01343_;
	assign _04395_ = _04394_ | _01346_;
	assign _04396_ = _01349_ & ~_04395_;
	assign _04397_ = \mchip.design.owner.tokens [53] & ~_04352_;
	assign _04398_ = _04397_ | _04396_;
	assign _04399_ = (_06005_ ? _04393_ : _04398_);
	assign _04400_ = _02771_ | _01377_;
	assign _04402_ = _04400_ | _01380_;
	assign _04403_ = _01382_ & ~_04402_;
	assign _04404_ = \mchip.design.owner.tokens [53] & ~_04362_;
	assign _04405_ = _04404_ | _04403_;
	assign _04406_ = (_05934_ ? _04399_ : _04405_);
	assign _04407_ = _02778_ | _01407_;
	assign _04408_ = _04407_ | _01398_;
	assign _04409_ = _01410_ & ~_04408_;
	assign _04410_ = \mchip.design.owner.tokens [53] & ~_04372_;
	assign _04411_ = _04410_ | _04409_;
	assign _00060_ = (_05827_ ? _04406_ : _04411_);
	assign _04413_ = _02785_ | _01257_;
	assign _04414_ = _04413_ | _01261_;
	assign _04415_ = _01243_ & ~_04414_;
	assign _04416_ = _02789_ | _01257_;
	assign _04417_ = _04416_ | _01261_;
	assign _04418_ = _01243_ & ~_04417_;
	assign _04419_ = \mchip.design.owner.tokens [54] & ~_04418_;
	assign _04420_ = _04419_ | _04415_;
	assign _04421_ = _02796_ | _01284_;
	assign _04423_ = _04421_ | _01288_;
	assign _04424_ = _01274_ & ~_04423_;
	assign _04425_ = _02800_ | _01284_;
	assign _04426_ = _04425_ | _01288_;
	assign _04427_ = _01274_ & ~_04426_;
	assign _04428_ = \mchip.design.owner.tokens [54] & ~_04427_;
	assign _04429_ = _04428_ | _04424_;
	assign _04430_ = (_00199_ ? _04420_ : _04429_);
	assign _04431_ = _02808_ | _01314_;
	assign _04432_ = _04431_ | _01318_;
	assign _04434_ = _01303_ & ~_04432_;
	assign _04435_ = _02813_ | _01314_;
	assign _04436_ = _04435_ | _01318_;
	assign _04437_ = _01303_ & ~_04436_;
	assign _04438_ = \mchip.design.owner.tokens [54] & ~_04437_;
	assign _04439_ = _04438_ | _04434_;
	assign _04440_ = (_00131_ ? _04430_ : _04439_);
	assign _04441_ = _02820_ | _01343_;
	assign _04442_ = _04441_ | _01346_;
	assign _04443_ = _01349_ & ~_04442_;
	assign _04445_ = _02825_ | _01343_;
	assign _04446_ = _04445_ | _01346_;
	assign _04447_ = _01349_ & ~_04446_;
	assign _04448_ = \mchip.design.owner.tokens [54] & ~_04447_;
	assign _04449_ = _04448_ | _04443_;
	assign _04450_ = (_06005_ ? _04440_ : _04449_);
	assign _04451_ = _02832_ | _01377_;
	assign _04452_ = _04451_ | _01380_;
	assign _04453_ = _01382_ & ~_04452_;
	assign _04454_ = _02837_ | _01377_;
	assign _04456_ = _04454_ | _01380_;
	assign _04457_ = _01382_ & ~_04456_;
	assign _04458_ = \mchip.design.owner.tokens [54] & ~_04457_;
	assign _04459_ = _04458_ | _04453_;
	assign _04460_ = (_05934_ ? _04450_ : _04459_);
	assign _04461_ = _02844_ | _01407_;
	assign _04462_ = _04461_ | _01398_;
	assign _04463_ = _01410_ & ~_04462_;
	assign _04464_ = _02849_ | _01407_;
	assign _04465_ = _04464_ | _01398_;
	assign _04467_ = _01410_ & ~_04465_;
	assign _04468_ = \mchip.design.owner.tokens [54] & ~_04467_;
	assign _04469_ = _04468_ | _04463_;
	assign _00061_ = (_05827_ ? _04460_ : _04469_);
	assign _04470_ = _02856_ | _01257_;
	assign _04471_ = _04470_ | _01261_;
	assign _04472_ = _01243_ & ~_04471_;
	assign _04473_ = \mchip.design.owner.tokens [55] & ~_04418_;
	assign _04474_ = _04473_ | _04472_;
	assign _04475_ = _02862_ | _01284_;
	assign _04477_ = _04475_ | _01288_;
	assign _04478_ = _01274_ & ~_04477_;
	assign _04479_ = \mchip.design.owner.tokens [55] & ~_04427_;
	assign _04480_ = _04479_ | _04478_;
	assign _04481_ = (_00199_ ? _04474_ : _04480_);
	assign _04482_ = _02870_ | _01314_;
	assign _04483_ = _04482_ | _01318_;
	assign _04484_ = _01303_ & ~_04483_;
	assign _04485_ = \mchip.design.owner.tokens [55] & ~_04437_;
	assign _04486_ = _04485_ | _04484_;
	assign _04488_ = (_00131_ ? _04481_ : _04486_);
	assign _04489_ = _02878_ | _01343_;
	assign _04490_ = _04489_ | _01346_;
	assign _04491_ = _01349_ & ~_04490_;
	assign _04492_ = \mchip.design.owner.tokens [55] & ~_04447_;
	assign _04493_ = _04492_ | _04491_;
	assign _04494_ = (_06005_ ? _04488_ : _04493_);
	assign _04495_ = _02885_ | _01377_;
	assign _04496_ = _04495_ | _01380_;
	assign _04497_ = _01382_ & ~_04496_;
	assign _04499_ = \mchip.design.owner.tokens [55] & ~_04457_;
	assign _04500_ = _04499_ | _04497_;
	assign _04501_ = (_05934_ ? _04494_ : _04500_);
	assign _04502_ = _02893_ | _01407_;
	assign _04503_ = _04502_ | _01398_;
	assign _04504_ = _01410_ & ~_04503_;
	assign _04505_ = \mchip.design.owner.tokens [55] & ~_04467_;
	assign _04506_ = _04505_ | _04504_;
	assign _00062_ = (_05827_ ? _04501_ : _04506_);
	assign _04507_ = _02900_ | _01257_;
	assign _04509_ = _04507_ | _01261_;
	assign _04510_ = _01243_ & ~_04509_;
	assign _04511_ = _02904_ | _01257_;
	assign _04512_ = _04511_ | _01261_;
	assign _04513_ = _01243_ & ~_04512_;
	assign _04514_ = \mchip.design.owner.tokens [56] & ~_04513_;
	assign _04515_ = _04514_ | _04510_;
	assign _04516_ = _02911_ | _01284_;
	assign _04517_ = _04516_ | _01288_;
	assign _04518_ = _01274_ & ~_04517_;
	assign _04520_ = _02915_ | _01284_;
	assign _04521_ = _04520_ | _01288_;
	assign _04522_ = _01274_ & ~_04521_;
	assign _04523_ = \mchip.design.owner.tokens [56] & ~_04522_;
	assign _04524_ = _04523_ | _04518_;
	assign _04525_ = (_00199_ ? _04515_ : _04524_);
	assign _04526_ = _02923_ | _01314_;
	assign _04527_ = _04526_ | _01318_;
	assign _04528_ = _01303_ & ~_04527_;
	assign _04529_ = _02927_ | _01314_;
	assign _04531_ = _04529_ | _01318_;
	assign _04532_ = _01303_ & ~_04531_;
	assign _04533_ = \mchip.design.owner.tokens [56] & ~_04532_;
	assign _04534_ = _04533_ | _04528_;
	assign _04535_ = (_00131_ ? _04525_ : _04534_);
	assign _04536_ = _02935_ | _01343_;
	assign _04537_ = _04536_ | _01346_;
	assign _04538_ = _01349_ & ~_04537_;
	assign _04539_ = _02939_ | _01343_;
	assign _04540_ = _04539_ | _01346_;
	assign _04542_ = _01349_ & ~_04540_;
	assign _04543_ = \mchip.design.owner.tokens [56] & ~_04542_;
	assign _04544_ = _04543_ | _04538_;
	assign _04545_ = (_06005_ ? _04535_ : _04544_);
	assign _04546_ = _02947_ | _01377_;
	assign _04547_ = _04546_ | _01380_;
	assign _04548_ = _01382_ & ~_04547_;
	assign _04549_ = _02951_ | _01377_;
	assign _04550_ = _04549_ | _01380_;
	assign _04551_ = _01382_ & ~_04550_;
	assign _04553_ = \mchip.design.owner.tokens [56] & ~_04551_;
	assign _04554_ = _04553_ | _04548_;
	assign _04555_ = (_05934_ ? _04545_ : _04554_);
	assign _04556_ = _02959_ | _01407_;
	assign _04557_ = _04556_ | _01398_;
	assign _04558_ = _01410_ & ~_04557_;
	assign _04559_ = _02963_ | _01407_;
	assign _04560_ = _04559_ | _01398_;
	assign _04561_ = _01410_ & ~_04560_;
	assign _04562_ = \mchip.design.owner.tokens [56] & ~_04561_;
	assign _04564_ = _04562_ | _04558_;
	assign _00063_ = (_05827_ ? _04555_ : _04564_);
	assign _04565_ = _02970_ | _01257_;
	assign _04566_ = _04565_ | _01261_;
	assign _04567_ = _01243_ & ~_04566_;
	assign _04568_ = \mchip.design.owner.tokens [57] & ~_04513_;
	assign _04569_ = _04568_ | _04567_;
	assign _04570_ = _02977_ | _01284_;
	assign _04571_ = _04570_ | _01288_;
	assign _04572_ = _01274_ & ~_04571_;
	assign _04574_ = \mchip.design.owner.tokens [57] & ~_04522_;
	assign _04575_ = _04574_ | _04572_;
	assign _04576_ = (_00199_ ? _04569_ : _04575_);
	assign _04577_ = _02984_ | _01314_;
	assign _04578_ = _04577_ | _01318_;
	assign _04579_ = _01303_ & ~_04578_;
	assign _04580_ = \mchip.design.owner.tokens [57] & ~_04532_;
	assign _04581_ = _04580_ | _04579_;
	assign _04582_ = (_00131_ ? _04576_ : _04581_);
	assign _04583_ = _02992_ | _01343_;
	assign _04585_ = _04583_ | _01346_;
	assign _04586_ = _01349_ & ~_04585_;
	assign _04587_ = \mchip.design.owner.tokens [57] & ~_04542_;
	assign _04588_ = _04587_ | _04586_;
	assign _04589_ = (_06005_ ? _04582_ : _04588_);
	assign _04590_ = _03000_ | _01377_;
	assign _04591_ = _04590_ | _01380_;
	assign _04592_ = _01382_ & ~_04591_;
	assign _04593_ = \mchip.design.owner.tokens [57] & ~_04551_;
	assign _04594_ = _04593_ | _04592_;
	assign _04596_ = (_05934_ ? _04589_ : _04594_);
	assign _04597_ = _03008_ | _01407_;
	assign _04598_ = _04597_ | _01398_;
	assign _04599_ = _01410_ & ~_04598_;
	assign _04600_ = \mchip.design.owner.tokens [57] & ~_04561_;
	assign _04601_ = _04600_ | _04599_;
	assign _00064_ = (_05827_ ? _04596_ : _04601_);
	assign _04602_ = _03014_ | _01257_;
	assign _04603_ = _04602_ | _01261_;
	assign _04604_ = _01243_ & ~_04603_;
	assign _04606_ = _03019_ | _01257_;
	assign _04607_ = _04606_ | _01261_;
	assign _04608_ = _01243_ & ~_04607_;
	assign _04609_ = \mchip.design.owner.tokens [58] & ~_04608_;
	assign _04610_ = _04609_ | _04604_;
	assign _04611_ = _03025_ | _01284_;
	assign _04612_ = _04611_ | _01288_;
	assign _04613_ = _01274_ & ~_04612_;
	assign _04614_ = _03030_ | _01284_;
	assign _04615_ = _04614_ | _01288_;
	assign _04617_ = _01274_ & ~_04615_;
	assign _04618_ = \mchip.design.owner.tokens [58] & ~_04617_;
	assign _04619_ = _04618_ | _04613_;
	assign _04620_ = (_00199_ ? _04610_ : _04619_);
	assign _04621_ = _03037_ | _01314_;
	assign _04622_ = _04621_ | _01318_;
	assign _04623_ = _01303_ & ~_04622_;
	assign _04624_ = _03042_ | _01314_;
	assign _04625_ = _04624_ | _01318_;
	assign _04626_ = _01303_ & ~_04625_;
	assign _04628_ = \mchip.design.owner.tokens [58] & ~_04626_;
	assign _04629_ = _04628_ | _04623_;
	assign _04630_ = (_00131_ ? _04620_ : _04629_);
	assign _04631_ = _03049_ | _01343_;
	assign _04632_ = _04631_ | _01346_;
	assign _04633_ = _01349_ & ~_04632_;
	assign _04634_ = _03054_ | _01343_;
	assign _04635_ = _04634_ | _01346_;
	assign _04636_ = _01349_ & ~_04635_;
	assign _04637_ = \mchip.design.owner.tokens [58] & ~_04636_;
	assign _04639_ = _04637_ | _04633_;
	assign _04640_ = (_06005_ ? _04630_ : _04639_);
	assign _04641_ = _03062_ | _01377_;
	assign _04642_ = _04641_ | _01380_;
	assign _04643_ = _01382_ & ~_04642_;
	assign _04644_ = _03066_ | _01377_;
	assign _04645_ = _04644_ | _01380_;
	assign _04646_ = _01382_ & ~_04645_;
	assign _04647_ = \mchip.design.owner.tokens [58] & ~_04646_;
	assign _04648_ = _04647_ | _04643_;
	assign _04650_ = (_05934_ ? _04640_ : _04648_);
	assign _04651_ = _03074_ | _01407_;
	assign _04652_ = _04651_ | _01398_;
	assign _04653_ = _01410_ & ~_04652_;
	assign _04654_ = _03078_ | _01407_;
	assign _04655_ = _04654_ | _01398_;
	assign _04656_ = _01410_ & ~_04655_;
	assign _04657_ = \mchip.design.owner.tokens [58] & ~_04656_;
	assign _04658_ = _04657_ | _04653_;
	assign _00065_ = (_05827_ ? _04650_ : _04658_);
	assign _04660_ = _03085_ | _01257_;
	assign _04661_ = _04660_ | _01261_;
	assign _04662_ = _01243_ & ~_04661_;
	assign _04663_ = \mchip.design.owner.tokens [59] & ~_04608_;
	assign _04664_ = _04663_ | _04662_;
	assign _04665_ = _03091_ | _01284_;
	assign _04666_ = _04665_ | _01288_;
	assign _04667_ = _01274_ & ~_04666_;
	assign _04668_ = \mchip.design.owner.tokens [59] & ~_04617_;
	assign _04669_ = _04668_ | _04667_;
	assign _04671_ = (_00199_ ? _04664_ : _04669_);
	assign _04672_ = _03099_ | _01314_;
	assign _04673_ = _04672_ | _01318_;
	assign _04674_ = _01303_ & ~_04673_;
	assign _04675_ = \mchip.design.owner.tokens [59] & ~_04626_;
	assign _04676_ = _04675_ | _04674_;
	assign _04677_ = (_00131_ ? _04671_ : _04676_);
	assign _04678_ = _03107_ | _01343_;
	assign _04679_ = _04678_ | _01346_;
	assign _04680_ = _01349_ & ~_04679_;
	assign _04682_ = \mchip.design.owner.tokens [59] & ~_04636_;
	assign _04683_ = _04682_ | _04680_;
	assign _04684_ = (_06005_ ? _04677_ : _04683_);
	assign _04685_ = _03114_ | _01377_;
	assign _04686_ = _04685_ | _01380_;
	assign _04687_ = _01382_ & ~_04686_;
	assign _04688_ = \mchip.design.owner.tokens [59] & ~_04646_;
	assign _04689_ = _04688_ | _04687_;
	assign _04690_ = (_05934_ ? _04684_ : _04689_);
	assign _04691_ = _03122_ | _01407_;
	assign _04693_ = _04691_ | _01398_;
	assign _04694_ = _01410_ & ~_04693_;
	assign _04695_ = \mchip.design.owner.tokens [59] & ~_04656_;
	assign _04696_ = _04695_ | _04694_;
	assign _00066_ = (_05827_ ? _04690_ : _04696_);
	assign _04697_ = _03128_ | _01257_;
	assign _04698_ = _04697_ | _01261_;
	assign _04699_ = _01243_ & ~_04698_;
	assign _04700_ = _03132_ | _01257_;
	assign _04701_ = _04700_ | _01261_;
	assign _04703_ = _01243_ & ~_04701_;
	assign _04704_ = \mchip.design.owner.tokens [60] & ~_04703_;
	assign _04705_ = _04704_ | _04699_;
	assign _04706_ = _03139_ | _01284_;
	assign _04707_ = _04706_ | _01288_;
	assign _04708_ = _01274_ & ~_04707_;
	assign _04709_ = _03143_ | _01284_;
	assign _04710_ = _04709_ | _01288_;
	assign _04711_ = _01274_ & ~_04710_;
	assign _04712_ = \mchip.design.owner.tokens [60] & ~_04711_;
	assign _04714_ = _04712_ | _04708_;
	assign _04715_ = (_00199_ ? _04705_ : _04714_);
	assign _04716_ = _03151_ | _01314_;
	assign _04717_ = _04716_ | _01318_;
	assign _04718_ = _01303_ & ~_04717_;
	assign _04719_ = _03155_ | _01314_;
	assign _04720_ = _04719_ | _01318_;
	assign _04721_ = _01303_ & ~_04720_;
	assign _04722_ = \mchip.design.owner.tokens [60] & ~_04721_;
	assign _04723_ = _04722_ | _04718_;
	assign _04725_ = (_00131_ ? _04715_ : _04723_);
	assign _04726_ = _03163_ | _01343_;
	assign _04727_ = _04726_ | _01346_;
	assign _04728_ = _01349_ & ~_04727_;
	assign _04729_ = _03167_ | _01343_;
	assign _04730_ = _04729_ | _01346_;
	assign _04731_ = _01349_ & ~_04730_;
	assign _04732_ = \mchip.design.owner.tokens [60] & ~_04731_;
	assign _04733_ = _04732_ | _04728_;
	assign _04734_ = (_06005_ ? _04725_ : _04733_);
	assign _04736_ = _03175_ | _01377_;
	assign _04737_ = _04736_ | _01380_;
	assign _04738_ = _01382_ & ~_04737_;
	assign _04739_ = _03180_ | _01377_;
	assign _04740_ = _04739_ | _01380_;
	assign _04741_ = _01382_ & ~_04740_;
	assign _04742_ = \mchip.design.owner.tokens [60] & ~_04741_;
	assign _04743_ = _04742_ | _04738_;
	assign _04744_ = (_05934_ ? _04734_ : _04743_);
	assign _04745_ = _03187_ | _01407_;
	assign _04747_ = _04745_ | _01398_;
	assign _04748_ = _01410_ & ~_04747_;
	assign _04749_ = _03192_ | _01407_;
	assign _04750_ = _04749_ | _01398_;
	assign _04751_ = _01410_ & ~_04750_;
	assign _04752_ = \mchip.design.owner.tokens [60] & ~_04751_;
	assign _04753_ = _04752_ | _04748_;
	assign _00068_ = (_05827_ ? _04744_ : _04753_);
	assign _04754_ = _03198_ | _01257_;
	assign _04755_ = _04754_ | _01261_;
	assign _04757_ = _01243_ & ~_04755_;
	assign _04758_ = \mchip.design.owner.tokens [61] & ~_04703_;
	assign _04759_ = _04758_ | _04757_;
	assign _04760_ = _03205_ | _01284_;
	assign _04761_ = _04760_ | _01288_;
	assign _04762_ = _01274_ & ~_04761_;
	assign _04763_ = \mchip.design.owner.tokens [61] & ~_04711_;
	assign _04764_ = _04763_ | _04762_;
	assign _04765_ = (_00199_ ? _04759_ : _04764_);
	assign _04766_ = _03213_ | _01314_;
	assign _04768_ = _04766_ | _01318_;
	assign _04769_ = _01303_ & ~_04768_;
	assign _04770_ = \mchip.design.owner.tokens [61] & ~_04721_;
	assign _04771_ = _04770_ | _04769_;
	assign _04772_ = (_00131_ ? _04765_ : _04771_);
	assign _04773_ = _03220_ | _01343_;
	assign _04774_ = _04773_ | _01346_;
	assign _04775_ = _01349_ & ~_04774_;
	assign _04776_ = \mchip.design.owner.tokens [61] & ~_04731_;
	assign _04777_ = _04776_ | _04775_;
	assign _04779_ = (_06005_ ? _04772_ : _04777_);
	assign _04780_ = _03228_ | _01377_;
	assign _04781_ = _04780_ | _01380_;
	assign _04782_ = _01382_ & ~_04781_;
	assign _04783_ = \mchip.design.owner.tokens [61] & ~_04741_;
	assign _04784_ = _04783_ | _04782_;
	assign _04785_ = (_05934_ ? _04779_ : _04784_);
	assign _04786_ = _03236_ | _01407_;
	assign _04787_ = _04786_ | _01398_;
	assign _04788_ = _01410_ & ~_04787_;
	assign _04790_ = \mchip.design.owner.tokens [61] & ~_04751_;
	assign _04791_ = _04790_ | _04788_;
	assign _00069_ = (_05827_ ? _04785_ : _04791_);
	assign _04792_ = _03242_ | _01257_;
	assign _04793_ = _04792_ | _01261_;
	assign _04794_ = _01243_ & ~_04793_;
	assign _04795_ = _03247_ | _01257_;
	assign _04796_ = _04795_ | _01261_;
	assign _04797_ = _01243_ & ~_04796_;
	assign _04798_ = \mchip.design.owner.tokens [62] & ~_04797_;
	assign _04800_ = _04798_ | _04794_;
	assign _04801_ = _03253_ | _01284_;
	assign _04802_ = _04801_ | _01288_;
	assign _04803_ = _01274_ & ~_04802_;
	assign _04804_ = _03258_ | _01284_;
	assign _04805_ = _04804_ | _01288_;
	assign _04806_ = _01274_ & ~_04805_;
	assign _04807_ = \mchip.design.owner.tokens [62] & ~_04806_;
	assign _04808_ = _04807_ | _04803_;
	assign _04809_ = (_00199_ ? _04800_ : _04808_);
	assign _04811_ = _03266_ | _01314_;
	assign _04812_ = _04811_ | _01318_;
	assign _04813_ = _01303_ & ~_04812_;
	assign _04814_ = _03270_ | _01314_;
	assign _04815_ = _04814_ | _01318_;
	assign _04816_ = _01303_ & ~_04815_;
	assign _04817_ = \mchip.design.owner.tokens [62] & ~_04816_;
	assign _04818_ = _04817_ | _04813_;
	assign _04819_ = (_00131_ ? _04809_ : _04818_);
	assign _04820_ = _03278_ | _01343_;
	assign _04822_ = _04820_ | _01346_;
	assign _04823_ = _01349_ & ~_04822_;
	assign _04824_ = _03282_ | _01343_;
	assign _04825_ = _04824_ | _01346_;
	assign _04826_ = _01349_ & ~_04825_;
	assign _04827_ = \mchip.design.owner.tokens [62] & ~_04826_;
	assign _04828_ = _04827_ | _04823_;
	assign _04829_ = (_06005_ ? _04819_ : _04828_);
	assign _04830_ = _03290_ | _01377_;
	assign _04831_ = _04830_ | _01380_;
	assign _04833_ = _01382_ & ~_04831_;
	assign _04834_ = _03294_ | _01377_;
	assign _04835_ = _04834_ | _01380_;
	assign _04836_ = _01382_ & ~_04835_;
	assign _04837_ = \mchip.design.owner.tokens [62] & ~_04836_;
	assign _04838_ = _04837_ | _04833_;
	assign _04839_ = (_05934_ ? _04829_ : _04838_);
	assign _04840_ = _03302_ | _01407_;
	assign _04841_ = _04840_ | _01398_;
	assign _04842_ = _01410_ & ~_04841_;
	assign _04844_ = _03306_ | _01407_;
	assign _04845_ = _04844_ | _01398_;
	assign _04846_ = _01410_ & ~_04845_;
	assign _04847_ = \mchip.design.owner.tokens [62] & ~_04846_;
	assign _04848_ = _04847_ | _04842_;
	assign _00070_ = (_05827_ ? _04839_ : _04848_);
	assign _04849_ = _03313_ | _01257_;
	assign _04850_ = _04849_ | _01261_;
	assign _04851_ = _01243_ & ~_04850_;
	assign _04852_ = \mchip.design.owner.tokens [63] & ~_04797_;
	assign _04854_ = _04852_ | _04851_;
	assign _04855_ = _03320_ | _01284_;
	assign _04856_ = _04855_ | _01288_;
	assign _04857_ = _01274_ & ~_04856_;
	assign _04858_ = \mchip.design.owner.tokens [63] & ~_04806_;
	assign _04859_ = _04858_ | _04857_;
	assign _04860_ = (_00199_ ? _04854_ : _04859_);
	assign _04861_ = _03327_ | _01314_;
	assign _04862_ = _04861_ | _01318_;
	assign _04863_ = _01303_ & ~_04862_;
	assign _04865_ = \mchip.design.owner.tokens [63] & ~_04816_;
	assign _04866_ = _04865_ | _04863_;
	assign _04867_ = (_00131_ ? _04860_ : _04866_);
	assign _04868_ = _03335_ | _01343_;
	assign _04869_ = _04868_ | _01346_;
	assign _04870_ = _01349_ & ~_04869_;
	assign _04871_ = \mchip.design.owner.tokens [63] & ~_04826_;
	assign _04872_ = _04871_ | _04870_;
	assign _04873_ = (_06005_ ? _04867_ : _04872_);
	assign _04874_ = _03343_ | _01377_;
	assign _04876_ = _04874_ | _01380_;
	assign _04877_ = _01382_ & ~_04876_;
	assign _04878_ = \mchip.design.owner.tokens [63] & ~_04836_;
	assign _04879_ = _04878_ | _04877_;
	assign _04880_ = (_05934_ ? _04873_ : _04879_);
	assign _04881_ = _03350_ | _01407_;
	assign _04882_ = _04881_ | _01398_;
	assign _04883_ = _01410_ & ~_04882_;
	assign _04884_ = \mchip.design.owner.tokens [63] & ~_04846_;
	assign _04885_ = _04884_ | _04883_;
	assign _00071_ = (_05827_ ? _04880_ : _04885_);
	assign _04887_ = _03357_ | _01257_;
	assign _04888_ = _04887_ | _01261_;
	assign _04889_ = _01243_ & ~_04888_;
	assign _04890_ = _03361_ | _01257_;
	assign _04891_ = _04890_ | _01261_;
	assign _04892_ = _01243_ & ~_04891_;
	assign _04893_ = \mchip.design.owner.tokens [64] & ~_04892_;
	assign _04894_ = _04893_ | _04889_;
	assign _04895_ = _03368_ | _01284_;
	assign _04897_ = _04895_ | _01288_;
	assign _04898_ = _01274_ & ~_04897_;
	assign _04899_ = _03372_ | _01284_;
	assign _04900_ = _04899_ | _01288_;
	assign _04901_ = _01274_ & ~_04900_;
	assign _04902_ = \mchip.design.owner.tokens [64] & ~_04901_;
	assign _04903_ = _04902_ | _04898_;
	assign _04904_ = (_00199_ ? _04894_ : _04903_);
	assign _04905_ = _03380_ | _01314_;
	assign _04906_ = _04905_ | _01318_;
	assign _04908_ = _01303_ & ~_04906_;
	assign _04909_ = _03385_ | _01314_;
	assign _04910_ = _04909_ | _01318_;
	assign _04911_ = _01303_ & ~_04910_;
	assign _04912_ = \mchip.design.owner.tokens [64] & ~_04911_;
	assign _04913_ = _04912_ | _04908_;
	assign _04914_ = (_00131_ ? _04904_ : _04913_);
	assign _04915_ = _03392_ | _01343_;
	assign _04916_ = _04915_ | _01346_;
	assign _04917_ = _01349_ & ~_04916_;
	assign _04919_ = _03397_ | _01343_;
	assign _04920_ = _04919_ | _01346_;
	assign _04921_ = _01349_ & ~_04920_;
	assign _04922_ = \mchip.design.owner.tokens [64] & ~_04921_;
	assign _04923_ = _04922_ | _04917_;
	assign _04924_ = (_06005_ ? _04914_ : _04923_);
	assign _04925_ = _03404_ | _01377_;
	assign _04926_ = _04925_ | _01380_;
	assign _04927_ = _01382_ & ~_04926_;
	assign _04928_ = _03409_ | _01377_;
	assign _04930_ = _04928_ | _01380_;
	assign _04931_ = _01382_ & ~_04930_;
	assign _04932_ = \mchip.design.owner.tokens [64] & ~_04931_;
	assign _04933_ = _04932_ | _04927_;
	assign _04934_ = (_05934_ ? _04924_ : _04933_);
	assign _04935_ = _03416_ | _01407_;
	assign _04936_ = _04935_ | _01398_;
	assign _04937_ = _01410_ & ~_04936_;
	assign _04938_ = _03421_ | _01407_;
	assign _04939_ = _04938_ | _01398_;
	assign _04941_ = _01410_ & ~_04939_;
	assign _04942_ = \mchip.design.owner.tokens [64] & ~_04941_;
	assign _04943_ = _04942_ | _04937_;
	assign _00072_ = (_05827_ ? _04934_ : _04943_);
	assign _04944_ = _03428_ | _01257_;
	assign _04945_ = _04944_ | _01261_;
	assign _04946_ = _01243_ & ~_04945_;
	assign _04947_ = \mchip.design.owner.tokens [65] & ~_04892_;
	assign _04948_ = _04947_ | _04946_;
	assign _04949_ = _03434_ | _01284_;
	assign _04951_ = _04949_ | _01288_;
	assign _04952_ = _01274_ & ~_04951_;
	assign _04953_ = \mchip.design.owner.tokens [65] & ~_04901_;
	assign _04954_ = _04953_ | _04952_;
	assign _04955_ = (_00199_ ? _04948_ : _04954_);
	assign _04956_ = _03442_ | _01314_;
	assign _04957_ = _04956_ | _01318_;
	assign _04958_ = _01303_ & ~_04957_;
	assign _04959_ = \mchip.design.owner.tokens [65] & ~_04911_;
	assign _04960_ = _04959_ | _04958_;
	assign _04962_ = (_00131_ ? _04955_ : _04960_);
	assign _04963_ = _03450_ | _01343_;
	assign _04964_ = _04963_ | _01346_;
	assign _04965_ = _01349_ & ~_04964_;
	assign _04966_ = \mchip.design.owner.tokens [65] & ~_04921_;
	assign _04967_ = _04966_ | _04965_;
	assign _04968_ = (_06005_ ? _04962_ : _04967_);
	assign _04969_ = _03457_ | _01377_;
	assign _04970_ = _04969_ | _01380_;
	assign _04971_ = _01382_ & ~_04970_;
	assign _04973_ = \mchip.design.owner.tokens [65] & ~_04931_;
	assign _04974_ = _04973_ | _04971_;
	assign _04975_ = (_05934_ ? _04968_ : _04974_);
	assign _04976_ = _03465_ | _01407_;
	assign _04977_ = _04976_ | _01398_;
	assign _04978_ = _01410_ & ~_04977_;
	assign _04979_ = \mchip.design.owner.tokens [65] & ~_04941_;
	assign _04980_ = _04979_ | _04978_;
	assign _00073_ = (_05827_ ? _04975_ : _04980_);
	assign _04981_ = _01496_ | ~_01261_;
	assign _04983_ = _01243_ & ~_04981_;
	assign _04984_ = _01501_ | ~_01261_;
	assign _04985_ = _01243_ & ~_04984_;
	assign _04986_ = \mchip.design.owner.tokens [66] & ~_04985_;
	assign _04987_ = _04986_ | _04983_;
	assign _04988_ = _01512_ | ~_01288_;
	assign _04989_ = _01274_ & ~_04988_;
	assign _04990_ = _01517_ | ~_01288_;
	assign _04991_ = _01274_ & ~_04990_;
	assign _04992_ = \mchip.design.owner.tokens [66] & ~_04991_;
	assign _04994_ = _04992_ | _04989_;
	assign _04995_ = (_00199_ ? _04987_ : _04994_);
	assign _04996_ = _01529_ | ~_01318_;
	assign _04997_ = _01303_ & ~_04996_;
	assign _04998_ = _01534_ | ~_01318_;
	assign _04999_ = _01303_ & ~_04998_;
	assign _05000_ = \mchip.design.owner.tokens [66] & ~_04999_;
	assign _05001_ = _05000_ | _04997_;
	assign _05002_ = (_00131_ ? _04995_ : _05001_);
	assign _05003_ = _01547_ | ~_01346_;
	assign _05005_ = _01349_ & ~_05003_;
	assign _05006_ = _01552_ | ~_01346_;
	assign _05007_ = _01349_ & ~_05006_;
	assign _05008_ = \mchip.design.owner.tokens [66] & ~_05007_;
	assign _05009_ = _05008_ | _05005_;
	assign _05010_ = (_06005_ ? _05002_ : _05009_);
	assign _05011_ = _01564_ | ~_01380_;
	assign _05012_ = _01382_ & ~_05011_;
	assign _05013_ = _01569_ | ~_01380_;
	assign _05014_ = _01382_ & ~_05013_;
	assign _05016_ = \mchip.design.owner.tokens [66] & ~_05014_;
	assign _05017_ = _05016_ | _05012_;
	assign _05018_ = (_05934_ ? _05010_ : _05017_);
	assign _05019_ = _01581_ | ~_01398_;
	assign _05020_ = _01410_ & ~_05019_;
	assign _05021_ = _01588_ | ~_01398_;
	assign _05022_ = _01410_ & ~_05021_;
	assign _05023_ = \mchip.design.owner.tokens [66] & ~_05022_;
	assign _05024_ = _05023_ | _05020_;
	assign _00074_ = (_05827_ ? _05018_ : _05024_);
	assign _05026_ = _01598_ | ~_01261_;
	assign _05027_ = _01243_ & ~_05026_;
	assign _05028_ = \mchip.design.owner.tokens [67] & ~_04985_;
	assign _05029_ = _05028_ | _05027_;
	assign _05030_ = _01608_ | ~_01288_;
	assign _05031_ = _01274_ & ~_05030_;
	assign _05032_ = \mchip.design.owner.tokens [67] & ~_04991_;
	assign _05033_ = _05032_ | _05031_;
	assign _05034_ = (_00199_ ? _05029_ : _05033_);
	assign _05035_ = _01619_ | ~_01318_;
	assign _05037_ = _01303_ & ~_05035_;
	assign _05038_ = \mchip.design.owner.tokens [67] & ~_04999_;
	assign _05039_ = _05038_ | _05037_;
	assign _05040_ = (_00131_ ? _05034_ : _05039_);
	assign _05041_ = _01630_ | ~_01346_;
	assign _05042_ = _01349_ & ~_05041_;
	assign _05043_ = \mchip.design.owner.tokens [67] & ~_05007_;
	assign _05044_ = _05043_ | _05042_;
	assign _05045_ = (_06005_ ? _05040_ : _05044_);
	assign _05046_ = _01641_ | ~_01380_;
	assign _05048_ = _01382_ & ~_05046_;
	assign _05049_ = \mchip.design.owner.tokens [67] & ~_05014_;
	assign _05050_ = _05049_ | _05048_;
	assign _05051_ = (_05934_ ? _05045_ : _05050_);
	assign _05052_ = _01652_ | ~_01398_;
	assign _05053_ = _01410_ & ~_05052_;
	assign _05054_ = \mchip.design.owner.tokens [67] & ~_05022_;
	assign _05055_ = _05054_ | _05053_;
	assign _00075_ = (_05827_ ? _05051_ : _05055_);
	assign _05056_ = _01661_ | ~_01261_;
	assign _05058_ = _01243_ & ~_05056_;
	assign _05059_ = _01666_ | ~_01261_;
	assign _05060_ = _01243_ & ~_05059_;
	assign _05061_ = \mchip.design.owner.tokens [68] & ~_05060_;
	assign _05062_ = _05061_ | _05058_;
	assign _05063_ = _01675_ | ~_01288_;
	assign _05064_ = _01274_ & ~_05063_;
	assign _05065_ = _01680_ | ~_01288_;
	assign _05066_ = _01274_ & ~_05065_;
	assign _05067_ = \mchip.design.owner.tokens [68] & ~_05066_;
	assign _05069_ = _05067_ | _05064_;
	assign _05070_ = (_00199_ ? _05062_ : _05069_);
	assign _05071_ = _01690_ | ~_01318_;
	assign _05072_ = _01303_ & ~_05071_;
	assign _05073_ = _01695_ | ~_01318_;
	assign _05074_ = _01303_ & ~_05073_;
	assign _05075_ = \mchip.design.owner.tokens [68] & ~_05074_;
	assign _05076_ = _05075_ | _05072_;
	assign _05077_ = (_00131_ ? _05070_ : _05076_);
	assign _05078_ = _01705_ | ~_01346_;
	assign _05080_ = _01349_ & ~_05078_;
	assign _05081_ = _01710_ | ~_01346_;
	assign _05082_ = _01349_ & ~_05081_;
	assign _05083_ = \mchip.design.owner.tokens [68] & ~_05082_;
	assign _05084_ = _05083_ | _05080_;
	assign _05085_ = (_06005_ ? _05077_ : _05084_);
	assign _05086_ = _01720_ | ~_01380_;
	assign _05087_ = _01382_ & ~_05086_;
	assign _05088_ = _01728_ | ~_01380_;
	assign _05089_ = _01382_ & ~_05088_;
	assign _05091_ = \mchip.design.owner.tokens [68] & ~_05089_;
	assign _05092_ = _05091_ | _05087_;
	assign _05093_ = (_05934_ ? _05085_ : _05092_);
	assign _05094_ = _01738_ | ~_01398_;
	assign _05095_ = _01410_ & ~_05094_;
	assign _05096_ = _01745_ | ~_01398_;
	assign _05097_ = _01410_ & ~_05096_;
	assign _05098_ = \mchip.design.owner.tokens [68] & ~_05097_;
	assign _05099_ = _05098_ | _05095_;
	assign _00076_ = (_05827_ ? _05093_ : _05099_);
	assign _05101_ = _01754_ | ~_01261_;
	assign _05102_ = _01243_ & ~_05101_;
	assign _05103_ = \mchip.design.owner.tokens [69] & ~_05060_;
	assign _05104_ = _05103_ | _05102_;
	assign _05105_ = _01763_ | ~_01288_;
	assign _05106_ = _01274_ & ~_05105_;
	assign _05107_ = \mchip.design.owner.tokens [69] & ~_05066_;
	assign _05108_ = _05107_ | _05106_;
	assign _05109_ = (_00199_ ? _05104_ : _05108_);
	assign _05110_ = _01773_ | ~_01318_;
	assign _05112_ = _01303_ & ~_05110_;
	assign _05113_ = \mchip.design.owner.tokens [69] & ~_05074_;
	assign _05114_ = _05113_ | _05112_;
	assign _05115_ = (_00131_ ? _05109_ : _05114_);
	assign _05116_ = _01783_ | ~_01346_;
	assign _05117_ = _01349_ & ~_05116_;
	assign _05118_ = \mchip.design.owner.tokens [69] & ~_05082_;
	assign _05119_ = _05118_ | _05117_;
	assign _05120_ = (_06005_ ? _05115_ : _05119_);
	assign _05121_ = _01793_ | ~_01380_;
	assign _05123_ = _01382_ & ~_05121_;
	assign _05124_ = \mchip.design.owner.tokens [69] & ~_05089_;
	assign _05125_ = _05124_ | _05123_;
	assign _05126_ = (_05934_ ? _05120_ : _05125_);
	assign _05127_ = _01803_ | ~_01398_;
	assign _05128_ = _01410_ & ~_05127_;
	assign _05129_ = \mchip.design.owner.tokens [69] & ~_05097_;
	assign _05130_ = _05129_ | _05128_;
	assign _00077_ = (_05827_ ? _05126_ : _05130_);
	assign _05131_ = _01811_ | ~_01261_;
	assign _05133_ = _01243_ & ~_05131_;
	assign _05134_ = _01816_ | ~_01261_;
	assign _05135_ = _01243_ & ~_05134_;
	assign _05136_ = \mchip.design.owner.tokens [70] & ~_05135_;
	assign _05137_ = _05136_ | _05133_;
	assign _05138_ = _01824_ | ~_01288_;
	assign _05139_ = _01274_ & ~_05138_;
	assign _05140_ = _01829_ | ~_01288_;
	assign _05141_ = _01274_ & ~_05140_;
	assign _05142_ = \mchip.design.owner.tokens [70] & ~_05141_;
	assign _05144_ = _05142_ | _05139_;
	assign _05145_ = (_00199_ ? _05137_ : _05144_);
	assign _05146_ = _01838_ | ~_01318_;
	assign _05147_ = _01303_ & ~_05146_;
	assign _05148_ = _01843_ | ~_01318_;
	assign _05149_ = _01303_ & ~_05148_;
	assign _05150_ = \mchip.design.owner.tokens [70] & ~_05149_;
	assign _05151_ = _05150_ | _05147_;
	assign _05152_ = (_00131_ ? _05145_ : _05151_);
	assign _05153_ = _01852_ | ~_01346_;
	assign _05155_ = _01349_ & ~_05153_;
	assign _05156_ = _01857_ | ~_01346_;
	assign _05157_ = _01349_ & ~_05156_;
	assign _05158_ = \mchip.design.owner.tokens [70] & ~_05157_;
	assign _05159_ = _05158_ | _05155_;
	assign _05160_ = (_06005_ ? _05152_ : _05159_);
	assign _05161_ = _01866_ | ~_01380_;
	assign _05162_ = _01382_ & ~_05161_;
	assign _05163_ = _01873_ | ~_01380_;
	assign _05164_ = _01382_ & ~_05163_;
	assign _05166_ = \mchip.design.owner.tokens [70] & ~_05164_;
	assign _05167_ = _05166_ | _05162_;
	assign _05168_ = (_05934_ ? _05160_ : _05167_);
	assign _05169_ = _01882_ | ~_01398_;
	assign _05170_ = _01410_ & ~_05169_;
	assign _05171_ = _01888_ | ~_01398_;
	assign _05172_ = _01410_ & ~_05171_;
	assign _05173_ = \mchip.design.owner.tokens [70] & ~_05172_;
	assign _05174_ = _05173_ | _05170_;
	assign _00079_ = (_05827_ ? _05168_ : _05174_);
	assign _05175_ = _01896_ | ~_01261_;
	assign _05176_ = _01243_ & ~_05175_;
	assign _05177_ = \mchip.design.owner.tokens [71] & ~_05135_;
	assign _05178_ = _05177_ | _05176_;
	assign _05179_ = _01904_ | ~_01288_;
	assign _05180_ = _01274_ & ~_05179_;
	assign _05181_ = \mchip.design.owner.tokens [71] & ~_05141_;
	assign _05182_ = _05181_ | _05180_;
	assign _05183_ = (_00199_ ? _05178_ : _05182_);
	assign _05184_ = _01913_ | ~_01318_;
	assign _05186_ = _01303_ & ~_05184_;
	assign _05187_ = \mchip.design.owner.tokens [71] & ~_05149_;
	assign _05188_ = _05187_ | _05186_;
	assign _05189_ = (_00131_ ? _05183_ : _05188_);
	assign _05190_ = _01922_ | ~_01346_;
	assign _05191_ = _01349_ & ~_05190_;
	assign _05192_ = \mchip.design.owner.tokens [71] & ~_05157_;
	assign _05193_ = _05192_ | _05191_;
	assign _05194_ = (_06005_ ? _05189_ : _05193_);
	assign _05195_ = _01931_ | ~_01380_;
	assign _05197_ = _01382_ & ~_05195_;
	assign _05198_ = \mchip.design.owner.tokens [71] & ~_05164_;
	assign _05199_ = _05198_ | _05197_;
	assign _05200_ = (_05934_ ? _05194_ : _05199_);
	assign _05201_ = _01940_ | ~_01398_;
	assign _05202_ = _01410_ & ~_05201_;
	assign _05203_ = \mchip.design.owner.tokens [71] & ~_05172_;
	assign _05204_ = _05203_ | _05202_;
	assign _00080_ = (_05827_ ? _05200_ : _05204_);
	assign _05205_ = _01948_ | ~_01261_;
	assign _05207_ = _01243_ & ~_05205_;
	assign _05208_ = _01953_ | ~_01261_;
	assign _05209_ = _01243_ & ~_05208_;
	assign _05210_ = \mchip.design.owner.tokens [72] & ~_05209_;
	assign _05211_ = _05210_ | _05207_;
	assign _05212_ = _01961_ | ~_01288_;
	assign _05213_ = _01274_ & ~_05212_;
	assign _05214_ = _01966_ | ~_01288_;
	assign _05215_ = _01274_ & ~_05214_;
	assign _05216_ = \mchip.design.owner.tokens [72] & ~_05215_;
	assign _05218_ = _05216_ | _05213_;
	assign _05219_ = (_00199_ ? _05211_ : _05218_);
	assign _05220_ = _01975_ | ~_01318_;
	assign _05221_ = _01303_ & ~_05220_;
	assign _05222_ = _01980_ | ~_01318_;
	assign _05223_ = _01303_ & ~_05222_;
	assign _05224_ = \mchip.design.owner.tokens [72] & ~_05223_;
	assign _05225_ = _05224_ | _05221_;
	assign _05226_ = (_00131_ ? _05219_ : _05225_);
	assign _05227_ = _01989_ | ~_01346_;
	assign _05229_ = _01349_ & ~_05227_;
	assign _05230_ = _01994_ | ~_01346_;
	assign _05231_ = _01349_ & ~_05230_;
	assign _05232_ = \mchip.design.owner.tokens [72] & ~_05231_;
	assign _05233_ = _05232_ | _05229_;
	assign _05234_ = (_06005_ ? _05226_ : _05233_);
	assign _05235_ = _02003_ | ~_01380_;
	assign _05236_ = _01382_ & ~_05235_;
	assign _05237_ = _02009_ | ~_01380_;
	assign _05238_ = _01382_ & ~_05237_;
	assign _05240_ = \mchip.design.owner.tokens [72] & ~_05238_;
	assign _05241_ = _05240_ | _05236_;
	assign _05242_ = (_05934_ ? _05234_ : _05241_);
	assign _05243_ = _02018_ | ~_01398_;
	assign _05244_ = _01410_ & ~_05243_;
	assign _05245_ = _02024_ | ~_01398_;
	assign _05246_ = _01410_ & ~_05245_;
	assign _05247_ = \mchip.design.owner.tokens [72] & ~_05246_;
	assign _05248_ = _05247_ | _05244_;
	assign _00081_ = (_05827_ ? _05242_ : _05248_);
	assign _05250_ = _02032_ | ~_01261_;
	assign _05251_ = _01243_ & ~_05250_;
	assign _05252_ = \mchip.design.owner.tokens [73] & ~_05209_;
	assign _05253_ = _05252_ | _05251_;
	assign _05254_ = _02040_ | ~_01288_;
	assign _05255_ = _01274_ & ~_05254_;
	assign _05256_ = \mchip.design.owner.tokens [73] & ~_05215_;
	assign _05257_ = _05256_ | _05255_;
	assign _05258_ = (_00199_ ? _05253_ : _05257_);
	assign _05259_ = _02049_ | ~_01318_;
	assign _05261_ = _01303_ & ~_05259_;
	assign _05262_ = \mchip.design.owner.tokens [73] & ~_05223_;
	assign _05263_ = _05262_ | _05261_;
	assign _05264_ = (_00131_ ? _05258_ : _05263_);
	assign _05265_ = _02058_ | ~_01346_;
	assign _05266_ = _01349_ & ~_05265_;
	assign _05267_ = \mchip.design.owner.tokens [73] & ~_05231_;
	assign _05268_ = _05267_ | _05266_;
	assign _05269_ = (_06005_ ? _05264_ : _05268_);
	assign _05270_ = _02067_ | ~_01380_;
	assign _05272_ = _01382_ & ~_05270_;
	assign _05273_ = \mchip.design.owner.tokens [73] & ~_05238_;
	assign _05274_ = _05273_ | _05272_;
	assign _05275_ = (_05934_ ? _05269_ : _05274_);
	assign _05276_ = _02076_ | ~_01398_;
	assign _05277_ = _01410_ & ~_05276_;
	assign _05278_ = \mchip.design.owner.tokens [73] & ~_05246_;
	assign _05279_ = _05278_ | _05277_;
	assign _00082_ = (_05827_ ? _05275_ : _05279_);
	assign _05280_ = _02083_ | ~_01261_;
	assign _05282_ = _01243_ & ~_05280_;
	assign _05283_ = _02088_ | ~_01261_;
	assign _05284_ = _01243_ & ~_05283_;
	assign _05285_ = \mchip.design.owner.tokens [74] & ~_05284_;
	assign _05286_ = _05285_ | _05282_;
	assign _05287_ = _02095_ | ~_01288_;
	assign _05288_ = _01274_ & ~_05287_;
	assign _05289_ = _02099_ | ~_01288_;
	assign _05290_ = _01274_ & ~_05289_;
	assign _05291_ = \mchip.design.owner.tokens [74] & ~_05290_;
	assign _05293_ = _05291_ | _05288_;
	assign _05294_ = (_00199_ ? _05286_ : _05293_);
	assign _05295_ = _02107_ | ~_01318_;
	assign _05296_ = _01303_ & ~_05295_;
	assign _05297_ = _02111_ | ~_01318_;
	assign _05298_ = _01303_ & ~_05297_;
	assign _05299_ = \mchip.design.owner.tokens [74] & ~_05298_;
	assign _05300_ = _05299_ | _05296_;
	assign _05301_ = (_00131_ ? _05294_ : _05300_);
	assign _05302_ = _02119_ | ~_01346_;
	assign _05304_ = _01349_ & ~_05302_;
	assign _05305_ = _02124_ | ~_01346_;
	assign _05306_ = _01349_ & ~_05305_;
	assign _05307_ = \mchip.design.owner.tokens [74] & ~_05306_;
	assign _05308_ = _05307_ | _05304_;
	assign _05309_ = (_06005_ ? _05301_ : _05308_);
	assign _05310_ = _02132_ | ~_01380_;
	assign _05311_ = _01382_ & ~_05310_;
	assign _05312_ = _02137_ | ~_01380_;
	assign _05313_ = _01382_ & ~_05312_;
	assign _05315_ = \mchip.design.owner.tokens [74] & ~_05313_;
	assign _05316_ = _05315_ | _05311_;
	assign _05317_ = (_05934_ ? _05309_ : _05316_);
	assign _05318_ = _02145_ | ~_01398_;
	assign _05319_ = _01410_ & ~_05318_;
	assign _05320_ = _02150_ | ~_01398_;
	assign _05321_ = _01410_ & ~_05320_;
	assign _05322_ = \mchip.design.owner.tokens [74] & ~_05321_;
	assign _05323_ = _05322_ | _05319_;
	assign _00083_ = (_05827_ ? _05317_ : _05323_);
	assign _05325_ = _02157_ | ~_01261_;
	assign _05326_ = _01243_ & ~_05325_;
	assign _05327_ = \mchip.design.owner.tokens [75] & ~_05284_;
	assign _05328_ = _05327_ | _05326_;
	assign _05329_ = _02164_ | ~_01288_;
	assign _05330_ = _01274_ & ~_05329_;
	assign _05331_ = \mchip.design.owner.tokens [75] & ~_05290_;
	assign _05332_ = _05331_ | _05330_;
	assign _05333_ = (_00199_ ? _05328_ : _05332_);
	assign _05334_ = _02172_ | ~_01318_;
	assign _05336_ = _01303_ & ~_05334_;
	assign _05337_ = \mchip.design.owner.tokens [75] & ~_05298_;
	assign _05338_ = _05337_ | _05336_;
	assign _05339_ = (_00131_ ? _05333_ : _05338_);
	assign _05340_ = _02180_ | ~_01346_;
	assign _05341_ = _01349_ & ~_05340_;
	assign _05342_ = \mchip.design.owner.tokens [75] & ~_05306_;
	assign _05343_ = _05342_ | _05341_;
	assign _05344_ = (_06005_ ? _05339_ : _05343_);
	assign _05345_ = _02188_ | ~_01380_;
	assign _05347_ = _01382_ & ~_05345_;
	assign _05348_ = \mchip.design.owner.tokens [75] & ~_05313_;
	assign _05349_ = _05348_ | _05347_;
	assign _05350_ = (_05934_ ? _05344_ : _05349_);
	assign _05351_ = _02196_ | ~_01398_;
	assign _05352_ = _01410_ & ~_05351_;
	assign _05353_ = \mchip.design.owner.tokens [75] & ~_05321_;
	assign _05354_ = _05353_ | _05352_;
	assign _00084_ = (_05827_ ? _05350_ : _05354_);
	assign _05355_ = _02203_ | ~_01261_;
	assign _05357_ = _01243_ & ~_05355_;
	assign _05358_ = _02208_ | ~_01261_;
	assign _05359_ = _01243_ & ~_05358_;
	assign _05360_ = \mchip.design.owner.tokens [76] & ~_05359_;
	assign _05361_ = _05360_ | _05357_;
	assign _05362_ = _02215_ | ~_01288_;
	assign _05363_ = _01274_ & ~_05362_;
	assign _05364_ = _02220_ | ~_01288_;
	assign _05365_ = _01274_ & ~_05364_;
	assign _05366_ = \mchip.design.owner.tokens [76] & ~_05365_;
	assign _05368_ = _05366_ | _05363_;
	assign _05369_ = (_00199_ ? _05361_ : _05368_);
	assign _05370_ = _02228_ | ~_01318_;
	assign _05371_ = _01303_ & ~_05370_;
	assign _05372_ = _02233_ | ~_01318_;
	assign _05373_ = _01303_ & ~_05372_;
	assign _05374_ = \mchip.design.owner.tokens [76] & ~_05373_;
	assign _05375_ = _05374_ | _05371_;
	assign _05376_ = (_00131_ ? _05369_ : _05375_);
	assign _05377_ = _02241_ | ~_01346_;
	assign _05379_ = _01349_ & ~_05377_;
	assign _05380_ = _02246_ | ~_01346_;
	assign _05381_ = _01349_ & ~_05380_;
	assign _05382_ = \mchip.design.owner.tokens [76] & ~_05381_;
	assign _05383_ = _05382_ | _05379_;
	assign _05384_ = (_06005_ ? _05376_ : _05383_);
	assign _05385_ = _02254_ | ~_01380_;
	assign _05386_ = _01382_ & ~_05385_;
	assign _05387_ = _02259_ | ~_01380_;
	assign _05388_ = _01382_ & ~_05387_;
	assign _05390_ = \mchip.design.owner.tokens [76] & ~_05388_;
	assign _05391_ = _05390_ | _05386_;
	assign _05392_ = (_05934_ ? _05384_ : _05391_);
	assign _05393_ = _02267_ | ~_01398_;
	assign _05394_ = _01410_ & ~_05393_;
	assign _05395_ = _02272_ | ~_01398_;
	assign _05396_ = _01410_ & ~_05395_;
	assign _05397_ = \mchip.design.owner.tokens [76] & ~_05396_;
	assign _05398_ = _05397_ | _05394_;
	assign _00085_ = (_05827_ ? _05392_ : _05398_);
	assign _05400_ = _02279_ | ~_01261_;
	assign _05401_ = _01243_ & ~_05400_;
	assign _05402_ = \mchip.design.owner.tokens [77] & ~_05359_;
	assign _05403_ = _05402_ | _05401_;
	assign _05404_ = _02286_ | ~_01288_;
	assign _05405_ = _01274_ & ~_05404_;
	assign _05406_ = \mchip.design.owner.tokens [77] & ~_05365_;
	assign _05407_ = _05406_ | _05405_;
	assign _05408_ = (_00199_ ? _05403_ : _05407_);
	assign _05409_ = _02294_ | ~_01318_;
	assign _05411_ = _01303_ & ~_05409_;
	assign _05412_ = \mchip.design.owner.tokens [77] & ~_05373_;
	assign _05413_ = _05412_ | _05411_;
	assign _05414_ = (_00131_ ? _05408_ : _05413_);
	assign _05415_ = _02302_ | ~_01346_;
	assign _05416_ = _01349_ & ~_05415_;
	assign _05417_ = \mchip.design.owner.tokens [77] & ~_05381_;
	assign _05418_ = _05417_ | _05416_;
	assign _05419_ = (_06005_ ? _05414_ : _05418_);
	assign _05420_ = _02310_ | ~_01380_;
	assign _05422_ = _01382_ & ~_05420_;
	assign _05423_ = \mchip.design.owner.tokens [77] & ~_05388_;
	assign _05424_ = _05423_ | _05422_;
	assign _05425_ = (_05934_ ? _05419_ : _05424_);
	assign _05426_ = _02318_ | ~_01398_;
	assign _05427_ = _01410_ & ~_05426_;
	assign _05428_ = \mchip.design.owner.tokens [77] & ~_05396_;
	assign _05429_ = _05428_ | _05427_;
	assign _00086_ = (_05827_ ? _05425_ : _05429_);
	assign _05430_ = _02325_ | ~_01261_;
	assign _05432_ = _01243_ & ~_05430_;
	assign _05433_ = _02330_ | ~_01261_;
	assign _05434_ = _01243_ & ~_05433_;
	assign _05435_ = \mchip.design.owner.tokens [78] & ~_05434_;
	assign _05436_ = _05435_ | _05432_;
	assign _05437_ = _02337_ | ~_01288_;
	assign _05438_ = _01274_ & ~_05437_;
	assign _05439_ = _02342_ | ~_01288_;
	assign _05440_ = _01274_ & ~_05439_;
	assign _05441_ = \mchip.design.owner.tokens [78] & ~_05440_;
	assign _05443_ = _05441_ | _05438_;
	assign _05444_ = (_00199_ ? _05436_ : _05443_);
	assign _05445_ = _02350_ | ~_01318_;
	assign _05446_ = _01303_ & ~_05445_;
	assign _05447_ = _02355_ | ~_01318_;
	assign _05448_ = _01303_ & ~_05447_;
	assign _05449_ = \mchip.design.owner.tokens [78] & ~_05448_;
	assign _05450_ = _05449_ | _05446_;
	assign _05451_ = (_00131_ ? _05444_ : _05450_);
	assign _05452_ = _02363_ | ~_01346_;
	assign _05454_ = _01349_ & ~_05452_;
	assign _05455_ = _02368_ | ~_01346_;
	assign _05456_ = _01349_ & ~_05455_;
	assign _05457_ = \mchip.design.owner.tokens [78] & ~_05456_;
	assign _05458_ = _05457_ | _05454_;
	assign _05459_ = (_06005_ ? _05451_ : _05458_);
	assign _05460_ = _02376_ | ~_01380_;
	assign _05461_ = _01382_ & ~_05460_;
	assign _05462_ = _02381_ | ~_01380_;
	assign _05463_ = _01382_ & ~_05462_;
	assign _05465_ = \mchip.design.owner.tokens [78] & ~_05463_;
	assign _05466_ = _05465_ | _05461_;
	assign _05467_ = (_05934_ ? _05459_ : _05466_);
	assign _05468_ = _02389_ | ~_01398_;
	assign _05469_ = _01410_ & ~_05468_;
	assign _05470_ = _02394_ | ~_01398_;
	assign _05471_ = _01410_ & ~_05470_;
	assign _05472_ = \mchip.design.owner.tokens [78] & ~_05471_;
	assign _05473_ = _05472_ | _05469_;
	assign _00087_ = (_05827_ ? _05467_ : _05473_);
	assign _05475_ = _02401_ | ~_01261_;
	assign _05476_ = _01243_ & ~_05475_;
	assign _05477_ = \mchip.design.owner.tokens [79] & ~_05434_;
	assign _05478_ = _05477_ | _05476_;
	assign _05479_ = _02408_ | ~_01288_;
	assign _05480_ = _01274_ & ~_05479_;
	assign _05481_ = \mchip.design.owner.tokens [79] & ~_05440_;
	assign _05482_ = _05481_ | _05480_;
	assign _05483_ = (_00199_ ? _05478_ : _05482_);
	assign _05484_ = _02416_ | ~_01318_;
	assign _05486_ = _01303_ & ~_05484_;
	assign _05487_ = \mchip.design.owner.tokens [79] & ~_05448_;
	assign _05488_ = _05487_ | _05486_;
	assign _05489_ = (_00131_ ? _05483_ : _05488_);
	assign _05490_ = _02424_ | ~_01346_;
	assign _05491_ = _01349_ & ~_05490_;
	assign _05492_ = \mchip.design.owner.tokens [79] & ~_05456_;
	assign _05493_ = _05492_ | _05491_;
	assign _05494_ = (_06005_ ? _05489_ : _05493_);
	assign _05495_ = _02432_ | ~_01380_;
	assign _05496_ = _01382_ & ~_05495_;
	assign _05497_ = \mchip.design.owner.tokens [79] & ~_05463_;
	assign _05498_ = _05497_ | _05496_;
	assign _05499_ = (_05934_ ? _05494_ : _05498_);
	assign _05500_ = _02440_ | ~_01398_;
	assign _05501_ = _01410_ & ~_05500_;
	assign _05502_ = \mchip.design.owner.tokens [79] & ~_05471_;
	assign _05503_ = _05502_ | _05501_;
	assign _00088_ = (_05827_ ? _05499_ : _05503_);
	assign _05504_ = _02447_ | ~_01261_;
	assign _05506_ = _01243_ & ~_05504_;
	assign _05507_ = _02451_ | ~_01261_;
	assign _05508_ = _01243_ & ~_05507_;
	assign _05509_ = \mchip.design.owner.tokens [80] & ~_05508_;
	assign _05510_ = _05509_ | _05506_;
	assign _05511_ = _02458_ | ~_01288_;
	assign _05512_ = _01274_ & ~_05511_;
	assign _05513_ = _02462_ | ~_01288_;
	assign _05514_ = _01274_ & ~_05513_;
	assign _05515_ = \mchip.design.owner.tokens [80] & ~_05514_;
	assign _05517_ = _05515_ | _05512_;
	assign _05518_ = (_00199_ ? _05510_ : _05517_);
	assign _05519_ = _02470_ | ~_01318_;
	assign _05520_ = _01303_ & ~_05519_;
	assign _05521_ = _02475_ | ~_01318_;
	assign _05522_ = _01303_ & ~_05521_;
	assign _05523_ = \mchip.design.owner.tokens [80] & ~_05522_;
	assign _05524_ = _05523_ | _05520_;
	assign _05525_ = (_00131_ ? _05518_ : _05524_);
	assign _05526_ = _02483_ | ~_01346_;
	assign _05528_ = _01349_ & ~_05526_;
	assign _05529_ = _02488_ | ~_01346_;
	assign _05530_ = _01349_ & ~_05529_;
	assign _05531_ = \mchip.design.owner.tokens [80] & ~_05530_;
	assign _05532_ = _05531_ | _05528_;
	assign _05533_ = (_06005_ ? _05525_ : _05532_);
	assign _05534_ = _02496_ | ~_01380_;
	assign _05535_ = _01382_ & ~_05534_;
	assign _05536_ = _02501_ | ~_01380_;
	assign _05537_ = _01382_ & ~_05536_;
	assign _05539_ = \mchip.design.owner.tokens [80] & ~_05537_;
	assign _05540_ = _05539_ | _05535_;
	assign _05541_ = (_05934_ ? _05533_ : _05540_);
	assign _05542_ = _02509_ | ~_01398_;
	assign _05543_ = _01410_ & ~_05542_;
	assign _05544_ = _02514_ | ~_01398_;
	assign _05545_ = _01410_ & ~_05544_;
	assign _05546_ = \mchip.design.owner.tokens [80] & ~_05545_;
	assign _05547_ = _05546_ | _05543_;
	assign _00090_ = (_05827_ ? _05541_ : _05547_);
	assign _05549_ = _02521_ | ~_01261_;
	assign _05550_ = _01243_ & ~_05549_;
	assign _05551_ = \mchip.design.owner.tokens [81] & ~_05508_;
	assign _05552_ = _05551_ | _05550_;
	assign _05553_ = _02528_ | ~_01288_;
	assign _05554_ = _01274_ & ~_05553_;
	assign _05555_ = \mchip.design.owner.tokens [81] & ~_05514_;
	assign _05556_ = _05555_ | _05554_;
	assign _05557_ = (_00199_ ? _05552_ : _05556_);
	assign _05558_ = _02536_ | ~_01318_;
	assign _05560_ = _01303_ & ~_05558_;
	assign _05561_ = \mchip.design.owner.tokens [81] & ~_05522_;
	assign _05562_ = _05561_ | _05560_;
	assign _05563_ = (_00131_ ? _05557_ : _05562_);
	assign _05564_ = _02544_ | ~_01346_;
	assign _05565_ = _01349_ & ~_05564_;
	assign _05566_ = \mchip.design.owner.tokens [81] & ~_05530_;
	assign _05567_ = _05566_ | _05565_;
	assign _05568_ = (_06005_ ? _05563_ : _05567_);
	assign _05569_ = _02552_ | ~_01380_;
	assign _05571_ = _01382_ & ~_05569_;
	assign _05572_ = \mchip.design.owner.tokens [81] & ~_05537_;
	assign _05573_ = _05572_ | _05571_;
	assign _05574_ = (_05934_ ? _05568_ : _05573_);
	assign _05575_ = _02560_ | ~_01398_;
	assign _05576_ = _01410_ & ~_05575_;
	assign _05577_ = \mchip.design.owner.tokens [81] & ~_05545_;
	assign _05578_ = _05577_ | _05576_;
	assign _00091_ = (_05827_ ? _05574_ : _05578_);
	assign _05579_ = _02566_ | ~_01261_;
	assign _05581_ = _01243_ & ~_05579_;
	assign _05582_ = _02570_ | ~_01261_;
	assign _05583_ = _01243_ & ~_05582_;
	assign _05584_ = \mchip.design.owner.tokens [82] & ~_05583_;
	assign _05585_ = _05584_ | _05581_;
	assign _05586_ = _02576_ | ~_01288_;
	assign _05587_ = _01274_ & ~_05586_;
	assign _05588_ = _02580_ | ~_01288_;
	assign _05589_ = _01274_ & ~_05588_;
	assign _05590_ = \mchip.design.owner.tokens [82] & ~_05589_;
	assign _05592_ = _05590_ | _05587_;
	assign _05593_ = (_00199_ ? _05585_ : _05592_);
	assign _05594_ = _02587_ | ~_01318_;
	assign _05595_ = _01303_ & ~_05594_;
	assign _05596_ = _02591_ | ~_01318_;
	assign _05597_ = _01303_ & ~_05596_;
	assign _05598_ = \mchip.design.owner.tokens [82] & ~_05597_;
	assign _05599_ = _05598_ | _05595_;
	assign _05600_ = (_00131_ ? _05593_ : _05599_);
	assign _05601_ = _02598_ | ~_01346_;
	assign _05603_ = _01349_ & ~_05601_;
	assign _05604_ = _02602_ | ~_01346_;
	assign _05605_ = _01349_ & ~_05604_;
	assign _05606_ = \mchip.design.owner.tokens [82] & ~_05605_;
	assign _05607_ = _05606_ | _05603_;
	assign _05608_ = (_06005_ ? _05600_ : _05607_);
	assign _05609_ = _02609_ | ~_01380_;
	assign _05610_ = _01382_ & ~_05609_;
	assign _05611_ = _02613_ | ~_01380_;
	assign _05612_ = _01382_ & ~_05611_;
	assign _05614_ = \mchip.design.owner.tokens [82] & ~_05612_;
	assign _05615_ = _05614_ | _05610_;
	assign _05616_ = (_05934_ ? _05608_ : _05615_);
	assign _05617_ = _02620_ | ~_01398_;
	assign _05618_ = _01410_ & ~_05617_;
	assign _05619_ = _02624_ | ~_01398_;
	assign _05620_ = _01410_ & ~_05619_;
	assign _05621_ = \mchip.design.owner.tokens [82] & ~_05620_;
	assign _05622_ = _05621_ | _05618_;
	assign _00092_ = (_05827_ ? _05616_ : _05622_);
	assign _05624_ = _02630_ | ~_01261_;
	assign _05625_ = _01243_ & ~_05624_;
	assign _05626_ = \mchip.design.owner.tokens [83] & ~_05583_;
	assign _05627_ = _05626_ | _05625_;
	assign _05628_ = _02636_ | ~_01288_;
	assign _05629_ = _01274_ & ~_05628_;
	assign _05630_ = \mchip.design.owner.tokens [83] & ~_05589_;
	assign _05631_ = _05630_ | _05629_;
	assign _05632_ = (_00199_ ? _05627_ : _05631_);
	assign _05633_ = _02643_ | ~_01318_;
	assign _05635_ = _01303_ & ~_05633_;
	assign _05636_ = \mchip.design.owner.tokens [83] & ~_05597_;
	assign _05637_ = _05636_ | _05635_;
	assign _05638_ = (_00131_ ? _05632_ : _05637_);
	assign _05639_ = _02650_ | ~_01346_;
	assign _05640_ = _01349_ & ~_05639_;
	assign _05641_ = \mchip.design.owner.tokens [83] & ~_05605_;
	assign _05642_ = _05641_ | _05640_;
	assign _05643_ = (_06005_ ? _05638_ : _05642_);
	assign _05644_ = _02657_ | ~_01380_;
	assign _05646_ = _01382_ & ~_05644_;
	assign _05647_ = \mchip.design.owner.tokens [83] & ~_05612_;
	assign _05648_ = _05647_ | _05646_;
	assign _05649_ = (_05934_ ? _05643_ : _05648_);
	assign _05650_ = _02665_ | ~_01398_;
	assign _05651_ = _01410_ & ~_05650_;
	assign _05652_ = \mchip.design.owner.tokens [83] & ~_05620_;
	assign _05653_ = _05652_ | _05651_;
	assign _00093_ = (_05827_ ? _05649_ : _05653_);
	assign _06061_[0] = ~\mchip.design.vga.h_idx [0];
	assign _05655_ = _00449_ | _00303_;
	assign _05656_ = _00297_ & ~_05655_;
	assign _05657_ = ~_00308_;
	assign _05658_ = ~_00305_;
	assign _05659_ = ~(_00315_ & _00298_);
	assign _05660_ = _05659_ & ~_00303_;
	assign _05661_ = _05658_ & ~_05660_;
	assign _05662_ = _00297_ & ~_05661_;
	assign _05663_ = _05657_ & ~_05662_;
	assign _05664_ = _05663_ | _05656_;
	assign _05666_ = ~(_00828_ | _00303_);
	assign _05667_ = ~(_05666_ & _00297_);
	assign _05668_ = ~(_00832_ | _00303_);
	assign _05669_ = _05658_ & ~_05668_;
	assign _05670_ = _00297_ & ~_05669_;
	assign _05671_ = _05657_ & ~_05670_;
	assign _05672_ = _05667_ & ~_05671_;
	assign _00107_ = _05672_ | _05664_;
	assign _05673_ = _00505_ & ~_00533_;
	assign _05674_ = _05673_ | _03750_;
	assign _05676_ = _00564_ | _00509_;
	assign _05677_ = _05676_ | _03814_;
	assign _05678_ = _05677_ | ~_00505_;
	assign _05679_ = ~(_00599_ | _00564_);
	assign _05680_ = _00532_ & ~_05679_;
	assign _05681_ = _00505_ & ~_05680_;
	assign _05682_ = _05681_ | _03750_;
	assign _05683_ = _05678_ & ~_05682_;
	assign _00096_ = _05683_ | _05674_;
	assign _06065_[1] = \mchip.design.pve.fsm.timeOut [1] ^ \mchip.design.pve.fsm.timeOut [0];
	assign _05685_ = \mchip.design.pve.fsm.timeOut [1] & \mchip.design.pve.fsm.timeOut [0];
	assign _06065_[2] = _05685_ ^ \mchip.design.pve.fsm.timeOut [2];
	assign _05686_ = _05685_ & \mchip.design.pve.fsm.timeOut [2];
	assign _06065_[3] = _05686_ ^ \mchip.design.pve.fsm.timeOut [3];
	assign _05687_ = ~(\mchip.design.pve.fsm.timeOut [2] & \mchip.design.pve.fsm.timeOut [3]);
	assign _05688_ = _05685_ & ~_05687_;
	assign _06065_[4] = _05688_ ^ \mchip.design.pve.fsm.timeOut [4];
	assign _05689_ = _05688_ & \mchip.design.pve.fsm.timeOut [4];
	assign _06065_[5] = _05689_ ^ \mchip.design.pve.fsm.timeOut [5];
	assign _05690_ = ~(\mchip.design.pve.fsm.timeOut [5] & \mchip.design.pve.fsm.timeOut [4]);
	assign _05692_ = _05688_ & ~_05690_;
	assign _06065_[6] = _05692_ ^ \mchip.design.pve.fsm.timeOut [6];
	assign _05693_ = _05692_ & \mchip.design.pve.fsm.timeOut [6];
	assign _06065_[7] = _05693_ ^ \mchip.design.pve.fsm.timeOut [7];
	assign _05694_ = ~(\mchip.design.pve.fsm.timeOut [6] & \mchip.design.pve.fsm.timeOut [7]);
	assign _05695_ = ~(_05694_ | _05690_);
	assign _05696_ = ~(_05695_ & _05688_);
	assign _06065_[8] = ~(_05696_ ^ \mchip.design.pve.fsm.timeOut [8]);
	assign _05697_ = \mchip.design.pve.fsm.timeOut [8] & ~_05696_;
	assign _06065_[9] = _05697_ ^ \mchip.design.pve.fsm.timeOut [9];
	assign _05699_ = ~(_05696_ | _02953_);
	assign _06065_[10] = _05699_ ^ \mchip.design.pve.fsm.timeOut [10];
	assign _05700_ = _05699_ & \mchip.design.pve.fsm.timeOut [10];
	assign _06065_[11] = _05700_ ^ \mchip.design.pve.fsm.timeOut [11];
	assign _05701_ = ~(_05696_ | _02964_);
	assign _06065_[12] = _05701_ ^ \mchip.design.pve.fsm.timeOut [12];
	assign _05702_ = _05701_ & \mchip.design.pve.fsm.timeOut [12];
	assign _06065_[13] = _05702_ ^ \mchip.design.pve.fsm.timeOut [13];
	assign _05703_ = ~(\mchip.design.pve.fsm.timeOut [12] & \mchip.design.pve.fsm.timeOut [13]);
	assign _05704_ = _05701_ & ~_05703_;
	assign _06065_[14] = _05704_ ^ \mchip.design.pve.fsm.timeOut [14];
	assign _05706_ = _05704_ & \mchip.design.pve.fsm.timeOut [14];
	assign _06065_[15] = _05706_ ^ \mchip.design.pve.fsm.timeOut [15];
	assign _05707_ = ~(\mchip.design.pve.fsm.timeOut [14] & \mchip.design.pve.fsm.timeOut [15]);
	assign _05708_ = _05707_ | _05703_;
	assign _05709_ = _05708_ | _02964_;
	assign _05710_ = _05709_ | _05696_;
	assign _06065_[16] = ~(_05710_ ^ \mchip.design.pve.fsm.timeOut [16]);
	assign _05711_ = \mchip.design.pve.fsm.timeOut [16] & ~_05710_;
	assign _06065_[17] = _05711_ ^ \mchip.design.pve.fsm.timeOut [17];
	assign _05713_ = _02693_ & ~_05710_;
	assign _06065_[18] = _05713_ ^ \mchip.design.pve.fsm.timeOut [18];
	assign _05714_ = _05713_ & \mchip.design.pve.fsm.timeOut [18];
	assign _06065_[19] = _05714_ ^ \mchip.design.pve.fsm.timeOut [19];
	assign _05715_ = ~(_05710_ | _02715_);
	assign _06065_[20] = _05715_ ^ \mchip.design.pve.fsm.timeOut [20];
	assign _05716_ = _05715_ & \mchip.design.pve.fsm.timeOut [20];
	assign _06065_[21] = _05716_ ^ \mchip.design.pve.fsm.timeOut [21];
	assign _05717_ = ~(\mchip.design.pve.fsm.timeOut [21] & \mchip.design.pve.fsm.timeOut [20]);
	assign _05718_ = _05715_ & ~_05717_;
	assign _06065_[22] = _05718_ ^ \mchip.design.pve.fsm.timeOut [22];
	assign _06066_[2] = ~(_00511_ ^ \mchip.design.vga.h_idx [2]);
	assign _05720_ = \mchip.design.vga.h_idx [2] & ~_00511_;
	assign _06066_[3] = _05720_ ^ \mchip.design.vga.h_idx [3];
	assign _06066_[4] = _00524_ ^ \mchip.design.vga.h_idx [4];
	assign _05721_ = _00524_ & ~_00548_;
	assign _06066_[5] = _05721_ ^ \mchip.design.vga.h_idx [5];
	assign _05722_ = _00524_ & _00521_;
	assign _06066_[6] = _05722_ ^ \mchip.design.vga.h_idx [6];
	assign _05723_ = _05722_ & \mchip.design.vga.h_idx [6];
	assign _06066_[7] = _05723_ ^ \mchip.design.vga.h_idx [7];
	assign _06066_[8] = _00616_ ^ \mchip.design.vga.h_idx [8];
	assign _05725_ = _00616_ & \mchip.design.vga.h_idx [8];
	assign _06066_[9] = _05725_ ^ \mchip.design.vga.h_idx [9];
	assign _06061_[1] = ~(_00562_ & _00530_);
	assign _05726_ = _03697_ | ~_03686_;
	assign _00001_ = \mchip.design.pve.fsm.currState [0] & ~_05726_;
	assign _05727_ = io_in[13] | ~\mchip.design.inputConfirmSync ;
	assign _00000_ = \mchip.design.currStateConfirm [0] & ~_05727_;
	assign \mchip.design.pve.rand0.inputFF [0] = \mchip.design.pve.rand0.outputFF [2] ^ \mchip.design.pve.rand0.outputFF [3];
	assign _06063_[1] = \mchip.design.debounceCount [0] ^ \mchip.design.debounceCount [1];
	assign _05729_ = \mchip.design.debounceCount [0] & \mchip.design.debounceCount [1];
	assign _06063_[2] = _05729_ ^ \mchip.design.debounceCount [2];
	assign _05730_ = _05729_ & \mchip.design.debounceCount [2];
	assign _06063_[3] = _05730_ ^ \mchip.design.debounceCount [3];
	assign _05731_ = ~(\mchip.design.debounceCount [2] & \mchip.design.debounceCount [3]);
	assign _05732_ = _05729_ & ~_05731_;
	assign _06063_[4] = _05732_ ^ \mchip.design.debounceCount [4];
	assign _05733_ = _05732_ & \mchip.design.debounceCount [4];
	assign _06063_[5] = _05733_ ^ \mchip.design.debounceCount [5];
	assign _05735_ = ~(\mchip.design.debounceCount [5] & \mchip.design.debounceCount [4]);
	assign _05736_ = _05732_ & ~_05735_;
	assign _06063_[6] = _05736_ ^ \mchip.design.debounceCount [6];
	assign _05737_ = _05736_ & \mchip.design.debounceCount [6];
	assign _06063_[7] = _05737_ ^ \mchip.design.debounceCount [7];
	assign _05738_ = ~(\mchip.design.debounceCount [6] & \mchip.design.debounceCount [7]);
	assign _05739_ = ~(_05738_ | _05735_);
	assign _05740_ = ~(_05739_ & _05732_);
	assign _06063_[8] = ~(_05740_ ^ \mchip.design.debounceCount [8]);
	assign _05741_ = \mchip.design.debounceCount [8] & ~_05740_;
	assign _06063_[9] = _05741_ ^ \mchip.design.debounceCount [9];
	assign _05743_ = ~(_05740_ | _00276_);
	assign _06063_[10] = _05743_ ^ \mchip.design.debounceCount [10];
	assign _05744_ = _05743_ & \mchip.design.debounceCount [10];
	assign _06063_[11] = _05744_ ^ \mchip.design.debounceCount [11];
	assign _05745_ = ~(_05740_ | _00277_);
	assign _06063_[12] = _05745_ ^ \mchip.design.debounceCount [12];
	assign _05746_ = _05745_ & \mchip.design.debounceCount [12];
	assign _06063_[13] = _05746_ ^ \mchip.design.debounceCount [13];
	assign _05747_ = ~(\mchip.design.debounceCount [12] & \mchip.design.debounceCount [13]);
	assign _05749_ = _05745_ & ~_05747_;
	assign _06063_[14] = _05749_ ^ \mchip.design.debounceCount [14];
	assign _05750_ = _05749_ & \mchip.design.debounceCount [14];
	assign _06063_[15] = _05750_ ^ \mchip.design.debounceCount [15];
	assign _05751_ = ~(\mchip.design.debounceCount [14] & \mchip.design.debounceCount [15]);
	assign _05752_ = _05751_ | _05747_;
	assign _05753_ = _05752_ | _00277_;
	assign _05754_ = _05753_ | _05740_;
	assign _06063_[16] = ~(_05754_ ^ \mchip.design.debounceCount [16]);
	assign _05755_ = \mchip.design.debounceCount [16] & ~_05754_;
	assign _06063_[17] = _05755_ ^ \mchip.design.debounceCount [17];
	assign _05757_ = _00252_ & ~_05754_;
	assign _06063_[18] = _05757_ ^ \mchip.design.debounceCount [18];
	assign _05758_ = _05757_ & \mchip.design.debounceCount [18];
	assign _06063_[19] = _05758_ ^ \mchip.design.debounceCount [19];
	assign _05759_ = ~(_05754_ | _00254_);
	assign _06063_[20] = _05759_ ^ \mchip.design.debounceCount [20];
	assign _05760_ = _05759_ & \mchip.design.debounceCount [20];
	assign _06063_[21] = _05760_ ^ \mchip.design.debounceCount [21];
	assign _05761_ = ~(\mchip.design.debounceCount [21] & \mchip.design.debounceCount [20]);
	assign _05762_ = _05759_ & ~_05761_;
	assign _06063_[22] = _05762_ ^ \mchip.design.debounceCount [22];
	assign \mchip.design.pve.rand6.inputFF [0] = \mchip.design.pve.rand6.outputFF [2] ^ \mchip.design.pve.rand6.outputFF [3];
	assign \mchip.design.pve.rand5.inputFF [0] = \mchip.design.pve.rand5.outputFF [2] ^ \mchip.design.pve.rand5.outputFF [3];
	assign \mchip.design.pve.rand4.inputFF [0] = \mchip.design.pve.rand4.outputFF [2] ^ \mchip.design.pve.rand4.outputFF [3];
	assign \mchip.design.pve.rand3.inputFF [0] = \mchip.design.pve.rand3.outputFF [2] ^ \mchip.design.pve.rand3.outputFF [3];
	assign \mchip.design.pve.rand2.inputFF [0] = \mchip.design.pve.rand2.outputFF [2] ^ \mchip.design.pve.rand2.outputFF [3];
	assign \mchip.design.pve.rand1.inputFF [0] = \mchip.design.pve.rand1.outputFF [2] ^ \mchip.design.pve.rand1.outputFF [3];
	always @(posedge io_in[12]) \mchip.design.currStateConfirm [0] <= _00002_;
	always @(posedge io_in[12]) \mchip.design.currStateConfirm [1] <= _00000_;
	always @(posedge io_in[12]) \mchip.design.currStateConfirm [2] <= _00003_;
	always @(posedge io_in[12]) \mchip.design.pve.fsm.currState [0] <= _00004_;
	always @(posedge io_in[12]) \mchip.design.pve.fsm.currState [1] <= _00005_;
	always @(posedge io_in[12]) \mchip.design.pve.fsm.currState [2] <= _00001_;
	always @(posedge io_in[12]) \mchip.design.inputNewGameSync  <= \mchip.design.inputNewGameHalf ;
	always @(posedge io_in[12]) \mchip.design.inputNewGameHalf  <= io_in[10];
	always @(posedge io_in[12]) \mchip.design.inputMovesHalf [0] <= io_in[0];
	always @(posedge io_in[12]) \mchip.design.inputMovesHalf [1] <= io_in[1];
	always @(posedge io_in[12]) \mchip.design.inputMovesHalf [2] <= io_in[2];
	always @(posedge io_in[12]) \mchip.design.inputMovesHalf [3] <= io_in[3];
	always @(posedge io_in[12]) \mchip.design.inputMovesHalf [4] <= io_in[4];
	always @(posedge io_in[12]) \mchip.design.inputMovesHalf [5] <= io_in[5];
	always @(posedge io_in[12]) \mchip.design.inputMovesHalf [6] <= io_in[6];
	always @(posedge io_in[12]) \mchip.design.inputMovesSync [0] <= \mchip.design.inputMovesHalf [0];
	always @(posedge io_in[12]) \mchip.design.inputMovesSync [1] <= \mchip.design.inputMovesHalf [1];
	always @(posedge io_in[12]) \mchip.design.inputMovesSync [2] <= \mchip.design.inputMovesHalf [2];
	always @(posedge io_in[12]) \mchip.design.inputMovesSync [3] <= \mchip.design.inputMovesHalf [3];
	always @(posedge io_in[12]) \mchip.design.inputMovesSync [4] <= \mchip.design.inputMovesHalf [4];
	always @(posedge io_in[12]) \mchip.design.inputMovesSync [5] <= \mchip.design.inputMovesHalf [5];
	always @(posedge io_in[12]) \mchip.design.inputMovesSync [6] <= \mchip.design.inputMovesHalf [6];
	always @(posedge io_in[12]) \mchip.design.inputConfirmHalf  <= io_in[7];
	always @(posedge io_in[12]) \mchip.design.inputConfirmSync  <= \mchip.design.inputConfirmHalf ;
	always @(posedge io_in[12]) \mchip.design.inputSwitchPlayerHalf  <= io_in[8];
	always @(posedge io_in[12]) \mchip.design.inputSwitchPlayerSync  <= \mchip.design.inputSwitchPlayerHalf ;
	always @(posedge io_in[12]) \mchip.design.inputSwitchPVPHalf  <= io_in[9];
	always @(posedge io_in[12]) \mchip.design.inputSwitchPVPSync  <= \mchip.design.inputSwitchPVPHalf ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.hsync  <= 1'h1;
		else
			\mchip.design.vga.hsync  <= _00096_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [0] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [0] <= _00097_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [1] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [1] <= _00098_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [2] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [2] <= _00099_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [3] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [3] <= _00100_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [4] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [4] <= _00101_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [5] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [5] <= _00102_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [6] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [6] <= _00103_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [7] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [7] <= _00104_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [8] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [8] <= _00105_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.v_idx [9] <= 1'h0;
		else if (_00011_)
			\mchip.design.vga.v_idx [9] <= _00106_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.vga.vsync  <= 1'h1;
		else if (_00011_)
			\mchip.design.vga.vsync  <= _00107_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand6.outputFF [0] <= 1'h1;
		else
			\mchip.design.pve.rand6.outputFF [0] <= \mchip.design.pve.rand6.inputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand6.outputFF [1] <= 1'h0;
		else
			\mchip.design.pve.rand6.outputFF [1] <= \mchip.design.pve.rand6.outputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand6.outputFF [2] <= 1'h1;
		else
			\mchip.design.pve.rand6.outputFF [2] <= \mchip.design.pve.rand6.outputFF [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand6.outputFF [3] <= 1'h0;
		else
			\mchip.design.pve.rand6.outputFF [3] <= \mchip.design.pve.rand6.outputFF [2];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [0] <= 1'h0;
		else
			\mchip.design.debounceCount [0] <= _06062_[0];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [1] <= 1'h0;
		else
			\mchip.design.debounceCount [1] <= _06063_[1];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [2] <= 1'h0;
		else
			\mchip.design.debounceCount [2] <= _06063_[2];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [3] <= 1'h0;
		else
			\mchip.design.debounceCount [3] <= _06063_[3];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [4] <= 1'h0;
		else
			\mchip.design.debounceCount [4] <= _06063_[4];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [5] <= 1'h0;
		else
			\mchip.design.debounceCount [5] <= _06063_[5];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [6] <= 1'h0;
		else
			\mchip.design.debounceCount [6] <= _06063_[6];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [7] <= 1'h0;
		else
			\mchip.design.debounceCount [7] <= _06063_[7];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [8] <= 1'h0;
		else
			\mchip.design.debounceCount [8] <= _06063_[8];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [9] <= 1'h0;
		else
			\mchip.design.debounceCount [9] <= _06063_[9];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [10] <= 1'h0;
		else
			\mchip.design.debounceCount [10] <= _06063_[10];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [11] <= 1'h0;
		else
			\mchip.design.debounceCount [11] <= _06063_[11];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [12] <= 1'h0;
		else
			\mchip.design.debounceCount [12] <= _06063_[12];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [13] <= 1'h0;
		else
			\mchip.design.debounceCount [13] <= _06063_[13];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [14] <= 1'h0;
		else
			\mchip.design.debounceCount [14] <= _06063_[14];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [15] <= 1'h0;
		else
			\mchip.design.debounceCount [15] <= _06063_[15];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [16] <= 1'h0;
		else
			\mchip.design.debounceCount [16] <= _06063_[16];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [17] <= 1'h0;
		else
			\mchip.design.debounceCount [17] <= _06063_[17];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [18] <= 1'h0;
		else
			\mchip.design.debounceCount [18] <= _06063_[18];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [19] <= 1'h0;
		else
			\mchip.design.debounceCount [19] <= _06063_[19];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [20] <= 1'h0;
		else
			\mchip.design.debounceCount [20] <= _06063_[20];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [21] <= 1'h0;
		else
			\mchip.design.debounceCount [21] <= _06063_[21];
	always @(posedge io_in[12])
		if (_00010_)
			\mchip.design.debounceCount [22] <= 1'h0;
		else
			\mchip.design.debounceCount [22] <= _06063_[22];
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [0] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [0] <= _00012_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [1] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [1] <= _00023_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [2] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [2] <= _00034_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [3] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [3] <= _00045_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [4] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [4] <= _00056_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [5] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [5] <= _00067_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [6] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [6] <= _00078_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [7] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [7] <= _00089_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [8] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [8] <= _00094_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [9] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [9] <= _00095_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [10] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [10] <= _00013_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [11] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [11] <= _00014_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [12] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [12] <= _00015_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [13] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [13] <= _00016_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [14] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [14] <= _00017_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [15] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [15] <= _00018_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [16] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [16] <= _00019_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [17] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [17] <= _00020_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [18] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [18] <= _00021_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [19] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [19] <= _00022_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [20] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [20] <= _00024_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [21] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [21] <= _00025_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [22] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [22] <= _00026_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [23] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [23] <= _00027_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [24] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [24] <= _00028_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [25] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [25] <= _00029_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [26] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [26] <= _00030_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [27] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [27] <= _00031_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [28] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [28] <= _00032_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [29] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [29] <= _00033_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [30] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [30] <= _00035_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [31] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [31] <= _00036_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [32] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [32] <= _00037_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [33] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [33] <= _00038_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [34] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [34] <= _00039_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [35] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [35] <= _00040_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [36] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [36] <= _00041_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [37] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [37] <= _00042_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [38] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [38] <= _00043_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [39] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [39] <= _00044_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [40] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [40] <= _00046_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [41] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [41] <= _00047_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [42] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [42] <= _00048_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [43] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [43] <= _00049_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [44] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [44] <= _00050_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [45] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [45] <= _00051_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [46] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [46] <= _00052_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [47] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [47] <= _00053_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [48] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [48] <= _00054_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [49] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [49] <= _00055_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [50] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [50] <= _00057_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [51] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [51] <= _00058_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [52] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [52] <= _00059_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [53] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [53] <= _00060_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [54] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [54] <= _00061_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [55] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [55] <= _00062_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [56] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [56] <= _00063_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [57] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [57] <= _00064_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [58] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [58] <= _00065_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [59] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [59] <= _00066_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [60] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [60] <= _00068_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [61] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [61] <= _00069_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [62] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [62] <= _00070_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [63] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [63] <= _00071_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [64] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [64] <= _00072_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [65] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [65] <= _00073_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [66] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [66] <= _00074_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [67] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [67] <= _00075_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [68] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [68] <= _00076_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [69] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [69] <= _00077_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [70] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [70] <= _00079_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [71] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [71] <= _00080_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [72] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [72] <= _00081_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [73] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [73] <= _00082_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [74] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [74] <= _00083_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [75] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [75] <= _00084_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [76] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [76] <= _00085_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [77] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [77] <= _00086_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [78] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [78] <= _00087_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [79] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [79] <= _00088_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [80] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [80] <= _00090_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [81] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [81] <= _00091_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [82] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [82] <= _00092_;
	always @(posedge io_in[12])
		if (_00009_)
			\mchip.design.owner.tokens [83] <= 1'h0;
		else if (_00006_)
			\mchip.design.owner.tokens [83] <= _00093_;
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [0] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [0] <= _06064_[0];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [1] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [1] <= _06065_[1];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [2] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [2] <= _06065_[2];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [3] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [3] <= _06065_[3];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [4] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [4] <= _06065_[4];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [5] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [5] <= _06065_[5];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [6] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [6] <= _06065_[6];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [7] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [7] <= _06065_[7];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [8] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [8] <= _06065_[8];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [9] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [9] <= _06065_[9];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [10] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [10] <= _06065_[10];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [11] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [11] <= _06065_[11];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [12] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [12] <= _06065_[12];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [13] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [13] <= _06065_[13];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [14] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [14] <= _06065_[14];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [15] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [15] <= _06065_[15];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [16] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [16] <= _06065_[16];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [17] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [17] <= _06065_[17];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [18] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [18] <= _06065_[18];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [19] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [19] <= _06065_[19];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [20] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [20] <= _06065_[20];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [21] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [21] <= _06065_[21];
	always @(posedge io_in[12])
		if (_00008_)
			\mchip.design.pve.fsm.timeOut [22] <= 1'h0;
		else if (\mchip.design.pve.fsm.currState [1])
			\mchip.design.pve.fsm.timeOut [22] <= _06065_[22];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [0] <= 1'h0;
		else
			\mchip.design.vga.h_idx [0] <= _06061_[0];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [1] <= 1'h0;
		else
			\mchip.design.vga.h_idx [1] <= _06061_[1];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [2] <= 1'h0;
		else
			\mchip.design.vga.h_idx [2] <= _06066_[2];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [3] <= 1'h0;
		else
			\mchip.design.vga.h_idx [3] <= _06066_[3];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [4] <= 1'h0;
		else
			\mchip.design.vga.h_idx [4] <= _06066_[4];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [5] <= 1'h0;
		else
			\mchip.design.vga.h_idx [5] <= _06066_[5];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [6] <= 1'h0;
		else
			\mchip.design.vga.h_idx [6] <= _06066_[6];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [7] <= 1'h0;
		else
			\mchip.design.vga.h_idx [7] <= _06066_[7];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [8] <= 1'h0;
		else
			\mchip.design.vga.h_idx [8] <= _06066_[8];
	always @(posedge io_in[12])
		if (_00007_)
			\mchip.design.vga.h_idx [9] <= 1'h0;
		else
			\mchip.design.vga.h_idx [9] <= _06066_[9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand5.outputFF [0] <= 1'h1;
		else
			\mchip.design.pve.rand5.outputFF [0] <= \mchip.design.pve.rand5.inputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand5.outputFF [1] <= 1'h1;
		else
			\mchip.design.pve.rand5.outputFF [1] <= \mchip.design.pve.rand5.outputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand5.outputFF [2] <= 1'h0;
		else
			\mchip.design.pve.rand5.outputFF [2] <= \mchip.design.pve.rand5.outputFF [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand5.outputFF [3] <= 1'h0;
		else
			\mchip.design.pve.rand5.outputFF [3] <= \mchip.design.pve.rand5.outputFF [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand4.outputFF [0] <= 1'h1;
		else
			\mchip.design.pve.rand4.outputFF [0] <= \mchip.design.pve.rand4.inputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand4.outputFF [1] <= 1'h0;
		else
			\mchip.design.pve.rand4.outputFF [1] <= \mchip.design.pve.rand4.outputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand4.outputFF [2] <= 1'h0;
		else
			\mchip.design.pve.rand4.outputFF [2] <= \mchip.design.pve.rand4.outputFF [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand4.outputFF [3] <= 1'h1;
		else
			\mchip.design.pve.rand4.outputFF [3] <= \mchip.design.pve.rand4.outputFF [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand3.outputFF [0] <= 1'h0;
		else
			\mchip.design.pve.rand3.outputFF [0] <= \mchip.design.pve.rand3.inputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand3.outputFF [1] <= 1'h0;
		else
			\mchip.design.pve.rand3.outputFF [1] <= \mchip.design.pve.rand3.outputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand3.outputFF [2] <= 1'h1;
		else
			\mchip.design.pve.rand3.outputFF [2] <= \mchip.design.pve.rand3.outputFF [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand3.outputFF [3] <= 1'h1;
		else
			\mchip.design.pve.rand3.outputFF [3] <= \mchip.design.pve.rand3.outputFF [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand2.outputFF [0] <= 1'h1;
		else
			\mchip.design.pve.rand2.outputFF [0] <= \mchip.design.pve.rand2.inputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand2.outputFF [1] <= 1'h0;
		else
			\mchip.design.pve.rand2.outputFF [1] <= \mchip.design.pve.rand2.outputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand2.outputFF [2] <= 1'h1;
		else
			\mchip.design.pve.rand2.outputFF [2] <= \mchip.design.pve.rand2.outputFF [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand2.outputFF [3] <= 1'h1;
		else
			\mchip.design.pve.rand2.outputFF [3] <= \mchip.design.pve.rand2.outputFF [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand1.outputFF [0] <= 1'h1;
		else
			\mchip.design.pve.rand1.outputFF [0] <= \mchip.design.pve.rand1.inputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand1.outputFF [1] <= 1'h1;
		else
			\mchip.design.pve.rand1.outputFF [1] <= \mchip.design.pve.rand1.outputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand1.outputFF [2] <= 1'h0;
		else
			\mchip.design.pve.rand1.outputFF [2] <= \mchip.design.pve.rand1.outputFF [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand1.outputFF [3] <= 1'h0;
		else
			\mchip.design.pve.rand1.outputFF [3] <= \mchip.design.pve.rand1.outputFF [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand0.outputFF [0] <= 1'h1;
		else
			\mchip.design.pve.rand0.outputFF [0] <= \mchip.design.pve.rand0.inputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand0.outputFF [1] <= 1'h1;
		else
			\mchip.design.pve.rand0.outputFF [1] <= \mchip.design.pve.rand0.outputFF [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand0.outputFF [2] <= 1'h1;
		else
			\mchip.design.pve.rand0.outputFF [2] <= \mchip.design.pve.rand0.outputFF [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.pve.rand0.outputFF [3] <= 1'h1;
		else
			\mchip.design.pve.rand0.outputFF [3] <= \mchip.design.pve.rand0.outputFF [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.design.owner.fsm.currState  <= 1'h0;
		else
			\mchip.design.owner.fsm.currState  <= \mchip.design.inputSwitchPlayerSync ;
	assign _06061_[9:2] = 8'h00;
	assign _06062_[22:1] = \mchip.design.debounceCount [22:1];
	assign _06063_[0] = _06062_[0];
	assign _06064_[22:1] = \mchip.design.pve.fsm.timeOut [22:1];
	assign _06065_[0] = _06064_[0];
	assign _06066_[1:0] = _06061_[1:0];
	assign {io_out[13:8], io_out[6], io_out[4:0]} = {4'h0, \mchip.design.board.is_board , \mchip.design.board.is_board , io_out[7], io_out[5], 1'h0, \mchip.design.blank , \mchip.design.vga.hsync , \mchip.design.vga.vsync };
	assign \mchip.clock  = io_in[12];
	assign \mchip.design.HS  = \mchip.design.vga.hsync ;
	assign \mchip.design.VGA_Blue  = {\mchip.design.board.is_board , \mchip.design.board.is_board };
	assign \mchip.design.VGA_Green  = {io_out[7], io_out[7]};
	assign \mchip.design.VGA_Red  = {io_out[5], io_out[5]};
	assign \mchip.design.VS  = \mchip.design.vga.vsync ;
	assign \mchip.design.board.col  = \mchip.design.vga.h_idx ;
	assign \mchip.design.board.level_0_H.high  = 9'h01d;
	assign \mchip.design.board.level_0_H.low  = 9'h000;
	assign \mchip.design.board.level_0_H.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.board.level_0_V.high  = 10'h02c;
	assign \mchip.design.board.level_0_V.low  = 10'h000;
	assign \mchip.design.board.level_0_V.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.board.level_1_H.high  = 9'h068;
	assign \mchip.design.board.level_1_H.low  = 9'h04b;
	assign \mchip.design.board.level_1_H.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.board.level_1_V.high  = 10'h081;
	assign \mchip.design.board.level_1_V.low  = 10'h055;
	assign \mchip.design.board.level_1_V.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.board.level_2_H.high  = 9'h0b3;
	assign \mchip.design.board.level_2_H.low  = 9'h096;
	assign \mchip.design.board.level_2_H.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.board.level_2_V.high  = 10'h0d6;
	assign \mchip.design.board.level_2_V.low  = 10'h0aa;
	assign \mchip.design.board.level_2_V.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.board.level_3_H.high  = 9'h0fe;
	assign \mchip.design.board.level_3_H.low  = 9'h0e1;
	assign \mchip.design.board.level_3_H.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.board.level_3_V.high  = 10'h12b;
	assign \mchip.design.board.level_3_V.low  = 10'h0ff;
	assign \mchip.design.board.level_3_V.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.board.level_4_H.high  = 9'h149;
	assign \mchip.design.board.level_4_H.low  = 9'h12c;
	assign \mchip.design.board.level_4_H.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.board.level_4_V.high  = 10'h180;
	assign \mchip.design.board.level_4_V.low  = 10'h154;
	assign \mchip.design.board.level_4_V.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.board.level_5_H.high  = 9'h194;
	assign \mchip.design.board.level_5_H.low  = 9'h177;
	assign \mchip.design.board.level_5_H.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.board.level_5_V.high  = 10'h1d5;
	assign \mchip.design.board.level_5_V.low  = 10'h1a9;
	assign \mchip.design.board.level_5_V.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.board.level_6_H.high  = 9'h1df;
	assign \mchip.design.board.level_6_H.low  = 9'h1c2;
	assign \mchip.design.board.level_6_H.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.board.level_6_V.high  = 10'h22a;
	assign \mchip.design.board.level_6_V.low  = 10'h1fe;
	assign \mchip.design.board.level_6_V.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.board.level_7_V.high  = 10'h27f;
	assign \mchip.design.board.level_7_V.low  = 10'h253;
	assign \mchip.design.board.level_7_V.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.board.row  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.bot_confirm  = \mchip.design.pve.fsm.currState [2];
	assign \mchip.design.clock  = io_in[12];
	assign \mchip.design.colFromVGA  = \mchip.design.vga.h_idx ;
	assign \mchip.design.colToModule  = \mchip.design.vga.h_idx ;
	assign \mchip.design.colors.blue  = {\mchip.design.board.is_board , \mchip.design.board.is_board };
	assign \mchip.design.colors.clock  = io_in[12];
	assign \mchip.design.colors.currentTokenCol  = 7'h00;
	assign \mchip.design.colors.currentTokenRow  = 6'h00;
	assign \mchip.design.colors.green  = {io_out[7], io_out[7]};
	assign \mchip.design.colors.is_board  = \mchip.design.board.is_board ;
	assign \mchip.design.colors.red  = {io_out[5], io_out[5]};
	assign \mchip.design.colors.reset  = io_in[13];
	assign \mchip.design.colors.tokens  = \mchip.design.owner.tokens ;
	assign \mchip.design.debounceClear  = 1'h1;
	assign \mchip.design.debounceCountEn  = \mchip.design.currStateConfirm [2];
	assign \mchip.design.debounceLimit  = 23'h5f5e10;
	assign \mchip.design.inputChangeDebug  = io_in[11];
	assign \mchip.design.inputConfirm  = io_in[7];
	assign \mchip.design.inputConfirmLimited  = \mchip.design.currStateConfirm [1];
	assign \mchip.design.inputMoves  = io_in[6:0];
	assign \mchip.design.inputNewGame  = io_in[10];
	assign \mchip.design.inputSwitchPVP  = io_in[9];
	assign \mchip.design.inputSwitchPlayer  = io_in[8];
	assign \mchip.design.is_board  = \mchip.design.board.is_board ;
	assign \mchip.design.outputs  = {2'h0, \mchip.design.board.is_board , \mchip.design.board.is_board , io_out[7], io_out[7], io_out[5], io_out[5], 1'h0, \mchip.design.blank , \mchip.design.vga.hsync , \mchip.design.vga.vsync };
	assign \mchip.design.owner.clock  = io_in[12];
	assign \mchip.design.owner.currentPlayer  = \mchip.design.owner.fsm.currState ;
	assign \mchip.design.owner.fsm.clock  = io_in[12];
	assign \mchip.design.owner.fsm.currentPlayer  = \mchip.design.owner.fsm.currState ;
	assign \mchip.design.owner.fsm.nextState  = \mchip.design.inputSwitchPlayerSync ;
	assign \mchip.design.owner.fsm.reset  = io_in[13];
	assign \mchip.design.owner.fsm.switchTurn  = \mchip.design.inputSwitchPlayerSync ;
	assign \mchip.design.owner.move  = 7'h00;
	assign \mchip.design.owner.newGame  = \mchip.design.inputNewGameSync ;
	assign \mchip.design.owner.player_1_confirm  = \mchip.design.currStateConfirm [1];
	assign \mchip.design.owner.player_1_input  = \mchip.design.inputMovesSync ;
	assign \mchip.design.owner.reset  = io_in[13];
	assign \mchip.design.owner.switchTurn  = \mchip.design.inputSwitchPlayerSync ;
	assign \mchip.design.pve.bot_confirm  = \mchip.design.pve.fsm.currState [2];
	assign \mchip.design.pve.bot_turn  = \mchip.design.inputSwitchPlayerSync ;
	assign \mchip.design.pve.clock  = io_in[12];
	assign \mchip.design.pve.fsm.bot_confirm  = \mchip.design.pve.fsm.currState [2];
	assign \mchip.design.pve.fsm.bot_turn  = \mchip.design.inputSwitchPlayerSync ;
	assign \mchip.design.pve.fsm.clock  = io_in[12];
	assign \mchip.design.pve.fsm.reset  = io_in[13];
	assign \mchip.design.pve.fsm.selectedMove  = 7'h00;
	assign \mchip.design.pve.fsm.timeOutDelay  = 23'h5f5e10;
	assign \mchip.design.pve.fsm.timeOutEn  = \mchip.design.pve.fsm.currState [1];
	assign \mchip.design.pve.rand0.clock  = io_in[12];
	assign \mchip.design.pve.rand0.inputFF [3:1] = \mchip.design.pve.rand0.outputFF [2:0];
	assign \mchip.design.pve.rand0.randomOut  = \mchip.design.pve.rand0.outputFF [3];
	assign \mchip.design.pve.rand0.reset  = io_in[13];
	assign \mchip.design.pve.rand1.clock  = io_in[12];
	assign \mchip.design.pve.rand1.inputFF [3:1] = \mchip.design.pve.rand1.outputFF [2:0];
	assign \mchip.design.pve.rand1.randomOut  = \mchip.design.pve.rand1.outputFF [3];
	assign \mchip.design.pve.rand1.reset  = io_in[13];
	assign \mchip.design.pve.rand2.clock  = io_in[12];
	assign \mchip.design.pve.rand2.inputFF [3:1] = \mchip.design.pve.rand2.outputFF [2:0];
	assign \mchip.design.pve.rand2.randomOut  = \mchip.design.pve.rand2.outputFF [3];
	assign \mchip.design.pve.rand2.reset  = io_in[13];
	assign \mchip.design.pve.rand3.clock  = io_in[12];
	assign \mchip.design.pve.rand3.inputFF [3:1] = \mchip.design.pve.rand3.outputFF [2:0];
	assign \mchip.design.pve.rand3.randomOut  = \mchip.design.pve.rand3.outputFF [3];
	assign \mchip.design.pve.rand3.reset  = io_in[13];
	assign \mchip.design.pve.rand4.clock  = io_in[12];
	assign \mchip.design.pve.rand4.inputFF [3:1] = \mchip.design.pve.rand4.outputFF [2:0];
	assign \mchip.design.pve.rand4.randomOut  = \mchip.design.pve.rand4.outputFF [3];
	assign \mchip.design.pve.rand4.reset  = io_in[13];
	assign \mchip.design.pve.rand5.clock  = io_in[12];
	assign \mchip.design.pve.rand5.inputFF [3:1] = \mchip.design.pve.rand5.outputFF [2:0];
	assign \mchip.design.pve.rand5.randomOut  = \mchip.design.pve.rand5.outputFF [3];
	assign \mchip.design.pve.rand5.reset  = io_in[13];
	assign \mchip.design.pve.rand6.clock  = io_in[12];
	assign \mchip.design.pve.rand6.inputFF [3:1] = \mchip.design.pve.rand6.outputFF [2:0];
	assign \mchip.design.pve.rand6.randomOut  = \mchip.design.pve.rand6.outputFF [3];
	assign \mchip.design.pve.rand6.reset  = io_in[13];
	assign \mchip.design.pve.random  = {\mchip.design.pve.rand6.outputFF [3], \mchip.design.pve.rand5.outputFF [3], \mchip.design.pve.rand4.outputFF [3], \mchip.design.pve.rand3.outputFF [3], \mchip.design.pve.rand2.outputFF [3], \mchip.design.pve.rand1.outputFF [3], \mchip.design.pve.rand0.outputFF [3]};
	assign \mchip.design.pve.reset  = io_in[13];
	assign \mchip.design.pve.tokens  = \mchip.design.owner.tokens ;
	assign \mchip.design.reset  = io_in[13];
	assign \mchip.design.rowFromVGA  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.rowToModule  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.col  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_0_H_0.high  = 10'h054;
	assign \mchip.design.token.level_0_H_0.low  = 10'h02d;
	assign \mchip.design.token.level_0_H_0.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_0_H_14.high  = 10'h054;
	assign \mchip.design.token.level_0_H_14.low  = 10'h02d;
	assign \mchip.design.token.level_0_H_14.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_0_H_21.high  = 10'h054;
	assign \mchip.design.token.level_0_H_21.low  = 10'h02d;
	assign \mchip.design.token.level_0_H_21.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_0_H_28.high  = 10'h054;
	assign \mchip.design.token.level_0_H_28.low  = 10'h02d;
	assign \mchip.design.token.level_0_H_28.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_0_H_35.high  = 10'h054;
	assign \mchip.design.token.level_0_H_35.low  = 10'h02d;
	assign \mchip.design.token.level_0_H_35.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_0_H_7.high  = 10'h054;
	assign \mchip.design.token.level_0_H_7.low  = 10'h02d;
	assign \mchip.design.token.level_0_H_7.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_0_V_0.high  = 9'h04a;
	assign \mchip.design.token.level_0_V_0.low  = 9'h01e;
	assign \mchip.design.token.level_0_V_0.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_0_V_1.high  = 9'h04a;
	assign \mchip.design.token.level_0_V_1.low  = 9'h01e;
	assign \mchip.design.token.level_0_V_1.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_0_V_2.high  = 9'h04a;
	assign \mchip.design.token.level_0_V_2.low  = 9'h01e;
	assign \mchip.design.token.level_0_V_2.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_0_V_3.high  = 9'h04a;
	assign \mchip.design.token.level_0_V_3.low  = 9'h01e;
	assign \mchip.design.token.level_0_V_3.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_0_V_4.high  = 9'h04a;
	assign \mchip.design.token.level_0_V_4.low  = 9'h01e;
	assign \mchip.design.token.level_0_V_4.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_0_V_5.high  = 9'h04a;
	assign \mchip.design.token.level_0_V_5.low  = 9'h01e;
	assign \mchip.design.token.level_0_V_5.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_0_V_6.high  = 9'h04a;
	assign \mchip.design.token.level_0_V_6.low  = 9'h01e;
	assign \mchip.design.token.level_0_V_6.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_1_H_1.high  = 10'h0a9;
	assign \mchip.design.token.level_1_H_1.low  = 10'h082;
	assign \mchip.design.token.level_1_H_1.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_1_H_15.high  = 10'h0a9;
	assign \mchip.design.token.level_1_H_15.low  = 10'h082;
	assign \mchip.design.token.level_1_H_15.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_1_H_22.high  = 10'h0a9;
	assign \mchip.design.token.level_1_H_22.low  = 10'h082;
	assign \mchip.design.token.level_1_H_22.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_1_H_29.high  = 10'h0a9;
	assign \mchip.design.token.level_1_H_29.low  = 10'h082;
	assign \mchip.design.token.level_1_H_29.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_1_H_36.high  = 10'h0a9;
	assign \mchip.design.token.level_1_H_36.low  = 10'h082;
	assign \mchip.design.token.level_1_H_36.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_1_H_8.high  = 10'h0a9;
	assign \mchip.design.token.level_1_H_8.low  = 10'h082;
	assign \mchip.design.token.level_1_H_8.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_1_V_10.high  = 9'h095;
	assign \mchip.design.token.level_1_V_10.low  = 9'h069;
	assign \mchip.design.token.level_1_V_10.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_1_V_11.high  = 9'h095;
	assign \mchip.design.token.level_1_V_11.low  = 9'h069;
	assign \mchip.design.token.level_1_V_11.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_1_V_12.high  = 9'h095;
	assign \mchip.design.token.level_1_V_12.low  = 9'h069;
	assign \mchip.design.token.level_1_V_12.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_1_V_13.high  = 9'h095;
	assign \mchip.design.token.level_1_V_13.low  = 9'h069;
	assign \mchip.design.token.level_1_V_13.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_1_V_7.high  = 9'h095;
	assign \mchip.design.token.level_1_V_7.low  = 9'h069;
	assign \mchip.design.token.level_1_V_7.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_1_V_8.high  = 9'h095;
	assign \mchip.design.token.level_1_V_8.low  = 9'h069;
	assign \mchip.design.token.level_1_V_8.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_1_V_9.high  = 9'h095;
	assign \mchip.design.token.level_1_V_9.low  = 9'h069;
	assign \mchip.design.token.level_1_V_9.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_2_H_16.high  = 10'h0fe;
	assign \mchip.design.token.level_2_H_16.low  = 10'h0d7;
	assign \mchip.design.token.level_2_H_16.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_2_H_2.high  = 10'h0fe;
	assign \mchip.design.token.level_2_H_2.low  = 10'h0d7;
	assign \mchip.design.token.level_2_H_2.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_2_H_23.high  = 10'h0fe;
	assign \mchip.design.token.level_2_H_23.low  = 10'h0d7;
	assign \mchip.design.token.level_2_H_23.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_2_H_30.high  = 10'h0fe;
	assign \mchip.design.token.level_2_H_30.low  = 10'h0d7;
	assign \mchip.design.token.level_2_H_30.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_2_H_37.high  = 10'h0fe;
	assign \mchip.design.token.level_2_H_37.low  = 10'h0d7;
	assign \mchip.design.token.level_2_H_37.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_2_H_9.high  = 10'h0fe;
	assign \mchip.design.token.level_2_H_9.low  = 10'h0d7;
	assign \mchip.design.token.level_2_H_9.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_2_V_14.high  = 9'h0e0;
	assign \mchip.design.token.level_2_V_14.low  = 9'h0b4;
	assign \mchip.design.token.level_2_V_14.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_2_V_15.high  = 9'h0e0;
	assign \mchip.design.token.level_2_V_15.low  = 9'h0b4;
	assign \mchip.design.token.level_2_V_15.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_2_V_16.high  = 9'h0e0;
	assign \mchip.design.token.level_2_V_16.low  = 9'h0b4;
	assign \mchip.design.token.level_2_V_16.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_2_V_17.high  = 9'h0e0;
	assign \mchip.design.token.level_2_V_17.low  = 9'h0b4;
	assign \mchip.design.token.level_2_V_17.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_2_V_18.high  = 9'h0e0;
	assign \mchip.design.token.level_2_V_18.low  = 9'h0b4;
	assign \mchip.design.token.level_2_V_18.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_2_V_19.high  = 9'h0e0;
	assign \mchip.design.token.level_2_V_19.low  = 9'h0b4;
	assign \mchip.design.token.level_2_V_19.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_2_V_20.high  = 9'h0e0;
	assign \mchip.design.token.level_2_V_20.low  = 9'h0b4;
	assign \mchip.design.token.level_2_V_20.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_3_H_10.high  = 10'h153;
	assign \mchip.design.token.level_3_H_10.low  = 10'h12c;
	assign \mchip.design.token.level_3_H_10.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_3_H_17.high  = 10'h153;
	assign \mchip.design.token.level_3_H_17.low  = 10'h12c;
	assign \mchip.design.token.level_3_H_17.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_3_H_24.high  = 10'h153;
	assign \mchip.design.token.level_3_H_24.low  = 10'h12c;
	assign \mchip.design.token.level_3_H_24.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_3_H_3.high  = 10'h153;
	assign \mchip.design.token.level_3_H_3.low  = 10'h12c;
	assign \mchip.design.token.level_3_H_3.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_3_H_31.high  = 10'h153;
	assign \mchip.design.token.level_3_H_31.low  = 10'h12c;
	assign \mchip.design.token.level_3_H_31.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_3_H_38.high  = 10'h153;
	assign \mchip.design.token.level_3_H_38.low  = 10'h12c;
	assign \mchip.design.token.level_3_H_38.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_3_V_21.high  = 9'h12b;
	assign \mchip.design.token.level_3_V_21.low  = 9'h0ff;
	assign \mchip.design.token.level_3_V_21.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_3_V_22.high  = 9'h12b;
	assign \mchip.design.token.level_3_V_22.low  = 9'h0ff;
	assign \mchip.design.token.level_3_V_22.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_3_V_23.high  = 9'h12b;
	assign \mchip.design.token.level_3_V_23.low  = 9'h0ff;
	assign \mchip.design.token.level_3_V_23.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_3_V_24.high  = 9'h12b;
	assign \mchip.design.token.level_3_V_24.low  = 9'h0ff;
	assign \mchip.design.token.level_3_V_24.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_3_V_25.high  = 9'h12b;
	assign \mchip.design.token.level_3_V_25.low  = 9'h0ff;
	assign \mchip.design.token.level_3_V_25.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_3_V_26.high  = 9'h12b;
	assign \mchip.design.token.level_3_V_26.low  = 9'h0ff;
	assign \mchip.design.token.level_3_V_26.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_3_V_27.high  = 9'h12b;
	assign \mchip.design.token.level_3_V_27.low  = 9'h0ff;
	assign \mchip.design.token.level_3_V_27.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_4_H_11.high  = 10'h1a8;
	assign \mchip.design.token.level_4_H_11.low  = 10'h181;
	assign \mchip.design.token.level_4_H_11.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_4_H_18.high  = 10'h1a8;
	assign \mchip.design.token.level_4_H_18.low  = 10'h181;
	assign \mchip.design.token.level_4_H_18.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_4_H_25.high  = 10'h1a8;
	assign \mchip.design.token.level_4_H_25.low  = 10'h181;
	assign \mchip.design.token.level_4_H_25.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_4_H_32.high  = 10'h1a8;
	assign \mchip.design.token.level_4_H_32.low  = 10'h181;
	assign \mchip.design.token.level_4_H_32.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_4_H_39.high  = 10'h1a8;
	assign \mchip.design.token.level_4_H_39.low  = 10'h181;
	assign \mchip.design.token.level_4_H_39.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_4_H_4.high  = 10'h1a8;
	assign \mchip.design.token.level_4_H_4.low  = 10'h181;
	assign \mchip.design.token.level_4_H_4.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_4_V_28.high  = 9'h176;
	assign \mchip.design.token.level_4_V_28.low  = 9'h14a;
	assign \mchip.design.token.level_4_V_28.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_4_V_29.high  = 9'h176;
	assign \mchip.design.token.level_4_V_29.low  = 9'h14a;
	assign \mchip.design.token.level_4_V_29.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_4_V_30.high  = 9'h176;
	assign \mchip.design.token.level_4_V_30.low  = 9'h14a;
	assign \mchip.design.token.level_4_V_30.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_4_V_31.high  = 9'h176;
	assign \mchip.design.token.level_4_V_31.low  = 9'h14a;
	assign \mchip.design.token.level_4_V_31.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_4_V_32.high  = 9'h176;
	assign \mchip.design.token.level_4_V_32.low  = 9'h14a;
	assign \mchip.design.token.level_4_V_32.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_4_V_33.high  = 9'h176;
	assign \mchip.design.token.level_4_V_33.low  = 9'h14a;
	assign \mchip.design.token.level_4_V_33.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_4_V_34.high  = 9'h176;
	assign \mchip.design.token.level_4_V_34.low  = 9'h14a;
	assign \mchip.design.token.level_4_V_34.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_5_H_12.high  = 10'h1fd;
	assign \mchip.design.token.level_5_H_12.low  = 10'h1d6;
	assign \mchip.design.token.level_5_H_12.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_5_H_19.high  = 10'h1fd;
	assign \mchip.design.token.level_5_H_19.low  = 10'h1d6;
	assign \mchip.design.token.level_5_H_19.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_5_H_26.high  = 10'h1fd;
	assign \mchip.design.token.level_5_H_26.low  = 10'h1d6;
	assign \mchip.design.token.level_5_H_26.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_5_H_33.high  = 10'h1fd;
	assign \mchip.design.token.level_5_H_33.low  = 10'h1d6;
	assign \mchip.design.token.level_5_H_33.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_5_H_40.high  = 10'h1fd;
	assign \mchip.design.token.level_5_H_40.low  = 10'h1d6;
	assign \mchip.design.token.level_5_H_40.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_5_H_5.high  = 10'h1fd;
	assign \mchip.design.token.level_5_H_5.low  = 10'h1d6;
	assign \mchip.design.token.level_5_H_5.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_5_V_35.high  = 9'h1c1;
	assign \mchip.design.token.level_5_V_35.low  = 9'h195;
	assign \mchip.design.token.level_5_V_35.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_5_V_36.high  = 9'h1c1;
	assign \mchip.design.token.level_5_V_36.low  = 9'h195;
	assign \mchip.design.token.level_5_V_36.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_5_V_37.high  = 9'h1c1;
	assign \mchip.design.token.level_5_V_37.low  = 9'h195;
	assign \mchip.design.token.level_5_V_37.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_5_V_38.high  = 9'h1c1;
	assign \mchip.design.token.level_5_V_38.low  = 9'h195;
	assign \mchip.design.token.level_5_V_38.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_5_V_39.high  = 9'h1c1;
	assign \mchip.design.token.level_5_V_39.low  = 9'h195;
	assign \mchip.design.token.level_5_V_39.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_5_V_40.high  = 9'h1c1;
	assign \mchip.design.token.level_5_V_40.low  = 9'h195;
	assign \mchip.design.token.level_5_V_40.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_5_V_41.high  = 9'h1c1;
	assign \mchip.design.token.level_5_V_41.low  = 9'h195;
	assign \mchip.design.token.level_5_V_41.val  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.token.level_6_H_13.high  = 10'h252;
	assign \mchip.design.token.level_6_H_13.low  = 10'h22b;
	assign \mchip.design.token.level_6_H_13.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_6_H_20.high  = 10'h252;
	assign \mchip.design.token.level_6_H_20.low  = 10'h22b;
	assign \mchip.design.token.level_6_H_20.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_6_H_27.high  = 10'h252;
	assign \mchip.design.token.level_6_H_27.low  = 10'h22b;
	assign \mchip.design.token.level_6_H_27.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_6_H_34.high  = 10'h252;
	assign \mchip.design.token.level_6_H_34.low  = 10'h22b;
	assign \mchip.design.token.level_6_H_34.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_6_H_41.high  = 10'h252;
	assign \mchip.design.token.level_6_H_41.low  = 10'h22b;
	assign \mchip.design.token.level_6_H_41.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.level_6_H_6.high  = 10'h252;
	assign \mchip.design.token.level_6_H_6.low  = 10'h22b;
	assign \mchip.design.token.level_6_H_6.val  = \mchip.design.vga.h_idx ;
	assign \mchip.design.token.row  = \mchip.design.vga.v_idx [8:0];
	assign \mchip.design.tokens  = \mchip.design.owner.tokens ;
	assign \mchip.design.vga.clk  = io_in[12];
	assign \mchip.design.vga.rst  = io_in[13];
	assign \mchip.design.vga.valid  = \mchip.design.blank ;
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {2'h0, \mchip.design.board.is_board , \mchip.design.board.is_board , io_out[7], io_out[7], io_out[5], io_out[5], 1'h0, \mchip.design.blank , \mchip.design.vga.hsync , \mchip.design.vga.vsync };
	assign \mchip.reset  = io_in[13];
endmodule
module d11_zhexic_i2cdriver (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	reg _027_;
	reg _028_;
	reg _029_;
	reg _030_;
	reg _031_;
	reg _032_;
	reg _033_;
	reg _034_;
	reg _035_;
	reg _036_;
	reg _037_;
	reg _038_;
	reg _039_;
	reg _040_;
	reg _041_;
	reg _042_;
	reg _043_;
	reg _044_;
	reg _045_;
	reg _046_;
	reg _047_;
	reg _048_;
	reg _049_;
	reg _050_;
	reg _051_;
	reg _052_;
	reg _053_;
	reg _054_;
	reg _055_;
	reg _056_;
	reg _057_;
	reg _058_;
	reg _059_;
	reg _060_;
	reg _061_;
	reg _062_;
	reg _063_;
	reg _064_;
	reg _065_;
	reg _066_;
	reg _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire _098_;
	wire _099_;
	wire _100_;
	wire _101_;
	wire _102_;
	wire _103_;
	wire _104_;
	wire _105_;
	wire _106_;
	wire _107_;
	wire _108_;
	wire _109_;
	wire _110_;
	wire _111_;
	wire _112_;
	wire _113_;
	wire _114_;
	wire _115_;
	wire _116_;
	wire _117_;
	wire _118_;
	wire _119_;
	wire _120_;
	wire _121_;
	wire _122_;
	wire _123_;
	wire _124_;
	wire _125_;
	wire _126_;
	wire _127_;
	wire _128_;
	wire _129_;
	wire _130_;
	wire _131_;
	wire _132_;
	wire _133_;
	wire _134_;
	wire _135_;
	wire _136_;
	wire _137_;
	wire _138_;
	wire _139_;
	wire _140_;
	wire _141_;
	wire _142_;
	wire _143_;
	wire _144_;
	wire _145_;
	wire _146_;
	wire _147_;
	wire _148_;
	wire _149_;
	wire _150_;
	wire _151_;
	wire _152_;
	wire _153_;
	wire _154_;
	wire _155_;
	wire _156_;
	wire _157_;
	wire _158_;
	wire _159_;
	wire _160_;
	wire _161_;
	wire _162_;
	wire _163_;
	wire _164_;
	wire _165_;
	wire _166_;
	wire _167_;
	wire _168_;
	wire _169_;
	wire _170_;
	wire _171_;
	wire _172_;
	wire _173_;
	wire _174_;
	wire _175_;
	wire _176_;
	wire _177_;
	wire _178_;
	wire _179_;
	wire _180_;
	wire _181_;
	wire _182_;
	wire _183_;
	wire _184_;
	wire _185_;
	wire _186_;
	wire _187_;
	wire _188_;
	wire _189_;
	wire _190_;
	wire _191_;
	wire _192_;
	wire _193_;
	wire _194_;
	wire _195_;
	wire _196_;
	wire _197_;
	wire _198_;
	wire _199_;
	wire _200_;
	wire _201_;
	wire _202_;
	wire _203_;
	wire _204_;
	wire _205_;
	wire _206_;
	wire _207_;
	wire _208_;
	wire _209_;
	wire _210_;
	wire _211_;
	wire _212_;
	wire _213_;
	wire _214_;
	wire _215_;
	wire _216_;
	wire _217_;
	wire _218_;
	wire _219_;
	wire _220_;
	wire _221_;
	wire _222_;
	wire _223_;
	wire _224_;
	wire _225_;
	wire _226_;
	wire _227_;
	wire _228_;
	wire _229_;
	wire _230_;
	wire _231_;
	wire _232_;
	wire _233_;
	wire _234_;
	wire _235_;
	wire _236_;
	wire _237_;
	wire _238_;
	wire _239_;
	wire _240_;
	wire _241_;
	wire _242_;
	wire _243_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire \mchip.slv.SCL ;
	wire \mchip.slv.SDA_in ;
	wire \mchip.slv.SDA_out ;
	wire \mchip.slv.clock ;
	wire [7:0] \mchip.slv.data_in ;
	wire \mchip.slv.data_incoming ;
	wire [7:0] \mchip.slv.data_out ;
	wire [3:0] \mchip.slv.nextstate ;
	wire \mchip.slv.r1w0 ;
	wire [7:0] \mchip.slv.register_out ;
	wire \mchip.slv.reset ;
	wire \mchip.slv.scl_high ;
	wire \mchip.slv.scl_nextstate ;
	wire \mchip.slv.sda_high ;
	wire \mchip.slv.sda_nextstate ;
	wire [7:0] \mchip.slv.sipo_out ;
	wire \mchip.slv.start_nextstate ;
	wire \mchip.slv.stop_nextstate ;
	wire \mchip.slv.store ;
	wire \mchip.slv.the_piso.clock ;
	wire [7:0] \mchip.slv.the_piso.data_in ;
	wire \mchip.slv.the_piso.reset ;
	wire \mchip.slv.the_reg.clock ;
	wire \mchip.slv.the_reg.enable ;
	wire [7:0] \mchip.slv.the_reg.in ;
	wire [7:0] \mchip.slv.the_reg.out ;
	wire \mchip.slv.the_reg.reset ;
	wire \mchip.slv.the_sipo.clock ;
	wire \mchip.slv.the_sipo.data_in ;
	wire [7:0] \mchip.slv.the_sipo.out ;
	wire \mchip.slv.the_sipo.reset ;
	wire \mchip.slv.wr_down ;
	wire \mchip.slv.wr_up ;
	wire \mchip.slv.writeOK ;
	assign _068_ = ~(_028_ & io_in[13]);
	assign _069_ = _029_ & io_in[13];
	assign _070_ = _068_ & ~_069_;
	assign _071_ = _031_ & io_in[13];
	assign _072_ = _030_ & io_in[13];
	assign _073_ = _071_ | ~_072_;
	assign _074_ = _070_ & ~_073_;
	assign _075_ = _069_ | _068_;
	assign _076_ = ~(_075_ | _073_);
	assign _077_ = ~(_069_ & _068_);
	assign _078_ = ~(_077_ | _073_);
	assign _079_ = _078_ | _076_;
	assign \mchip.slv.wr_down  = _079_ | _074_;
	assign _080_ = io_in[10] & ~\mchip.slv.wr_down ;
	assign _081_ = io_in[13] & ~_062_;
	assign _082_ = _061_ & io_in[13];
	assign _083_ = _082_ | _081_;
	assign _084_ = _060_ & io_in[13];
	assign _085_ = _059_ & io_in[13];
	assign _086_ = _085_ | _084_;
	assign _087_ = _086_ | _083_;
	assign _088_ = io_in[13] & ~_027_;
	assign _089_ = _088_ | io_in[1];
	assign _090_ = _072_ | ~_071_;
	assign _091_ = _070_ & ~_090_;
	assign _092_ = ~(_090_ | _075_);
	assign _093_ = ~(_092_ | _091_);
	assign _094_ = ~(_093_ | _089_);
	assign _095_ = _087_ & ~_089_;
	assign _096_ = ~(_090_ | _077_);
	assign _097_ = _096_ & _095_;
	assign _098_ = _097_ | _094_;
	assign _099_ = _093_ & ~_096_;
	assign _100_ = _098_ & ~_099_;
	assign _001_ = (_087_ ? _100_ : _080_);
	assign _101_ = _066_ & io_in[13];
	assign _102_ = ~(_067_ & io_in[13]);
	assign _103_ = _102_ | _101_;
	assign _104_ = _065_ & io_in[13];
	assign _105_ = _064_ & io_in[13];
	assign _106_ = _105_ | _104_;
	assign _107_ = _106_ | _103_;
	assign _108_ = ~(_088_ & io_in[1]);
	assign _109_ = _108_ | ~_107_;
	assign _110_ = ~(_107_ | _089_);
	assign _111_ = ~(_110_ & _109_);
	assign \mchip.slv.store  = _078_ & ~_111_;
	assign _112_ = _072_ | _071_;
	assign _113_ = _070_ & ~_112_;
	assign _114_ = _089_ | io_in[0];
	assign _115_ = ~(_033_ & io_in[13]);
	assign _116_ = _115_ | _114_;
	assign _117_ = _113_ & ~_116_;
	assign _118_ = _074_ & ~_089_;
	assign _119_ = _118_ | _117_;
	assign _120_ = _071_ | ~_070_;
	assign _121_ = _119_ & ~_120_;
	assign _122_ = ~(_112_ | _075_);
	assign _123_ = ~(_122_ | _078_);
	assign _124_ = _123_ & ~_076_;
	assign _125_ = _123_ | _109_;
	assign _126_ = _076_ & ~_108_;
	assign _127_ = _125_ & ~_126_;
	assign _128_ = _127_ | _124_;
	assign _129_ = _107_ & ~_128_;
	assign _000_ = _129_ | _121_;
	assign _130_ = _063_ & io_in[13];
	assign _131_ = ~_089_;
	assign _132_ = _068_ | ~_069_;
	assign _133_ = _132_ | _112_;
	assign _134_ = _132_ | _073_;
	assign _135_ = ~(_134_ & _133_);
	assign _136_ = _091_ | _074_;
	assign _137_ = (_089_ ? _136_ : _135_);
	assign _138_ = _137_ | \mchip.slv.store ;
	assign _139_ = ~(_136_ | _135_);
	assign _140_ = _139_ & ~_078_;
	assign _141_ = _138_ & ~_140_;
	assign \mchip.slv.SDA_out  = _130_ & ~_141_;
	assign _142_ = ~io_in[0];
	assign _143_ = _142_ & ~_108_;
	assign _144_ = _032_ & io_in[13];
	assign _145_ = _034_ | ~io_in[13];
	assign _146_ = _145_ | _142_;
	assign _147_ = (io_in[1] ? _146_ : _088_);
	assign \mchip.slv.stop_nextstate  = (_144_ ? _147_ : _143_);
	assign _148_ = ~(_145_ & _142_);
	assign _149_ = io_in[1] & ~_148_;
	assign _150_ = io_in[0] & ~_089_;
	assign _151_ = _114_ & ~_150_;
	assign \mchip.slv.start_nextstate  = (_115_ ? _149_ : _151_);
	assign _019_ = _129_ & ~_142_;
	assign _152_ = ~(_035_ & io_in[13]);
	assign \mchip.slv.r1w0  = ~_152_;
	assign _020_ = _129_ & ~_152_;
	assign \mchip.slv.the_sipo.out [1] = _036_ & io_in[13];
	assign _021_ = \mchip.slv.the_sipo.out [1] & _129_;
	assign \mchip.slv.the_sipo.out [2] = _037_ & io_in[13];
	assign _022_ = \mchip.slv.the_sipo.out [2] & _129_;
	assign \mchip.slv.the_sipo.out [3] = _038_ & io_in[13];
	assign _023_ = \mchip.slv.the_sipo.out [3] & _129_;
	assign _153_ = ~(_039_ & io_in[13]);
	assign \mchip.slv.the_sipo.out [4] = ~_153_;
	assign _024_ = _129_ & ~_153_;
	assign \mchip.slv.the_sipo.out [5] = _040_ & io_in[13];
	assign _025_ = \mchip.slv.the_sipo.out [5] & _129_;
	assign \mchip.slv.the_sipo.out [6] = _041_ & io_in[13];
	assign _026_ = \mchip.slv.the_sipo.out [6] & _129_;
	assign _015_ = _129_ & ~_105_;
	assign _154_ = _105_ & _104_;
	assign _155_ = _154_ | ~_106_;
	assign _016_ = _129_ & ~_155_;
	assign _156_ = ~_101_;
	assign _157_ = _154_ ^ _156_;
	assign _017_ = _129_ & ~_157_;
	assign _158_ = _154_ & ~_156_;
	assign _159_ = _158_ ^ _102_;
	assign _018_ = _129_ & ~_159_;
	assign _160_ = _080_ & ~_087_;
	assign _161_ = ~(_058_ & io_in[13]);
	assign _006_ = ~(_161_ | _160_);
	assign _002_ = ~(_160_ | _085_);
	assign _003_ = _085_ ^ _084_;
	assign _162_ = ~_082_;
	assign _163_ = _085_ & _084_;
	assign _164_ = _163_ ^ _162_;
	assign _004_ = ~(_164_ | _160_);
	assign _165_ = _163_ & ~_162_;
	assign _166_ = _165_ ^ _081_;
	assign _005_ = ~(_166_ | _160_);
	assign _007_ = _160_ & io_in[2];
	assign _167_ = _051_ & io_in[13];
	assign _008_ = (_160_ ? io_in[3] : _167_);
	assign _168_ = _052_ & io_in[13];
	assign _009_ = (_160_ ? io_in[4] : _168_);
	assign _169_ = _053_ & io_in[13];
	assign _010_ = (_160_ ? io_in[5] : _169_);
	assign _170_ = _054_ & io_in[13];
	assign _011_ = (_160_ ? io_in[6] : _170_);
	assign _171_ = _055_ & io_in[13];
	assign _012_ = (_160_ ? io_in[7] : _171_);
	assign _172_ = _056_ & io_in[13];
	assign _013_ = (_160_ ? io_in[8] : _172_);
	assign _173_ = _057_ & io_in[13];
	assign _014_ = (_160_ ? io_in[9] : _173_);
	assign _174_ = ~_096_;
	assign _175_ = _089_ | _087_;
	assign _176_ = _175_ & ~_174_;
	assign _177_ = _176_ | _094_;
	assign \mchip.slv.wr_up  = _177_ & ~_099_;
	assign _178_ = ~(_042_ & io_in[13]);
	assign \mchip.slv.the_sipo.out [7] = ~_178_;
	assign _179_ = ~_109_;
	assign _180_ = \mchip.slv.the_sipo.out [1] & ~\mchip.slv.the_sipo.out [2];
	assign _181_ = _153_ | \mchip.slv.the_sipo.out [3];
	assign _182_ = _180_ & ~_181_;
	assign _183_ = \mchip.slv.the_sipo.out [6] | \mchip.slv.the_sipo.out [5];
	assign _184_ = _183_ | _178_;
	assign _185_ = _182_ & ~_184_;
	assign _186_ = ~(_185_ | _107_);
	assign _187_ = _186_ & ~_179_;
	assign _188_ = _122_ & ~_187_;
	assign _189_ = _188_ | _117_;
	assign _190_ = _089_ & ~_133_;
	assign _191_ = _190_ | _189_;
	assign _192_ = _108_ & _076_;
	assign _193_ = _192_ | _118_;
	assign _194_ = _089_ & ~_134_;
	assign _195_ = _194_ | _193_;
	assign _196_ = (_089_ ? _092_ : _091_);
	assign _197_ = _096_ & ~_175_;
	assign _198_ = io_in[0] & ~_108_;
	assign _199_ = ~(_132_ | _090_);
	assign _200_ = _199_ & ~_198_;
	assign _201_ = _200_ | _197_;
	assign _202_ = _201_ | _196_;
	assign _203_ = _202_ | _195_;
	assign _204_ = _203_ | _191_;
	assign _205_ = ~(_072_ & _071_);
	assign \mchip.slv.nextstate [0] = _205_ & _204_;
	assign _206_ = _198_ | _143_;
	assign _207_ = _199_ & ~_206_;
	assign _208_ = _174_ & ~_207_;
	assign _209_ = _092_ & ~_089_;
	assign _210_ = _208_ & ~_209_;
	assign _211_ = _146_ | ~io_in[1];
	assign _212_ = _211_ & ~_110_;
	assign _213_ = _109_ & ~_212_;
	assign _214_ = _078_ & ~_213_;
	assign _215_ = _214_ | _194_;
	assign _216_ = _215_ | _126_;
	assign _217_ = _210_ & ~_216_;
	assign _218_ = _107_ | ~_109_;
	assign _219_ = _122_ & ~_218_;
	assign _220_ = ~(_112_ | _077_);
	assign _221_ = _144_ & ~_211_;
	assign _222_ = _220_ & ~_221_;
	assign _223_ = _222_ | _190_;
	assign _224_ = _223_ | _219_;
	assign _225_ = _217_ & ~_224_;
	assign \mchip.slv.nextstate [1] = _205_ & ~_225_;
	assign _226_ = ~(_076_ | _074_);
	assign _227_ = _211_ | _110_;
	assign _228_ = _109_ & ~_227_;
	assign _229_ = _078_ & ~_228_;
	assign _230_ = _229_ | _194_;
	assign _231_ = _226_ & ~_230_;
	assign _232_ = _107_ | ~_185_;
	assign _233_ = _232_ | _152_;
	assign _234_ = _233_ | _186_;
	assign _235_ = _234_ | _179_;
	assign _236_ = _122_ & ~_235_;
	assign _237_ = _131_ & ~_133_;
	assign _238_ = _237_ | _236_;
	assign _239_ = _231_ & ~_238_;
	assign \mchip.slv.nextstate [2] = _205_ & ~_239_;
	assign _240_ = _200_ | _096_;
	assign _241_ = _093_ & ~_240_;
	assign _242_ = _131_ & ~_134_;
	assign _243_ = _241_ & ~_242_;
	assign \mchip.slv.nextstate [3] = _205_ & ~_243_;
	assign \mchip.slv.writeOK  = ~(_087_ | \mchip.slv.wr_down );
	assign io_out[2] = _043_ & io_in[13];
	assign io_out[3] = _044_ & io_in[13];
	assign io_out[4] = _045_ & io_in[13];
	assign io_out[5] = _046_ & io_in[13];
	assign io_out[6] = _047_ & io_in[13];
	assign io_out[7] = _048_ & io_in[13];
	assign io_out[8] = _049_ & io_in[13];
	assign io_out[9] = _050_ & io_in[13];
	always @(posedge io_in[12])
		if (!io_in[13])
			_027_ <= 1'h1;
		else
			_027_ <= io_in[1];
	always @(posedge io_in[12])
		if (!io_in[13])
			_028_ <= 1'h0;
		else
			_028_ <= \mchip.slv.nextstate [0];
	always @(posedge io_in[12])
		if (!io_in[13])
			_029_ <= 1'h0;
		else
			_029_ <= \mchip.slv.nextstate [1];
	always @(posedge io_in[12])
		if (!io_in[13])
			_030_ <= 1'h0;
		else
			_030_ <= \mchip.slv.nextstate [2];
	always @(posedge io_in[12])
		if (!io_in[13])
			_031_ <= 1'h0;
		else
			_031_ <= \mchip.slv.nextstate [3];
	always @(posedge io_in[12])
		if (!io_in[13])
			_032_ <= 1'h0;
		else
			_032_ <= \mchip.slv.stop_nextstate ;
	always @(posedge io_in[12])
		if (!io_in[13])
			_033_ <= 1'h0;
		else
			_033_ <= \mchip.slv.start_nextstate ;
	always @(posedge io_in[12])
		if (!io_in[13])
			_034_ <= 1'h1;
		else
			_034_ <= io_in[0];
	always @(posedge io_in[12])
		if (!io_in[13])
			_035_ <= 1'h0;
		else if (_000_)
			_035_ <= _019_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_036_ <= 1'h0;
		else if (_000_)
			_036_ <= _020_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_037_ <= 1'h0;
		else if (_000_)
			_037_ <= _021_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_038_ <= 1'h0;
		else if (_000_)
			_038_ <= _022_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_039_ <= 1'h0;
		else if (_000_)
			_039_ <= _023_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_040_ <= 1'h0;
		else if (_000_)
			_040_ <= _024_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_041_ <= 1'h0;
		else if (_000_)
			_041_ <= _025_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_042_ <= 1'h0;
		else if (_000_)
			_042_ <= _026_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_043_ <= 1'h0;
		else if (\mchip.slv.store )
			_043_ <= \mchip.slv.r1w0 ;
	always @(posedge io_in[12])
		if (!io_in[13])
			_044_ <= 1'h0;
		else if (\mchip.slv.store )
			_044_ <= \mchip.slv.the_sipo.out [1];
	always @(posedge io_in[12])
		if (!io_in[13])
			_045_ <= 1'h0;
		else if (\mchip.slv.store )
			_045_ <= \mchip.slv.the_sipo.out [2];
	always @(posedge io_in[12])
		if (!io_in[13])
			_046_ <= 1'h0;
		else if (\mchip.slv.store )
			_046_ <= \mchip.slv.the_sipo.out [3];
	always @(posedge io_in[12])
		if (!io_in[13])
			_047_ <= 1'h0;
		else if (\mchip.slv.store )
			_047_ <= \mchip.slv.the_sipo.out [4];
	always @(posedge io_in[12])
		if (!io_in[13])
			_048_ <= 1'h0;
		else if (\mchip.slv.store )
			_048_ <= \mchip.slv.the_sipo.out [5];
	always @(posedge io_in[12])
		if (!io_in[13])
			_049_ <= 1'h0;
		else if (\mchip.slv.store )
			_049_ <= \mchip.slv.the_sipo.out [6];
	always @(posedge io_in[12])
		if (!io_in[13])
			_050_ <= 1'h0;
		else if (\mchip.slv.store )
			_050_ <= \mchip.slv.the_sipo.out [7];
	always @(posedge io_in[12])
		if (!io_in[13])
			_051_ <= 1'h0;
		else if (_001_)
			_051_ <= _007_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_052_ <= 1'h0;
		else if (_001_)
			_052_ <= _008_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_053_ <= 1'h0;
		else if (_001_)
			_053_ <= _009_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_054_ <= 1'h0;
		else if (_001_)
			_054_ <= _010_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_055_ <= 1'h0;
		else if (_001_)
			_055_ <= _011_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_056_ <= 1'h0;
		else if (_001_)
			_056_ <= _012_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_057_ <= 1'h0;
		else if (_001_)
			_057_ <= _013_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_058_ <= 1'h0;
		else if (_001_)
			_058_ <= _014_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_059_ <= 1'h0;
		else if (_001_)
			_059_ <= _002_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_060_ <= 1'h0;
		else if (_001_)
			_060_ <= _003_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_061_ <= 1'h0;
		else if (_001_)
			_061_ <= _004_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_062_ <= 1'h1;
		else if (_001_)
			_062_ <= _005_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_063_ <= 1'h0;
		else if (_001_)
			_063_ <= _006_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_064_ <= 1'h0;
		else if (_000_)
			_064_ <= _015_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_065_ <= 1'h0;
		else if (_000_)
			_065_ <= _016_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_066_ <= 1'h0;
		else if (_000_)
			_066_ <= _017_;
	always @(posedge io_in[12])
		if (!io_in[13])
			_067_ <= 1'h0;
		else if (_000_)
			_067_ <= _018_;
	assign {io_out[13:10], io_out[1:0]} = {2'h0, \mchip.slv.wr_down , \mchip.slv.writeOK , \mchip.slv.wr_up , \mchip.slv.SDA_out };
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.slv.wr_down , \mchip.slv.writeOK , io_out[9:2], \mchip.slv.wr_up , \mchip.slv.SDA_out };
	assign \mchip.reset  = io_in[13];
	assign \mchip.slv.SCL  = io_in[1];
	assign \mchip.slv.SDA_in  = io_in[0];
	assign \mchip.slv.clock  = io_in[12];
	assign \mchip.slv.data_in  = io_in[9:2];
	assign \mchip.slv.data_incoming  = io_in[10];
	assign \mchip.slv.data_out  = io_out[9:2];
	assign \mchip.slv.register_out  = io_out[9:2];
	assign \mchip.slv.reset  = io_in[13];
	assign \mchip.slv.scl_high  = io_in[1];
	assign \mchip.slv.scl_nextstate  = io_in[1];
	assign \mchip.slv.sda_high  = io_in[0];
	assign \mchip.slv.sda_nextstate  = io_in[0];
	assign \mchip.slv.sipo_out  = {\mchip.slv.the_sipo.out [7:1], \mchip.slv.r1w0 };
	assign \mchip.slv.the_piso.clock  = io_in[12];
	assign \mchip.slv.the_piso.data_in  = io_in[9:2];
	assign \mchip.slv.the_piso.reset  = io_in[13];
	assign \mchip.slv.the_reg.clock  = io_in[12];
	assign \mchip.slv.the_reg.enable  = \mchip.slv.store ;
	assign \mchip.slv.the_reg.in  = {\mchip.slv.the_sipo.out [7:1], \mchip.slv.r1w0 };
	assign \mchip.slv.the_reg.out  = io_out[9:2];
	assign \mchip.slv.the_reg.reset  = io_in[13];
	assign \mchip.slv.the_sipo.clock  = io_in[12];
	assign \mchip.slv.the_sipo.data_in  = io_in[0];
	assign \mchip.slv.the_sipo.out [0] = \mchip.slv.r1w0 ;
	assign \mchip.slv.the_sipo.reset  = io_in[13];
endmodule
module d12_sjg2_tiny_game_of_life (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire _2025_;
	wire _2026_;
	wire _2027_;
	wire _2028_;
	wire _2029_;
	wire _2030_;
	wire _2031_;
	wire _2032_;
	wire _2033_;
	wire _2034_;
	wire _2035_;
	wire _2036_;
	wire _2037_;
	wire _2038_;
	wire _2039_;
	wire _2040_;
	wire _2041_;
	wire _2042_;
	wire _2043_;
	wire _2044_;
	wire _2045_;
	wire _2046_;
	wire _2047_;
	wire _2048_;
	wire _2049_;
	wire _2050_;
	wire _2051_;
	wire _2052_;
	wire _2053_;
	wire _2054_;
	wire _2055_;
	wire _2056_;
	wire _2057_;
	wire _2058_;
	wire _2059_;
	wire _2060_;
	wire _2061_;
	wire _2062_;
	wire _2063_;
	wire _2064_;
	wire _2065_;
	wire _2066_;
	wire _2067_;
	wire _2068_;
	wire _2069_;
	wire _2070_;
	wire _2071_;
	wire _2072_;
	wire _2073_;
	wire _2074_;
	wire _2075_;
	wire _2076_;
	wire _2077_;
	wire _2078_;
	wire _2079_;
	wire _2080_;
	wire _2081_;
	wire _2082_;
	wire _2083_;
	wire _2084_;
	wire _2085_;
	wire _2086_;
	wire _2087_;
	wire _2088_;
	wire _2089_;
	wire _2090_;
	wire _2091_;
	wire _2092_;
	wire _2093_;
	wire _2094_;
	wire _2095_;
	wire _2096_;
	wire _2097_;
	wire _2098_;
	wire _2099_;
	wire _2100_;
	wire _2101_;
	wire _2102_;
	wire _2103_;
	wire _2104_;
	wire _2105_;
	wire _2106_;
	wire _2107_;
	wire _2108_;
	wire _2109_;
	wire _2110_;
	wire _2111_;
	wire _2112_;
	wire _2113_;
	wire _2114_;
	wire [9:0] _2115_;
	wire [9:0] _2116_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [31:0] \mchip.COLS ;
	wire [31:0] \mchip.ROWS ;
	wire [31:0] \mchip.TILE_COLS ;
	wire [31:0] \mchip.TILE_HEIGHT ;
	wire [31:0] \mchip.TILE_ROWS ;
	wire [31:0] \mchip.TILE_WIDTH ;
	wire [2:0] \mchip.blue ;
	wire [639:0] \mchip.bottom ;
	wire [6:0] \mchip.btn ;
	reg \mchip.btn3_sync ;
	reg \mchip.btn3_tmp ;
	reg \mchip.btn4_sync ;
	reg \mchip.btn4_tmp ;
	wire \mchip.clock ;
	reg [2:0] \mchip.focus_col ;
	reg [2:0] \mchip.focus_row ;
	wire \mchip.frame_end ;
	reg \mchip.fsm_state ;
	wire \mchip.gn14 ;
	wire \mchip.gn15 ;
	wire \mchip.gn16 ;
	wire \mchip.gn17 ;
	wire \mchip.gn21 ;
	wire \mchip.gn22 ;
	wire \mchip.gn23 ;
	wire \mchip.gn24 ;
	wire \mchip.gp16 ;
	wire \mchip.gp17 ;
	wire \mchip.gp21 ;
	wire \mchip.gp22 ;
	wire \mchip.gp23 ;
	wire \mchip.gp24 ;
	wire [2:0] \mchip.green ;
	wire [9:0] \mchip.h_idx ;
	wire \mchip.hsync ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire [639:0] \mchip.left ;
	reg \mchip.lock_state ;
	wire [2:0] \mchip.red ;
	wire \mchip.refresh ;
	wire \mchip.reset ;
	wire [639:0] \mchip.right ;
	wire [9:0] \mchip.row_sel[0].col_sel[0].tile.bottom ;
	wire [9:0] \mchip.row_sel[0].col_sel[0].tile.h_idx ;
	wire [9:0] \mchip.row_sel[0].col_sel[0].tile.left ;
	wire [9:0] \mchip.row_sel[0].col_sel[0].tile.right ;
	wire [9:0] \mchip.row_sel[0].col_sel[0].tile.top ;
	wire [9:0] \mchip.row_sel[0].col_sel[0].tile.v_idx ;
	wire \mchip.row_sel[0].col_sel[0].tile_state.clk ;
	wire [2:0] \mchip.row_sel[0].col_sel[0].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[0].col_sel[0].tile_state.focus_row ;
	wire \mchip.row_sel[0].col_sel[0].tile_state.fsm_state ;
	wire \mchip.row_sel[0].col_sel[0].tile_state.lock_state ;
	wire \mchip.row_sel[0].col_sel[0].tile_state.refresh ;
	wire \mchip.row_sel[0].col_sel[0].tile_state.rst ;
	reg \mchip.row_sel[0].col_sel[0].tile_state.state ;
	reg \mchip.row_sel[0].col_sel[0].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[0].col_sel[0].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[0].col_sel[1].tile.bottom ;
	wire [9:0] \mchip.row_sel[0].col_sel[1].tile.h_idx ;
	wire [9:0] \mchip.row_sel[0].col_sel[1].tile.left ;
	wire [9:0] \mchip.row_sel[0].col_sel[1].tile.right ;
	wire [9:0] \mchip.row_sel[0].col_sel[1].tile.top ;
	wire [9:0] \mchip.row_sel[0].col_sel[1].tile.v_idx ;
	wire \mchip.row_sel[0].col_sel[1].tile_state.clk ;
	wire [2:0] \mchip.row_sel[0].col_sel[1].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[0].col_sel[1].tile_state.focus_row ;
	wire \mchip.row_sel[0].col_sel[1].tile_state.fsm_state ;
	wire \mchip.row_sel[0].col_sel[1].tile_state.lock_state ;
	wire [1:0] \mchip.row_sel[0].col_sel[1].tile_state.neighbors_vert ;
	wire \mchip.row_sel[0].col_sel[1].tile_state.refresh ;
	wire \mchip.row_sel[0].col_sel[1].tile_state.rst ;
	reg \mchip.row_sel[0].col_sel[1].tile_state.state ;
	reg \mchip.row_sel[0].col_sel[1].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[0].col_sel[1].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[0].col_sel[2].tile.bottom ;
	wire [9:0] \mchip.row_sel[0].col_sel[2].tile.h_idx ;
	wire [9:0] \mchip.row_sel[0].col_sel[2].tile.left ;
	wire [9:0] \mchip.row_sel[0].col_sel[2].tile.right ;
	wire [9:0] \mchip.row_sel[0].col_sel[2].tile.top ;
	wire [9:0] \mchip.row_sel[0].col_sel[2].tile.v_idx ;
	wire \mchip.row_sel[0].col_sel[2].tile_state.clk ;
	wire [2:0] \mchip.row_sel[0].col_sel[2].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[0].col_sel[2].tile_state.focus_row ;
	wire \mchip.row_sel[0].col_sel[2].tile_state.fsm_state ;
	wire \mchip.row_sel[0].col_sel[2].tile_state.lock_state ;
	wire \mchip.row_sel[0].col_sel[2].tile_state.refresh ;
	wire \mchip.row_sel[0].col_sel[2].tile_state.rst ;
	reg \mchip.row_sel[0].col_sel[2].tile_state.state ;
	reg \mchip.row_sel[0].col_sel[2].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[0].col_sel[2].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[0].col_sel[3].tile.bottom ;
	wire [9:0] \mchip.row_sel[0].col_sel[3].tile.h_idx ;
	wire [9:0] \mchip.row_sel[0].col_sel[3].tile.left ;
	wire [9:0] \mchip.row_sel[0].col_sel[3].tile.right ;
	wire [9:0] \mchip.row_sel[0].col_sel[3].tile.top ;
	wire [9:0] \mchip.row_sel[0].col_sel[3].tile.v_idx ;
	wire \mchip.row_sel[0].col_sel[3].tile_state.clk ;
	wire [2:0] \mchip.row_sel[0].col_sel[3].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[0].col_sel[3].tile_state.focus_row ;
	wire \mchip.row_sel[0].col_sel[3].tile_state.fsm_state ;
	wire \mchip.row_sel[0].col_sel[3].tile_state.lock_state ;
	wire \mchip.row_sel[0].col_sel[3].tile_state.refresh ;
	wire \mchip.row_sel[0].col_sel[3].tile_state.rst ;
	reg \mchip.row_sel[0].col_sel[3].tile_state.state ;
	reg \mchip.row_sel[0].col_sel[3].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[0].col_sel[3].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[0].col_sel[4].tile.bottom ;
	wire [9:0] \mchip.row_sel[0].col_sel[4].tile.h_idx ;
	wire [9:0] \mchip.row_sel[0].col_sel[4].tile.left ;
	wire [9:0] \mchip.row_sel[0].col_sel[4].tile.right ;
	wire [9:0] \mchip.row_sel[0].col_sel[4].tile.top ;
	wire [9:0] \mchip.row_sel[0].col_sel[4].tile.v_idx ;
	wire \mchip.row_sel[0].col_sel[4].tile_state.clk ;
	wire [2:0] \mchip.row_sel[0].col_sel[4].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[0].col_sel[4].tile_state.focus_row ;
	wire \mchip.row_sel[0].col_sel[4].tile_state.fsm_state ;
	wire \mchip.row_sel[0].col_sel[4].tile_state.lock_state ;
	wire \mchip.row_sel[0].col_sel[4].tile_state.refresh ;
	wire \mchip.row_sel[0].col_sel[4].tile_state.rst ;
	reg \mchip.row_sel[0].col_sel[4].tile_state.state ;
	reg \mchip.row_sel[0].col_sel[4].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[0].col_sel[4].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[0].col_sel[5].tile.bottom ;
	wire [9:0] \mchip.row_sel[0].col_sel[5].tile.h_idx ;
	wire [9:0] \mchip.row_sel[0].col_sel[5].tile.left ;
	wire [9:0] \mchip.row_sel[0].col_sel[5].tile.right ;
	wire [9:0] \mchip.row_sel[0].col_sel[5].tile.top ;
	wire [9:0] \mchip.row_sel[0].col_sel[5].tile.v_idx ;
	wire \mchip.row_sel[0].col_sel[5].tile_state.clk ;
	wire [2:0] \mchip.row_sel[0].col_sel[5].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[0].col_sel[5].tile_state.focus_row ;
	wire \mchip.row_sel[0].col_sel[5].tile_state.fsm_state ;
	wire \mchip.row_sel[0].col_sel[5].tile_state.lock_state ;
	wire \mchip.row_sel[0].col_sel[5].tile_state.refresh ;
	wire \mchip.row_sel[0].col_sel[5].tile_state.rst ;
	reg \mchip.row_sel[0].col_sel[5].tile_state.state ;
	reg \mchip.row_sel[0].col_sel[5].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[0].col_sel[5].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[0].col_sel[6].tile.bottom ;
	wire [9:0] \mchip.row_sel[0].col_sel[6].tile.h_idx ;
	wire [9:0] \mchip.row_sel[0].col_sel[6].tile.left ;
	wire [9:0] \mchip.row_sel[0].col_sel[6].tile.right ;
	wire [9:0] \mchip.row_sel[0].col_sel[6].tile.top ;
	wire [9:0] \mchip.row_sel[0].col_sel[6].tile.v_idx ;
	wire \mchip.row_sel[0].col_sel[6].tile_state.clk ;
	wire [2:0] \mchip.row_sel[0].col_sel[6].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[0].col_sel[6].tile_state.focus_row ;
	wire \mchip.row_sel[0].col_sel[6].tile_state.fsm_state ;
	wire \mchip.row_sel[0].col_sel[6].tile_state.lock_state ;
	wire [1:0] \mchip.row_sel[0].col_sel[6].tile_state.neighbors_vert ;
	wire \mchip.row_sel[0].col_sel[6].tile_state.refresh ;
	wire \mchip.row_sel[0].col_sel[6].tile_state.rst ;
	reg \mchip.row_sel[0].col_sel[6].tile_state.state ;
	reg \mchip.row_sel[0].col_sel[6].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[0].col_sel[6].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[0].col_sel[7].tile.bottom ;
	wire [9:0] \mchip.row_sel[0].col_sel[7].tile.h_idx ;
	wire [9:0] \mchip.row_sel[0].col_sel[7].tile.left ;
	wire [9:0] \mchip.row_sel[0].col_sel[7].tile.right ;
	wire [9:0] \mchip.row_sel[0].col_sel[7].tile.top ;
	wire [9:0] \mchip.row_sel[0].col_sel[7].tile.v_idx ;
	wire \mchip.row_sel[0].col_sel[7].tile_state.clk ;
	wire [2:0] \mchip.row_sel[0].col_sel[7].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[0].col_sel[7].tile_state.focus_row ;
	wire \mchip.row_sel[0].col_sel[7].tile_state.fsm_state ;
	wire \mchip.row_sel[0].col_sel[7].tile_state.lock_state ;
	wire \mchip.row_sel[0].col_sel[7].tile_state.refresh ;
	wire \mchip.row_sel[0].col_sel[7].tile_state.rst ;
	reg \mchip.row_sel[0].col_sel[7].tile_state.state ;
	reg \mchip.row_sel[0].col_sel[7].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[0].col_sel[7].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[1].col_sel[0].tile.bottom ;
	wire [9:0] \mchip.row_sel[1].col_sel[0].tile.h_idx ;
	wire [9:0] \mchip.row_sel[1].col_sel[0].tile.left ;
	wire [9:0] \mchip.row_sel[1].col_sel[0].tile.right ;
	wire [9:0] \mchip.row_sel[1].col_sel[0].tile.top ;
	wire [9:0] \mchip.row_sel[1].col_sel[0].tile.v_idx ;
	wire \mchip.row_sel[1].col_sel[0].tile_state.clk ;
	wire [2:0] \mchip.row_sel[1].col_sel[0].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[1].col_sel[0].tile_state.focus_row ;
	wire \mchip.row_sel[1].col_sel[0].tile_state.fsm_state ;
	wire \mchip.row_sel[1].col_sel[0].tile_state.lock_state ;
	wire [1:0] \mchip.row_sel[1].col_sel[0].tile_state.neighbors_hori ;
	wire \mchip.row_sel[1].col_sel[0].tile_state.refresh ;
	wire \mchip.row_sel[1].col_sel[0].tile_state.rst ;
	reg \mchip.row_sel[1].col_sel[0].tile_state.state ;
	reg \mchip.row_sel[1].col_sel[0].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[1].col_sel[0].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[1].col_sel[1].tile.bottom ;
	wire [9:0] \mchip.row_sel[1].col_sel[1].tile.h_idx ;
	wire [9:0] \mchip.row_sel[1].col_sel[1].tile.left ;
	wire [9:0] \mchip.row_sel[1].col_sel[1].tile.right ;
	wire [9:0] \mchip.row_sel[1].col_sel[1].tile.top ;
	wire [9:0] \mchip.row_sel[1].col_sel[1].tile.v_idx ;
	wire \mchip.row_sel[1].col_sel[1].tile_state.clk ;
	wire [2:0] \mchip.row_sel[1].col_sel[1].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[1].col_sel[1].tile_state.focus_row ;
	wire \mchip.row_sel[1].col_sel[1].tile_state.fsm_state ;
	wire \mchip.row_sel[1].col_sel[1].tile_state.lock_state ;
	wire \mchip.row_sel[1].col_sel[1].tile_state.refresh ;
	wire \mchip.row_sel[1].col_sel[1].tile_state.rst ;
	reg \mchip.row_sel[1].col_sel[1].tile_state.state ;
	reg \mchip.row_sel[1].col_sel[1].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[1].col_sel[1].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[1].col_sel[2].tile.bottom ;
	wire [9:0] \mchip.row_sel[1].col_sel[2].tile.h_idx ;
	wire [9:0] \mchip.row_sel[1].col_sel[2].tile.left ;
	wire [9:0] \mchip.row_sel[1].col_sel[2].tile.right ;
	wire [9:0] \mchip.row_sel[1].col_sel[2].tile.top ;
	wire [9:0] \mchip.row_sel[1].col_sel[2].tile.v_idx ;
	wire \mchip.row_sel[1].col_sel[2].tile_state.clk ;
	wire [2:0] \mchip.row_sel[1].col_sel[2].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[1].col_sel[2].tile_state.focus_row ;
	wire \mchip.row_sel[1].col_sel[2].tile_state.fsm_state ;
	wire \mchip.row_sel[1].col_sel[2].tile_state.lock_state ;
	wire \mchip.row_sel[1].col_sel[2].tile_state.refresh ;
	wire \mchip.row_sel[1].col_sel[2].tile_state.rst ;
	reg \mchip.row_sel[1].col_sel[2].tile_state.state ;
	reg \mchip.row_sel[1].col_sel[2].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[1].col_sel[2].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[1].col_sel[3].tile.bottom ;
	wire [9:0] \mchip.row_sel[1].col_sel[3].tile.h_idx ;
	wire [9:0] \mchip.row_sel[1].col_sel[3].tile.left ;
	wire [9:0] \mchip.row_sel[1].col_sel[3].tile.right ;
	wire [9:0] \mchip.row_sel[1].col_sel[3].tile.top ;
	wire [9:0] \mchip.row_sel[1].col_sel[3].tile.v_idx ;
	wire \mchip.row_sel[1].col_sel[3].tile_state.clk ;
	wire [2:0] \mchip.row_sel[1].col_sel[3].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[1].col_sel[3].tile_state.focus_row ;
	wire \mchip.row_sel[1].col_sel[3].tile_state.fsm_state ;
	wire \mchip.row_sel[1].col_sel[3].tile_state.lock_state ;
	wire \mchip.row_sel[1].col_sel[3].tile_state.refresh ;
	wire \mchip.row_sel[1].col_sel[3].tile_state.rst ;
	reg \mchip.row_sel[1].col_sel[3].tile_state.state ;
	reg \mchip.row_sel[1].col_sel[3].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[1].col_sel[3].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[1].col_sel[4].tile.bottom ;
	wire [9:0] \mchip.row_sel[1].col_sel[4].tile.h_idx ;
	wire [9:0] \mchip.row_sel[1].col_sel[4].tile.left ;
	wire [9:0] \mchip.row_sel[1].col_sel[4].tile.right ;
	wire [9:0] \mchip.row_sel[1].col_sel[4].tile.top ;
	wire [9:0] \mchip.row_sel[1].col_sel[4].tile.v_idx ;
	wire \mchip.row_sel[1].col_sel[4].tile_state.clk ;
	wire [2:0] \mchip.row_sel[1].col_sel[4].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[1].col_sel[4].tile_state.focus_row ;
	wire \mchip.row_sel[1].col_sel[4].tile_state.fsm_state ;
	wire \mchip.row_sel[1].col_sel[4].tile_state.lock_state ;
	wire \mchip.row_sel[1].col_sel[4].tile_state.refresh ;
	wire \mchip.row_sel[1].col_sel[4].tile_state.rst ;
	reg \mchip.row_sel[1].col_sel[4].tile_state.state ;
	reg \mchip.row_sel[1].col_sel[4].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[1].col_sel[4].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[1].col_sel[5].tile.bottom ;
	wire [9:0] \mchip.row_sel[1].col_sel[5].tile.h_idx ;
	wire [9:0] \mchip.row_sel[1].col_sel[5].tile.left ;
	wire [9:0] \mchip.row_sel[1].col_sel[5].tile.right ;
	wire [9:0] \mchip.row_sel[1].col_sel[5].tile.top ;
	wire [9:0] \mchip.row_sel[1].col_sel[5].tile.v_idx ;
	wire \mchip.row_sel[1].col_sel[5].tile_state.clk ;
	wire [2:0] \mchip.row_sel[1].col_sel[5].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[1].col_sel[5].tile_state.focus_row ;
	wire \mchip.row_sel[1].col_sel[5].tile_state.fsm_state ;
	wire \mchip.row_sel[1].col_sel[5].tile_state.lock_state ;
	wire \mchip.row_sel[1].col_sel[5].tile_state.refresh ;
	wire \mchip.row_sel[1].col_sel[5].tile_state.rst ;
	reg \mchip.row_sel[1].col_sel[5].tile_state.state ;
	reg \mchip.row_sel[1].col_sel[5].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[1].col_sel[5].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[1].col_sel[6].tile.bottom ;
	wire [9:0] \mchip.row_sel[1].col_sel[6].tile.h_idx ;
	wire [9:0] \mchip.row_sel[1].col_sel[6].tile.left ;
	wire [9:0] \mchip.row_sel[1].col_sel[6].tile.right ;
	wire [9:0] \mchip.row_sel[1].col_sel[6].tile.top ;
	wire [9:0] \mchip.row_sel[1].col_sel[6].tile.v_idx ;
	wire \mchip.row_sel[1].col_sel[6].tile_state.clk ;
	wire [2:0] \mchip.row_sel[1].col_sel[6].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[1].col_sel[6].tile_state.focus_row ;
	wire \mchip.row_sel[1].col_sel[6].tile_state.fsm_state ;
	wire \mchip.row_sel[1].col_sel[6].tile_state.lock_state ;
	wire \mchip.row_sel[1].col_sel[6].tile_state.refresh ;
	wire \mchip.row_sel[1].col_sel[6].tile_state.rst ;
	reg \mchip.row_sel[1].col_sel[6].tile_state.state ;
	reg \mchip.row_sel[1].col_sel[6].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[1].col_sel[6].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[1].col_sel[7].tile.bottom ;
	wire [9:0] \mchip.row_sel[1].col_sel[7].tile.h_idx ;
	wire [9:0] \mchip.row_sel[1].col_sel[7].tile.left ;
	wire [9:0] \mchip.row_sel[1].col_sel[7].tile.right ;
	wire [9:0] \mchip.row_sel[1].col_sel[7].tile.top ;
	wire [9:0] \mchip.row_sel[1].col_sel[7].tile.v_idx ;
	wire \mchip.row_sel[1].col_sel[7].tile_state.clk ;
	wire [2:0] \mchip.row_sel[1].col_sel[7].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[1].col_sel[7].tile_state.focus_row ;
	wire \mchip.row_sel[1].col_sel[7].tile_state.fsm_state ;
	wire \mchip.row_sel[1].col_sel[7].tile_state.lock_state ;
	wire [1:0] \mchip.row_sel[1].col_sel[7].tile_state.neighbors_hori ;
	wire \mchip.row_sel[1].col_sel[7].tile_state.refresh ;
	wire \mchip.row_sel[1].col_sel[7].tile_state.rst ;
	reg \mchip.row_sel[1].col_sel[7].tile_state.state ;
	reg \mchip.row_sel[1].col_sel[7].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[1].col_sel[7].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[2].col_sel[0].tile.bottom ;
	wire [9:0] \mchip.row_sel[2].col_sel[0].tile.h_idx ;
	wire [9:0] \mchip.row_sel[2].col_sel[0].tile.left ;
	wire [9:0] \mchip.row_sel[2].col_sel[0].tile.right ;
	wire [9:0] \mchip.row_sel[2].col_sel[0].tile.top ;
	wire [9:0] \mchip.row_sel[2].col_sel[0].tile.v_idx ;
	wire \mchip.row_sel[2].col_sel[0].tile_state.clk ;
	wire [2:0] \mchip.row_sel[2].col_sel[0].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[2].col_sel[0].tile_state.focus_row ;
	wire \mchip.row_sel[2].col_sel[0].tile_state.fsm_state ;
	wire \mchip.row_sel[2].col_sel[0].tile_state.lock_state ;
	wire \mchip.row_sel[2].col_sel[0].tile_state.refresh ;
	wire \mchip.row_sel[2].col_sel[0].tile_state.rst ;
	reg \mchip.row_sel[2].col_sel[0].tile_state.state ;
	reg \mchip.row_sel[2].col_sel[0].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[2].col_sel[0].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[2].col_sel[1].tile.bottom ;
	wire [9:0] \mchip.row_sel[2].col_sel[1].tile.h_idx ;
	wire [9:0] \mchip.row_sel[2].col_sel[1].tile.left ;
	wire [9:0] \mchip.row_sel[2].col_sel[1].tile.right ;
	wire [9:0] \mchip.row_sel[2].col_sel[1].tile.top ;
	wire [9:0] \mchip.row_sel[2].col_sel[1].tile.v_idx ;
	wire \mchip.row_sel[2].col_sel[1].tile_state.clk ;
	wire [2:0] \mchip.row_sel[2].col_sel[1].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[2].col_sel[1].tile_state.focus_row ;
	wire \mchip.row_sel[2].col_sel[1].tile_state.fsm_state ;
	wire \mchip.row_sel[2].col_sel[1].tile_state.lock_state ;
	wire \mchip.row_sel[2].col_sel[1].tile_state.refresh ;
	wire \mchip.row_sel[2].col_sel[1].tile_state.rst ;
	reg \mchip.row_sel[2].col_sel[1].tile_state.state ;
	reg \mchip.row_sel[2].col_sel[1].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[2].col_sel[1].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[2].col_sel[2].tile.bottom ;
	wire [9:0] \mchip.row_sel[2].col_sel[2].tile.h_idx ;
	wire [9:0] \mchip.row_sel[2].col_sel[2].tile.left ;
	wire [9:0] \mchip.row_sel[2].col_sel[2].tile.right ;
	wire [9:0] \mchip.row_sel[2].col_sel[2].tile.top ;
	wire [9:0] \mchip.row_sel[2].col_sel[2].tile.v_idx ;
	wire \mchip.row_sel[2].col_sel[2].tile_state.clk ;
	wire [2:0] \mchip.row_sel[2].col_sel[2].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[2].col_sel[2].tile_state.focus_row ;
	wire \mchip.row_sel[2].col_sel[2].tile_state.fsm_state ;
	wire \mchip.row_sel[2].col_sel[2].tile_state.lock_state ;
	wire \mchip.row_sel[2].col_sel[2].tile_state.refresh ;
	wire \mchip.row_sel[2].col_sel[2].tile_state.rst ;
	reg \mchip.row_sel[2].col_sel[2].tile_state.state ;
	reg \mchip.row_sel[2].col_sel[2].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[2].col_sel[2].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[2].col_sel[3].tile.bottom ;
	wire [9:0] \mchip.row_sel[2].col_sel[3].tile.h_idx ;
	wire [9:0] \mchip.row_sel[2].col_sel[3].tile.left ;
	wire [9:0] \mchip.row_sel[2].col_sel[3].tile.right ;
	wire [9:0] \mchip.row_sel[2].col_sel[3].tile.top ;
	wire [9:0] \mchip.row_sel[2].col_sel[3].tile.v_idx ;
	wire \mchip.row_sel[2].col_sel[3].tile_state.clk ;
	wire [2:0] \mchip.row_sel[2].col_sel[3].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[2].col_sel[3].tile_state.focus_row ;
	wire \mchip.row_sel[2].col_sel[3].tile_state.fsm_state ;
	wire \mchip.row_sel[2].col_sel[3].tile_state.lock_state ;
	wire \mchip.row_sel[2].col_sel[3].tile_state.refresh ;
	wire \mchip.row_sel[2].col_sel[3].tile_state.rst ;
	reg \mchip.row_sel[2].col_sel[3].tile_state.state ;
	reg \mchip.row_sel[2].col_sel[3].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[2].col_sel[3].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[2].col_sel[4].tile.bottom ;
	wire [9:0] \mchip.row_sel[2].col_sel[4].tile.h_idx ;
	wire [9:0] \mchip.row_sel[2].col_sel[4].tile.left ;
	wire [9:0] \mchip.row_sel[2].col_sel[4].tile.right ;
	wire [9:0] \mchip.row_sel[2].col_sel[4].tile.top ;
	wire [9:0] \mchip.row_sel[2].col_sel[4].tile.v_idx ;
	wire \mchip.row_sel[2].col_sel[4].tile_state.clk ;
	wire [2:0] \mchip.row_sel[2].col_sel[4].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[2].col_sel[4].tile_state.focus_row ;
	wire \mchip.row_sel[2].col_sel[4].tile_state.fsm_state ;
	wire \mchip.row_sel[2].col_sel[4].tile_state.lock_state ;
	wire \mchip.row_sel[2].col_sel[4].tile_state.refresh ;
	wire \mchip.row_sel[2].col_sel[4].tile_state.rst ;
	reg \mchip.row_sel[2].col_sel[4].tile_state.state ;
	reg \mchip.row_sel[2].col_sel[4].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[2].col_sel[4].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[2].col_sel[5].tile.bottom ;
	wire [9:0] \mchip.row_sel[2].col_sel[5].tile.h_idx ;
	wire [9:0] \mchip.row_sel[2].col_sel[5].tile.left ;
	wire [9:0] \mchip.row_sel[2].col_sel[5].tile.right ;
	wire [9:0] \mchip.row_sel[2].col_sel[5].tile.top ;
	wire [9:0] \mchip.row_sel[2].col_sel[5].tile.v_idx ;
	wire \mchip.row_sel[2].col_sel[5].tile_state.clk ;
	wire [2:0] \mchip.row_sel[2].col_sel[5].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[2].col_sel[5].tile_state.focus_row ;
	wire \mchip.row_sel[2].col_sel[5].tile_state.fsm_state ;
	wire \mchip.row_sel[2].col_sel[5].tile_state.lock_state ;
	wire \mchip.row_sel[2].col_sel[5].tile_state.refresh ;
	wire \mchip.row_sel[2].col_sel[5].tile_state.rst ;
	reg \mchip.row_sel[2].col_sel[5].tile_state.state ;
	reg \mchip.row_sel[2].col_sel[5].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[2].col_sel[5].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[2].col_sel[6].tile.bottom ;
	wire [9:0] \mchip.row_sel[2].col_sel[6].tile.h_idx ;
	wire [9:0] \mchip.row_sel[2].col_sel[6].tile.left ;
	wire [9:0] \mchip.row_sel[2].col_sel[6].tile.right ;
	wire [9:0] \mchip.row_sel[2].col_sel[6].tile.top ;
	wire [9:0] \mchip.row_sel[2].col_sel[6].tile.v_idx ;
	wire \mchip.row_sel[2].col_sel[6].tile_state.clk ;
	wire [2:0] \mchip.row_sel[2].col_sel[6].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[2].col_sel[6].tile_state.focus_row ;
	wire \mchip.row_sel[2].col_sel[6].tile_state.fsm_state ;
	wire \mchip.row_sel[2].col_sel[6].tile_state.lock_state ;
	wire \mchip.row_sel[2].col_sel[6].tile_state.refresh ;
	wire \mchip.row_sel[2].col_sel[6].tile_state.rst ;
	reg \mchip.row_sel[2].col_sel[6].tile_state.state ;
	reg \mchip.row_sel[2].col_sel[6].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[2].col_sel[6].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[2].col_sel[7].tile.bottom ;
	wire [9:0] \mchip.row_sel[2].col_sel[7].tile.h_idx ;
	wire [9:0] \mchip.row_sel[2].col_sel[7].tile.left ;
	wire [9:0] \mchip.row_sel[2].col_sel[7].tile.right ;
	wire [9:0] \mchip.row_sel[2].col_sel[7].tile.top ;
	wire [9:0] \mchip.row_sel[2].col_sel[7].tile.v_idx ;
	wire \mchip.row_sel[2].col_sel[7].tile_state.clk ;
	wire [2:0] \mchip.row_sel[2].col_sel[7].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[2].col_sel[7].tile_state.focus_row ;
	wire \mchip.row_sel[2].col_sel[7].tile_state.fsm_state ;
	wire \mchip.row_sel[2].col_sel[7].tile_state.lock_state ;
	wire \mchip.row_sel[2].col_sel[7].tile_state.refresh ;
	wire \mchip.row_sel[2].col_sel[7].tile_state.rst ;
	reg \mchip.row_sel[2].col_sel[7].tile_state.state ;
	reg \mchip.row_sel[2].col_sel[7].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[2].col_sel[7].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[3].col_sel[0].tile.bottom ;
	wire [9:0] \mchip.row_sel[3].col_sel[0].tile.h_idx ;
	wire [9:0] \mchip.row_sel[3].col_sel[0].tile.left ;
	wire [9:0] \mchip.row_sel[3].col_sel[0].tile.right ;
	wire [9:0] \mchip.row_sel[3].col_sel[0].tile.top ;
	wire [9:0] \mchip.row_sel[3].col_sel[0].tile.v_idx ;
	wire \mchip.row_sel[3].col_sel[0].tile_state.clk ;
	wire [2:0] \mchip.row_sel[3].col_sel[0].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[3].col_sel[0].tile_state.focus_row ;
	wire \mchip.row_sel[3].col_sel[0].tile_state.fsm_state ;
	wire \mchip.row_sel[3].col_sel[0].tile_state.lock_state ;
	wire \mchip.row_sel[3].col_sel[0].tile_state.refresh ;
	wire \mchip.row_sel[3].col_sel[0].tile_state.rst ;
	reg \mchip.row_sel[3].col_sel[0].tile_state.state ;
	reg \mchip.row_sel[3].col_sel[0].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[3].col_sel[0].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[3].col_sel[1].tile.bottom ;
	wire [9:0] \mchip.row_sel[3].col_sel[1].tile.h_idx ;
	wire [9:0] \mchip.row_sel[3].col_sel[1].tile.left ;
	wire [9:0] \mchip.row_sel[3].col_sel[1].tile.right ;
	wire [9:0] \mchip.row_sel[3].col_sel[1].tile.top ;
	wire [9:0] \mchip.row_sel[3].col_sel[1].tile.v_idx ;
	wire \mchip.row_sel[3].col_sel[1].tile_state.clk ;
	wire [2:0] \mchip.row_sel[3].col_sel[1].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[3].col_sel[1].tile_state.focus_row ;
	wire \mchip.row_sel[3].col_sel[1].tile_state.fsm_state ;
	wire \mchip.row_sel[3].col_sel[1].tile_state.lock_state ;
	wire \mchip.row_sel[3].col_sel[1].tile_state.refresh ;
	wire \mchip.row_sel[3].col_sel[1].tile_state.rst ;
	reg \mchip.row_sel[3].col_sel[1].tile_state.state ;
	reg \mchip.row_sel[3].col_sel[1].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[3].col_sel[1].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[3].col_sel[2].tile.bottom ;
	wire [9:0] \mchip.row_sel[3].col_sel[2].tile.h_idx ;
	wire [9:0] \mchip.row_sel[3].col_sel[2].tile.left ;
	wire [9:0] \mchip.row_sel[3].col_sel[2].tile.right ;
	wire [9:0] \mchip.row_sel[3].col_sel[2].tile.top ;
	wire [9:0] \mchip.row_sel[3].col_sel[2].tile.v_idx ;
	wire \mchip.row_sel[3].col_sel[2].tile_state.clk ;
	wire [2:0] \mchip.row_sel[3].col_sel[2].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[3].col_sel[2].tile_state.focus_row ;
	wire \mchip.row_sel[3].col_sel[2].tile_state.fsm_state ;
	wire \mchip.row_sel[3].col_sel[2].tile_state.lock_state ;
	wire \mchip.row_sel[3].col_sel[2].tile_state.refresh ;
	wire \mchip.row_sel[3].col_sel[2].tile_state.rst ;
	reg \mchip.row_sel[3].col_sel[2].tile_state.state ;
	reg \mchip.row_sel[3].col_sel[2].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[3].col_sel[2].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[3].col_sel[3].tile.bottom ;
	wire [9:0] \mchip.row_sel[3].col_sel[3].tile.h_idx ;
	wire [9:0] \mchip.row_sel[3].col_sel[3].tile.left ;
	wire [9:0] \mchip.row_sel[3].col_sel[3].tile.right ;
	wire [9:0] \mchip.row_sel[3].col_sel[3].tile.top ;
	wire [9:0] \mchip.row_sel[3].col_sel[3].tile.v_idx ;
	wire \mchip.row_sel[3].col_sel[3].tile_state.clk ;
	wire [2:0] \mchip.row_sel[3].col_sel[3].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[3].col_sel[3].tile_state.focus_row ;
	wire \mchip.row_sel[3].col_sel[3].tile_state.fsm_state ;
	wire \mchip.row_sel[3].col_sel[3].tile_state.lock_state ;
	wire \mchip.row_sel[3].col_sel[3].tile_state.refresh ;
	wire \mchip.row_sel[3].col_sel[3].tile_state.rst ;
	reg \mchip.row_sel[3].col_sel[3].tile_state.state ;
	reg \mchip.row_sel[3].col_sel[3].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[3].col_sel[3].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[3].col_sel[4].tile.bottom ;
	wire [9:0] \mchip.row_sel[3].col_sel[4].tile.h_idx ;
	wire [9:0] \mchip.row_sel[3].col_sel[4].tile.left ;
	wire [9:0] \mchip.row_sel[3].col_sel[4].tile.right ;
	wire [9:0] \mchip.row_sel[3].col_sel[4].tile.top ;
	wire [9:0] \mchip.row_sel[3].col_sel[4].tile.v_idx ;
	wire \mchip.row_sel[3].col_sel[4].tile_state.clk ;
	wire [2:0] \mchip.row_sel[3].col_sel[4].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[3].col_sel[4].tile_state.focus_row ;
	wire \mchip.row_sel[3].col_sel[4].tile_state.fsm_state ;
	wire \mchip.row_sel[3].col_sel[4].tile_state.lock_state ;
	wire \mchip.row_sel[3].col_sel[4].tile_state.refresh ;
	wire \mchip.row_sel[3].col_sel[4].tile_state.rst ;
	reg \mchip.row_sel[3].col_sel[4].tile_state.state ;
	reg \mchip.row_sel[3].col_sel[4].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[3].col_sel[4].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[3].col_sel[5].tile.bottom ;
	wire [9:0] \mchip.row_sel[3].col_sel[5].tile.h_idx ;
	wire [9:0] \mchip.row_sel[3].col_sel[5].tile.left ;
	wire [9:0] \mchip.row_sel[3].col_sel[5].tile.right ;
	wire [9:0] \mchip.row_sel[3].col_sel[5].tile.top ;
	wire [9:0] \mchip.row_sel[3].col_sel[5].tile.v_idx ;
	wire \mchip.row_sel[3].col_sel[5].tile_state.clk ;
	wire [2:0] \mchip.row_sel[3].col_sel[5].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[3].col_sel[5].tile_state.focus_row ;
	wire \mchip.row_sel[3].col_sel[5].tile_state.fsm_state ;
	wire \mchip.row_sel[3].col_sel[5].tile_state.lock_state ;
	wire \mchip.row_sel[3].col_sel[5].tile_state.refresh ;
	wire \mchip.row_sel[3].col_sel[5].tile_state.rst ;
	reg \mchip.row_sel[3].col_sel[5].tile_state.state ;
	reg \mchip.row_sel[3].col_sel[5].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[3].col_sel[5].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[3].col_sel[6].tile.bottom ;
	wire [9:0] \mchip.row_sel[3].col_sel[6].tile.h_idx ;
	wire [9:0] \mchip.row_sel[3].col_sel[6].tile.left ;
	wire [9:0] \mchip.row_sel[3].col_sel[6].tile.right ;
	wire [9:0] \mchip.row_sel[3].col_sel[6].tile.top ;
	wire [9:0] \mchip.row_sel[3].col_sel[6].tile.v_idx ;
	wire \mchip.row_sel[3].col_sel[6].tile_state.clk ;
	wire [2:0] \mchip.row_sel[3].col_sel[6].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[3].col_sel[6].tile_state.focus_row ;
	wire \mchip.row_sel[3].col_sel[6].tile_state.fsm_state ;
	wire \mchip.row_sel[3].col_sel[6].tile_state.lock_state ;
	wire \mchip.row_sel[3].col_sel[6].tile_state.refresh ;
	wire \mchip.row_sel[3].col_sel[6].tile_state.rst ;
	reg \mchip.row_sel[3].col_sel[6].tile_state.state ;
	reg \mchip.row_sel[3].col_sel[6].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[3].col_sel[6].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[3].col_sel[7].tile.bottom ;
	wire [9:0] \mchip.row_sel[3].col_sel[7].tile.h_idx ;
	wire [9:0] \mchip.row_sel[3].col_sel[7].tile.left ;
	wire [9:0] \mchip.row_sel[3].col_sel[7].tile.right ;
	wire [9:0] \mchip.row_sel[3].col_sel[7].tile.top ;
	wire [9:0] \mchip.row_sel[3].col_sel[7].tile.v_idx ;
	wire \mchip.row_sel[3].col_sel[7].tile_state.clk ;
	wire [2:0] \mchip.row_sel[3].col_sel[7].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[3].col_sel[7].tile_state.focus_row ;
	wire \mchip.row_sel[3].col_sel[7].tile_state.fsm_state ;
	wire \mchip.row_sel[3].col_sel[7].tile_state.lock_state ;
	wire \mchip.row_sel[3].col_sel[7].tile_state.refresh ;
	wire \mchip.row_sel[3].col_sel[7].tile_state.rst ;
	reg \mchip.row_sel[3].col_sel[7].tile_state.state ;
	reg \mchip.row_sel[3].col_sel[7].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[3].col_sel[7].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[4].col_sel[0].tile.bottom ;
	wire [9:0] \mchip.row_sel[4].col_sel[0].tile.h_idx ;
	wire [9:0] \mchip.row_sel[4].col_sel[0].tile.left ;
	wire [9:0] \mchip.row_sel[4].col_sel[0].tile.right ;
	wire [9:0] \mchip.row_sel[4].col_sel[0].tile.top ;
	wire [9:0] \mchip.row_sel[4].col_sel[0].tile.v_idx ;
	wire \mchip.row_sel[4].col_sel[0].tile_state.clk ;
	wire [2:0] \mchip.row_sel[4].col_sel[0].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[4].col_sel[0].tile_state.focus_row ;
	wire \mchip.row_sel[4].col_sel[0].tile_state.fsm_state ;
	wire \mchip.row_sel[4].col_sel[0].tile_state.lock_state ;
	wire \mchip.row_sel[4].col_sel[0].tile_state.refresh ;
	wire \mchip.row_sel[4].col_sel[0].tile_state.rst ;
	reg \mchip.row_sel[4].col_sel[0].tile_state.state ;
	reg \mchip.row_sel[4].col_sel[0].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[4].col_sel[0].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[4].col_sel[1].tile.bottom ;
	wire [9:0] \mchip.row_sel[4].col_sel[1].tile.h_idx ;
	wire [9:0] \mchip.row_sel[4].col_sel[1].tile.left ;
	wire [9:0] \mchip.row_sel[4].col_sel[1].tile.right ;
	wire [9:0] \mchip.row_sel[4].col_sel[1].tile.top ;
	wire [9:0] \mchip.row_sel[4].col_sel[1].tile.v_idx ;
	wire \mchip.row_sel[4].col_sel[1].tile_state.clk ;
	wire [2:0] \mchip.row_sel[4].col_sel[1].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[4].col_sel[1].tile_state.focus_row ;
	wire \mchip.row_sel[4].col_sel[1].tile_state.fsm_state ;
	wire \mchip.row_sel[4].col_sel[1].tile_state.lock_state ;
	wire \mchip.row_sel[4].col_sel[1].tile_state.refresh ;
	wire \mchip.row_sel[4].col_sel[1].tile_state.rst ;
	reg \mchip.row_sel[4].col_sel[1].tile_state.state ;
	reg \mchip.row_sel[4].col_sel[1].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[4].col_sel[1].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[4].col_sel[2].tile.bottom ;
	wire [9:0] \mchip.row_sel[4].col_sel[2].tile.h_idx ;
	wire [9:0] \mchip.row_sel[4].col_sel[2].tile.left ;
	wire [9:0] \mchip.row_sel[4].col_sel[2].tile.right ;
	wire [9:0] \mchip.row_sel[4].col_sel[2].tile.top ;
	wire [9:0] \mchip.row_sel[4].col_sel[2].tile.v_idx ;
	wire \mchip.row_sel[4].col_sel[2].tile_state.clk ;
	wire [2:0] \mchip.row_sel[4].col_sel[2].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[4].col_sel[2].tile_state.focus_row ;
	wire \mchip.row_sel[4].col_sel[2].tile_state.fsm_state ;
	wire \mchip.row_sel[4].col_sel[2].tile_state.lock_state ;
	wire \mchip.row_sel[4].col_sel[2].tile_state.refresh ;
	wire \mchip.row_sel[4].col_sel[2].tile_state.rst ;
	reg \mchip.row_sel[4].col_sel[2].tile_state.state ;
	reg \mchip.row_sel[4].col_sel[2].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[4].col_sel[2].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[4].col_sel[3].tile.bottom ;
	wire [9:0] \mchip.row_sel[4].col_sel[3].tile.h_idx ;
	wire [9:0] \mchip.row_sel[4].col_sel[3].tile.left ;
	wire [9:0] \mchip.row_sel[4].col_sel[3].tile.right ;
	wire [9:0] \mchip.row_sel[4].col_sel[3].tile.top ;
	wire [9:0] \mchip.row_sel[4].col_sel[3].tile.v_idx ;
	wire \mchip.row_sel[4].col_sel[3].tile_state.clk ;
	wire [2:0] \mchip.row_sel[4].col_sel[3].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[4].col_sel[3].tile_state.focus_row ;
	wire \mchip.row_sel[4].col_sel[3].tile_state.fsm_state ;
	wire \mchip.row_sel[4].col_sel[3].tile_state.lock_state ;
	wire \mchip.row_sel[4].col_sel[3].tile_state.refresh ;
	wire \mchip.row_sel[4].col_sel[3].tile_state.rst ;
	reg \mchip.row_sel[4].col_sel[3].tile_state.state ;
	reg \mchip.row_sel[4].col_sel[3].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[4].col_sel[3].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[4].col_sel[4].tile.bottom ;
	wire [9:0] \mchip.row_sel[4].col_sel[4].tile.h_idx ;
	wire [9:0] \mchip.row_sel[4].col_sel[4].tile.left ;
	wire [9:0] \mchip.row_sel[4].col_sel[4].tile.right ;
	wire [9:0] \mchip.row_sel[4].col_sel[4].tile.top ;
	wire [9:0] \mchip.row_sel[4].col_sel[4].tile.v_idx ;
	wire \mchip.row_sel[4].col_sel[4].tile_state.clk ;
	wire [2:0] \mchip.row_sel[4].col_sel[4].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[4].col_sel[4].tile_state.focus_row ;
	wire \mchip.row_sel[4].col_sel[4].tile_state.fsm_state ;
	wire \mchip.row_sel[4].col_sel[4].tile_state.lock_state ;
	wire \mchip.row_sel[4].col_sel[4].tile_state.refresh ;
	wire \mchip.row_sel[4].col_sel[4].tile_state.rst ;
	reg \mchip.row_sel[4].col_sel[4].tile_state.state ;
	reg \mchip.row_sel[4].col_sel[4].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[4].col_sel[4].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[4].col_sel[5].tile.bottom ;
	wire [9:0] \mchip.row_sel[4].col_sel[5].tile.h_idx ;
	wire [9:0] \mchip.row_sel[4].col_sel[5].tile.left ;
	wire [9:0] \mchip.row_sel[4].col_sel[5].tile.right ;
	wire [9:0] \mchip.row_sel[4].col_sel[5].tile.top ;
	wire [9:0] \mchip.row_sel[4].col_sel[5].tile.v_idx ;
	wire \mchip.row_sel[4].col_sel[5].tile_state.clk ;
	wire [2:0] \mchip.row_sel[4].col_sel[5].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[4].col_sel[5].tile_state.focus_row ;
	wire \mchip.row_sel[4].col_sel[5].tile_state.fsm_state ;
	wire \mchip.row_sel[4].col_sel[5].tile_state.lock_state ;
	wire \mchip.row_sel[4].col_sel[5].tile_state.refresh ;
	wire \mchip.row_sel[4].col_sel[5].tile_state.rst ;
	reg \mchip.row_sel[4].col_sel[5].tile_state.state ;
	reg \mchip.row_sel[4].col_sel[5].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[4].col_sel[5].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[4].col_sel[6].tile.bottom ;
	wire [9:0] \mchip.row_sel[4].col_sel[6].tile.h_idx ;
	wire [9:0] \mchip.row_sel[4].col_sel[6].tile.left ;
	wire [9:0] \mchip.row_sel[4].col_sel[6].tile.right ;
	wire [9:0] \mchip.row_sel[4].col_sel[6].tile.top ;
	wire [9:0] \mchip.row_sel[4].col_sel[6].tile.v_idx ;
	wire \mchip.row_sel[4].col_sel[6].tile_state.clk ;
	wire [2:0] \mchip.row_sel[4].col_sel[6].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[4].col_sel[6].tile_state.focus_row ;
	wire \mchip.row_sel[4].col_sel[6].tile_state.fsm_state ;
	wire \mchip.row_sel[4].col_sel[6].tile_state.lock_state ;
	wire \mchip.row_sel[4].col_sel[6].tile_state.refresh ;
	wire \mchip.row_sel[4].col_sel[6].tile_state.rst ;
	reg \mchip.row_sel[4].col_sel[6].tile_state.state ;
	reg \mchip.row_sel[4].col_sel[6].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[4].col_sel[6].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[4].col_sel[7].tile.bottom ;
	wire [9:0] \mchip.row_sel[4].col_sel[7].tile.h_idx ;
	wire [9:0] \mchip.row_sel[4].col_sel[7].tile.left ;
	wire [9:0] \mchip.row_sel[4].col_sel[7].tile.right ;
	wire [9:0] \mchip.row_sel[4].col_sel[7].tile.top ;
	wire [9:0] \mchip.row_sel[4].col_sel[7].tile.v_idx ;
	wire \mchip.row_sel[4].col_sel[7].tile_state.clk ;
	wire [2:0] \mchip.row_sel[4].col_sel[7].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[4].col_sel[7].tile_state.focus_row ;
	wire \mchip.row_sel[4].col_sel[7].tile_state.fsm_state ;
	wire \mchip.row_sel[4].col_sel[7].tile_state.lock_state ;
	wire \mchip.row_sel[4].col_sel[7].tile_state.refresh ;
	wire \mchip.row_sel[4].col_sel[7].tile_state.rst ;
	reg \mchip.row_sel[4].col_sel[7].tile_state.state ;
	reg \mchip.row_sel[4].col_sel[7].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[4].col_sel[7].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[5].col_sel[0].tile.bottom ;
	wire [9:0] \mchip.row_sel[5].col_sel[0].tile.h_idx ;
	wire [9:0] \mchip.row_sel[5].col_sel[0].tile.left ;
	wire [9:0] \mchip.row_sel[5].col_sel[0].tile.right ;
	wire [9:0] \mchip.row_sel[5].col_sel[0].tile.top ;
	wire [9:0] \mchip.row_sel[5].col_sel[0].tile.v_idx ;
	wire \mchip.row_sel[5].col_sel[0].tile_state.clk ;
	wire [2:0] \mchip.row_sel[5].col_sel[0].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[5].col_sel[0].tile_state.focus_row ;
	wire \mchip.row_sel[5].col_sel[0].tile_state.fsm_state ;
	wire \mchip.row_sel[5].col_sel[0].tile_state.lock_state ;
	wire \mchip.row_sel[5].col_sel[0].tile_state.refresh ;
	wire \mchip.row_sel[5].col_sel[0].tile_state.rst ;
	reg \mchip.row_sel[5].col_sel[0].tile_state.state ;
	reg \mchip.row_sel[5].col_sel[0].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[5].col_sel[0].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[5].col_sel[1].tile.bottom ;
	wire [9:0] \mchip.row_sel[5].col_sel[1].tile.h_idx ;
	wire [9:0] \mchip.row_sel[5].col_sel[1].tile.left ;
	wire [9:0] \mchip.row_sel[5].col_sel[1].tile.right ;
	wire [9:0] \mchip.row_sel[5].col_sel[1].tile.top ;
	wire [9:0] \mchip.row_sel[5].col_sel[1].tile.v_idx ;
	wire \mchip.row_sel[5].col_sel[1].tile_state.clk ;
	wire [2:0] \mchip.row_sel[5].col_sel[1].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[5].col_sel[1].tile_state.focus_row ;
	wire \mchip.row_sel[5].col_sel[1].tile_state.fsm_state ;
	wire \mchip.row_sel[5].col_sel[1].tile_state.lock_state ;
	wire \mchip.row_sel[5].col_sel[1].tile_state.refresh ;
	wire \mchip.row_sel[5].col_sel[1].tile_state.rst ;
	reg \mchip.row_sel[5].col_sel[1].tile_state.state ;
	reg \mchip.row_sel[5].col_sel[1].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[5].col_sel[1].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[5].col_sel[2].tile.bottom ;
	wire [9:0] \mchip.row_sel[5].col_sel[2].tile.h_idx ;
	wire [9:0] \mchip.row_sel[5].col_sel[2].tile.left ;
	wire [9:0] \mchip.row_sel[5].col_sel[2].tile.right ;
	wire [9:0] \mchip.row_sel[5].col_sel[2].tile.top ;
	wire [9:0] \mchip.row_sel[5].col_sel[2].tile.v_idx ;
	wire \mchip.row_sel[5].col_sel[2].tile_state.clk ;
	wire [2:0] \mchip.row_sel[5].col_sel[2].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[5].col_sel[2].tile_state.focus_row ;
	wire \mchip.row_sel[5].col_sel[2].tile_state.fsm_state ;
	wire \mchip.row_sel[5].col_sel[2].tile_state.lock_state ;
	wire \mchip.row_sel[5].col_sel[2].tile_state.refresh ;
	wire \mchip.row_sel[5].col_sel[2].tile_state.rst ;
	reg \mchip.row_sel[5].col_sel[2].tile_state.state ;
	reg \mchip.row_sel[5].col_sel[2].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[5].col_sel[2].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[5].col_sel[3].tile.bottom ;
	wire [9:0] \mchip.row_sel[5].col_sel[3].tile.h_idx ;
	wire [9:0] \mchip.row_sel[5].col_sel[3].tile.left ;
	wire [9:0] \mchip.row_sel[5].col_sel[3].tile.right ;
	wire [9:0] \mchip.row_sel[5].col_sel[3].tile.top ;
	wire [9:0] \mchip.row_sel[5].col_sel[3].tile.v_idx ;
	wire \mchip.row_sel[5].col_sel[3].tile_state.clk ;
	wire [2:0] \mchip.row_sel[5].col_sel[3].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[5].col_sel[3].tile_state.focus_row ;
	wire \mchip.row_sel[5].col_sel[3].tile_state.fsm_state ;
	wire \mchip.row_sel[5].col_sel[3].tile_state.lock_state ;
	wire \mchip.row_sel[5].col_sel[3].tile_state.refresh ;
	wire \mchip.row_sel[5].col_sel[3].tile_state.rst ;
	reg \mchip.row_sel[5].col_sel[3].tile_state.state ;
	reg \mchip.row_sel[5].col_sel[3].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[5].col_sel[3].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[5].col_sel[4].tile.bottom ;
	wire [9:0] \mchip.row_sel[5].col_sel[4].tile.h_idx ;
	wire [9:0] \mchip.row_sel[5].col_sel[4].tile.left ;
	wire [9:0] \mchip.row_sel[5].col_sel[4].tile.right ;
	wire [9:0] \mchip.row_sel[5].col_sel[4].tile.top ;
	wire [9:0] \mchip.row_sel[5].col_sel[4].tile.v_idx ;
	wire \mchip.row_sel[5].col_sel[4].tile_state.clk ;
	wire [2:0] \mchip.row_sel[5].col_sel[4].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[5].col_sel[4].tile_state.focus_row ;
	wire \mchip.row_sel[5].col_sel[4].tile_state.fsm_state ;
	wire \mchip.row_sel[5].col_sel[4].tile_state.lock_state ;
	wire \mchip.row_sel[5].col_sel[4].tile_state.refresh ;
	wire \mchip.row_sel[5].col_sel[4].tile_state.rst ;
	reg \mchip.row_sel[5].col_sel[4].tile_state.state ;
	reg \mchip.row_sel[5].col_sel[4].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[5].col_sel[4].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[5].col_sel[5].tile.bottom ;
	wire [9:0] \mchip.row_sel[5].col_sel[5].tile.h_idx ;
	wire [9:0] \mchip.row_sel[5].col_sel[5].tile.left ;
	wire [9:0] \mchip.row_sel[5].col_sel[5].tile.right ;
	wire [9:0] \mchip.row_sel[5].col_sel[5].tile.top ;
	wire [9:0] \mchip.row_sel[5].col_sel[5].tile.v_idx ;
	wire \mchip.row_sel[5].col_sel[5].tile_state.clk ;
	wire [2:0] \mchip.row_sel[5].col_sel[5].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[5].col_sel[5].tile_state.focus_row ;
	wire \mchip.row_sel[5].col_sel[5].tile_state.fsm_state ;
	wire \mchip.row_sel[5].col_sel[5].tile_state.lock_state ;
	wire \mchip.row_sel[5].col_sel[5].tile_state.refresh ;
	wire \mchip.row_sel[5].col_sel[5].tile_state.rst ;
	reg \mchip.row_sel[5].col_sel[5].tile_state.state ;
	reg \mchip.row_sel[5].col_sel[5].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[5].col_sel[5].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[5].col_sel[6].tile.bottom ;
	wire [9:0] \mchip.row_sel[5].col_sel[6].tile.h_idx ;
	wire [9:0] \mchip.row_sel[5].col_sel[6].tile.left ;
	wire [9:0] \mchip.row_sel[5].col_sel[6].tile.right ;
	wire [9:0] \mchip.row_sel[5].col_sel[6].tile.top ;
	wire [9:0] \mchip.row_sel[5].col_sel[6].tile.v_idx ;
	wire \mchip.row_sel[5].col_sel[6].tile_state.clk ;
	wire [2:0] \mchip.row_sel[5].col_sel[6].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[5].col_sel[6].tile_state.focus_row ;
	wire \mchip.row_sel[5].col_sel[6].tile_state.fsm_state ;
	wire \mchip.row_sel[5].col_sel[6].tile_state.lock_state ;
	wire \mchip.row_sel[5].col_sel[6].tile_state.refresh ;
	wire \mchip.row_sel[5].col_sel[6].tile_state.rst ;
	reg \mchip.row_sel[5].col_sel[6].tile_state.state ;
	reg \mchip.row_sel[5].col_sel[6].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[5].col_sel[6].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[5].col_sel[7].tile.bottom ;
	wire [9:0] \mchip.row_sel[5].col_sel[7].tile.h_idx ;
	wire [9:0] \mchip.row_sel[5].col_sel[7].tile.left ;
	wire [9:0] \mchip.row_sel[5].col_sel[7].tile.right ;
	wire [9:0] \mchip.row_sel[5].col_sel[7].tile.top ;
	wire [9:0] \mchip.row_sel[5].col_sel[7].tile.v_idx ;
	wire \mchip.row_sel[5].col_sel[7].tile_state.clk ;
	wire [2:0] \mchip.row_sel[5].col_sel[7].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[5].col_sel[7].tile_state.focus_row ;
	wire \mchip.row_sel[5].col_sel[7].tile_state.fsm_state ;
	wire \mchip.row_sel[5].col_sel[7].tile_state.lock_state ;
	wire \mchip.row_sel[5].col_sel[7].tile_state.refresh ;
	wire \mchip.row_sel[5].col_sel[7].tile_state.rst ;
	reg \mchip.row_sel[5].col_sel[7].tile_state.state ;
	reg \mchip.row_sel[5].col_sel[7].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[5].col_sel[7].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[6].col_sel[0].tile.bottom ;
	wire [9:0] \mchip.row_sel[6].col_sel[0].tile.h_idx ;
	wire [9:0] \mchip.row_sel[6].col_sel[0].tile.left ;
	wire [9:0] \mchip.row_sel[6].col_sel[0].tile.right ;
	wire [9:0] \mchip.row_sel[6].col_sel[0].tile.top ;
	wire [9:0] \mchip.row_sel[6].col_sel[0].tile.v_idx ;
	wire \mchip.row_sel[6].col_sel[0].tile_state.clk ;
	wire [2:0] \mchip.row_sel[6].col_sel[0].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[6].col_sel[0].tile_state.focus_row ;
	wire \mchip.row_sel[6].col_sel[0].tile_state.fsm_state ;
	wire \mchip.row_sel[6].col_sel[0].tile_state.lock_state ;
	wire [1:0] \mchip.row_sel[6].col_sel[0].tile_state.neighbors_hori ;
	wire \mchip.row_sel[6].col_sel[0].tile_state.refresh ;
	wire \mchip.row_sel[6].col_sel[0].tile_state.rst ;
	reg \mchip.row_sel[6].col_sel[0].tile_state.state ;
	reg \mchip.row_sel[6].col_sel[0].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[6].col_sel[0].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[6].col_sel[1].tile.bottom ;
	wire [9:0] \mchip.row_sel[6].col_sel[1].tile.h_idx ;
	wire [9:0] \mchip.row_sel[6].col_sel[1].tile.left ;
	wire [9:0] \mchip.row_sel[6].col_sel[1].tile.right ;
	wire [9:0] \mchip.row_sel[6].col_sel[1].tile.top ;
	wire [9:0] \mchip.row_sel[6].col_sel[1].tile.v_idx ;
	wire \mchip.row_sel[6].col_sel[1].tile_state.clk ;
	wire [2:0] \mchip.row_sel[6].col_sel[1].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[6].col_sel[1].tile_state.focus_row ;
	wire \mchip.row_sel[6].col_sel[1].tile_state.fsm_state ;
	wire \mchip.row_sel[6].col_sel[1].tile_state.lock_state ;
	wire \mchip.row_sel[6].col_sel[1].tile_state.refresh ;
	wire \mchip.row_sel[6].col_sel[1].tile_state.rst ;
	reg \mchip.row_sel[6].col_sel[1].tile_state.state ;
	reg \mchip.row_sel[6].col_sel[1].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[6].col_sel[1].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[6].col_sel[2].tile.bottom ;
	wire [9:0] \mchip.row_sel[6].col_sel[2].tile.h_idx ;
	wire [9:0] \mchip.row_sel[6].col_sel[2].tile.left ;
	wire [9:0] \mchip.row_sel[6].col_sel[2].tile.right ;
	wire [9:0] \mchip.row_sel[6].col_sel[2].tile.top ;
	wire [9:0] \mchip.row_sel[6].col_sel[2].tile.v_idx ;
	wire \mchip.row_sel[6].col_sel[2].tile_state.clk ;
	wire [2:0] \mchip.row_sel[6].col_sel[2].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[6].col_sel[2].tile_state.focus_row ;
	wire \mchip.row_sel[6].col_sel[2].tile_state.fsm_state ;
	wire \mchip.row_sel[6].col_sel[2].tile_state.lock_state ;
	wire \mchip.row_sel[6].col_sel[2].tile_state.refresh ;
	wire \mchip.row_sel[6].col_sel[2].tile_state.rst ;
	reg \mchip.row_sel[6].col_sel[2].tile_state.state ;
	reg \mchip.row_sel[6].col_sel[2].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[6].col_sel[2].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[6].col_sel[3].tile.bottom ;
	wire [9:0] \mchip.row_sel[6].col_sel[3].tile.h_idx ;
	wire [9:0] \mchip.row_sel[6].col_sel[3].tile.left ;
	wire [9:0] \mchip.row_sel[6].col_sel[3].tile.right ;
	wire [9:0] \mchip.row_sel[6].col_sel[3].tile.top ;
	wire [9:0] \mchip.row_sel[6].col_sel[3].tile.v_idx ;
	wire \mchip.row_sel[6].col_sel[3].tile_state.clk ;
	wire [2:0] \mchip.row_sel[6].col_sel[3].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[6].col_sel[3].tile_state.focus_row ;
	wire \mchip.row_sel[6].col_sel[3].tile_state.fsm_state ;
	wire \mchip.row_sel[6].col_sel[3].tile_state.lock_state ;
	wire \mchip.row_sel[6].col_sel[3].tile_state.refresh ;
	wire \mchip.row_sel[6].col_sel[3].tile_state.rst ;
	reg \mchip.row_sel[6].col_sel[3].tile_state.state ;
	reg \mchip.row_sel[6].col_sel[3].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[6].col_sel[3].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[6].col_sel[4].tile.bottom ;
	wire [9:0] \mchip.row_sel[6].col_sel[4].tile.h_idx ;
	wire [9:0] \mchip.row_sel[6].col_sel[4].tile.left ;
	wire [9:0] \mchip.row_sel[6].col_sel[4].tile.right ;
	wire [9:0] \mchip.row_sel[6].col_sel[4].tile.top ;
	wire [9:0] \mchip.row_sel[6].col_sel[4].tile.v_idx ;
	wire \mchip.row_sel[6].col_sel[4].tile_state.clk ;
	wire [2:0] \mchip.row_sel[6].col_sel[4].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[6].col_sel[4].tile_state.focus_row ;
	wire \mchip.row_sel[6].col_sel[4].tile_state.fsm_state ;
	wire \mchip.row_sel[6].col_sel[4].tile_state.lock_state ;
	wire \mchip.row_sel[6].col_sel[4].tile_state.refresh ;
	wire \mchip.row_sel[6].col_sel[4].tile_state.rst ;
	reg \mchip.row_sel[6].col_sel[4].tile_state.state ;
	reg \mchip.row_sel[6].col_sel[4].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[6].col_sel[4].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[6].col_sel[5].tile.bottom ;
	wire [9:0] \mchip.row_sel[6].col_sel[5].tile.h_idx ;
	wire [9:0] \mchip.row_sel[6].col_sel[5].tile.left ;
	wire [9:0] \mchip.row_sel[6].col_sel[5].tile.right ;
	wire [9:0] \mchip.row_sel[6].col_sel[5].tile.top ;
	wire [9:0] \mchip.row_sel[6].col_sel[5].tile.v_idx ;
	wire \mchip.row_sel[6].col_sel[5].tile_state.clk ;
	wire [2:0] \mchip.row_sel[6].col_sel[5].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[6].col_sel[5].tile_state.focus_row ;
	wire \mchip.row_sel[6].col_sel[5].tile_state.fsm_state ;
	wire \mchip.row_sel[6].col_sel[5].tile_state.lock_state ;
	wire \mchip.row_sel[6].col_sel[5].tile_state.refresh ;
	wire \mchip.row_sel[6].col_sel[5].tile_state.rst ;
	reg \mchip.row_sel[6].col_sel[5].tile_state.state ;
	reg \mchip.row_sel[6].col_sel[5].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[6].col_sel[5].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[6].col_sel[6].tile.bottom ;
	wire [9:0] \mchip.row_sel[6].col_sel[6].tile.h_idx ;
	wire [9:0] \mchip.row_sel[6].col_sel[6].tile.left ;
	wire [9:0] \mchip.row_sel[6].col_sel[6].tile.right ;
	wire [9:0] \mchip.row_sel[6].col_sel[6].tile.top ;
	wire [9:0] \mchip.row_sel[6].col_sel[6].tile.v_idx ;
	wire \mchip.row_sel[6].col_sel[6].tile_state.clk ;
	wire [2:0] \mchip.row_sel[6].col_sel[6].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[6].col_sel[6].tile_state.focus_row ;
	wire \mchip.row_sel[6].col_sel[6].tile_state.fsm_state ;
	wire \mchip.row_sel[6].col_sel[6].tile_state.lock_state ;
	wire \mchip.row_sel[6].col_sel[6].tile_state.refresh ;
	wire \mchip.row_sel[6].col_sel[6].tile_state.rst ;
	reg \mchip.row_sel[6].col_sel[6].tile_state.state ;
	reg \mchip.row_sel[6].col_sel[6].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[6].col_sel[6].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[6].col_sel[7].tile.bottom ;
	wire [9:0] \mchip.row_sel[6].col_sel[7].tile.h_idx ;
	wire [9:0] \mchip.row_sel[6].col_sel[7].tile.left ;
	wire [9:0] \mchip.row_sel[6].col_sel[7].tile.right ;
	wire [9:0] \mchip.row_sel[6].col_sel[7].tile.top ;
	wire [9:0] \mchip.row_sel[6].col_sel[7].tile.v_idx ;
	wire \mchip.row_sel[6].col_sel[7].tile_state.clk ;
	wire [2:0] \mchip.row_sel[6].col_sel[7].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[6].col_sel[7].tile_state.focus_row ;
	wire \mchip.row_sel[6].col_sel[7].tile_state.fsm_state ;
	wire \mchip.row_sel[6].col_sel[7].tile_state.lock_state ;
	wire [1:0] \mchip.row_sel[6].col_sel[7].tile_state.neighbors_hori ;
	wire \mchip.row_sel[6].col_sel[7].tile_state.refresh ;
	wire \mchip.row_sel[6].col_sel[7].tile_state.rst ;
	reg \mchip.row_sel[6].col_sel[7].tile_state.state ;
	reg \mchip.row_sel[6].col_sel[7].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[6].col_sel[7].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[7].col_sel[0].tile.bottom ;
	wire [9:0] \mchip.row_sel[7].col_sel[0].tile.h_idx ;
	wire [9:0] \mchip.row_sel[7].col_sel[0].tile.left ;
	wire [9:0] \mchip.row_sel[7].col_sel[0].tile.right ;
	wire [9:0] \mchip.row_sel[7].col_sel[0].tile.top ;
	wire [9:0] \mchip.row_sel[7].col_sel[0].tile.v_idx ;
	wire \mchip.row_sel[7].col_sel[0].tile_state.clk ;
	wire [2:0] \mchip.row_sel[7].col_sel[0].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[7].col_sel[0].tile_state.focus_row ;
	wire \mchip.row_sel[7].col_sel[0].tile_state.fsm_state ;
	wire \mchip.row_sel[7].col_sel[0].tile_state.lock_state ;
	wire \mchip.row_sel[7].col_sel[0].tile_state.refresh ;
	wire \mchip.row_sel[7].col_sel[0].tile_state.rst ;
	reg \mchip.row_sel[7].col_sel[0].tile_state.state ;
	reg \mchip.row_sel[7].col_sel[0].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[7].col_sel[0].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[7].col_sel[1].tile.bottom ;
	wire [9:0] \mchip.row_sel[7].col_sel[1].tile.h_idx ;
	wire [9:0] \mchip.row_sel[7].col_sel[1].tile.left ;
	wire [9:0] \mchip.row_sel[7].col_sel[1].tile.right ;
	wire [9:0] \mchip.row_sel[7].col_sel[1].tile.top ;
	wire [9:0] \mchip.row_sel[7].col_sel[1].tile.v_idx ;
	wire \mchip.row_sel[7].col_sel[1].tile_state.clk ;
	wire [2:0] \mchip.row_sel[7].col_sel[1].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[7].col_sel[1].tile_state.focus_row ;
	wire \mchip.row_sel[7].col_sel[1].tile_state.fsm_state ;
	wire \mchip.row_sel[7].col_sel[1].tile_state.lock_state ;
	wire [1:0] \mchip.row_sel[7].col_sel[1].tile_state.neighbors_vert ;
	wire \mchip.row_sel[7].col_sel[1].tile_state.refresh ;
	wire \mchip.row_sel[7].col_sel[1].tile_state.rst ;
	reg \mchip.row_sel[7].col_sel[1].tile_state.state ;
	reg \mchip.row_sel[7].col_sel[1].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[7].col_sel[1].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[7].col_sel[2].tile.bottom ;
	wire [9:0] \mchip.row_sel[7].col_sel[2].tile.h_idx ;
	wire [9:0] \mchip.row_sel[7].col_sel[2].tile.left ;
	wire [9:0] \mchip.row_sel[7].col_sel[2].tile.right ;
	wire [9:0] \mchip.row_sel[7].col_sel[2].tile.top ;
	wire [9:0] \mchip.row_sel[7].col_sel[2].tile.v_idx ;
	wire \mchip.row_sel[7].col_sel[2].tile_state.clk ;
	wire [2:0] \mchip.row_sel[7].col_sel[2].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[7].col_sel[2].tile_state.focus_row ;
	wire \mchip.row_sel[7].col_sel[2].tile_state.fsm_state ;
	wire \mchip.row_sel[7].col_sel[2].tile_state.lock_state ;
	wire \mchip.row_sel[7].col_sel[2].tile_state.refresh ;
	wire \mchip.row_sel[7].col_sel[2].tile_state.rst ;
	reg \mchip.row_sel[7].col_sel[2].tile_state.state ;
	reg \mchip.row_sel[7].col_sel[2].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[7].col_sel[2].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[7].col_sel[3].tile.bottom ;
	wire [9:0] \mchip.row_sel[7].col_sel[3].tile.h_idx ;
	wire [9:0] \mchip.row_sel[7].col_sel[3].tile.left ;
	wire [9:0] \mchip.row_sel[7].col_sel[3].tile.right ;
	wire [9:0] \mchip.row_sel[7].col_sel[3].tile.top ;
	wire [9:0] \mchip.row_sel[7].col_sel[3].tile.v_idx ;
	wire \mchip.row_sel[7].col_sel[3].tile_state.clk ;
	wire [2:0] \mchip.row_sel[7].col_sel[3].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[7].col_sel[3].tile_state.focus_row ;
	wire \mchip.row_sel[7].col_sel[3].tile_state.fsm_state ;
	wire \mchip.row_sel[7].col_sel[3].tile_state.lock_state ;
	wire \mchip.row_sel[7].col_sel[3].tile_state.refresh ;
	wire \mchip.row_sel[7].col_sel[3].tile_state.rst ;
	reg \mchip.row_sel[7].col_sel[3].tile_state.state ;
	reg \mchip.row_sel[7].col_sel[3].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[7].col_sel[3].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[7].col_sel[4].tile.bottom ;
	wire [9:0] \mchip.row_sel[7].col_sel[4].tile.h_idx ;
	wire [9:0] \mchip.row_sel[7].col_sel[4].tile.left ;
	wire [9:0] \mchip.row_sel[7].col_sel[4].tile.right ;
	wire [9:0] \mchip.row_sel[7].col_sel[4].tile.top ;
	wire [9:0] \mchip.row_sel[7].col_sel[4].tile.v_idx ;
	wire \mchip.row_sel[7].col_sel[4].tile_state.clk ;
	wire [2:0] \mchip.row_sel[7].col_sel[4].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[7].col_sel[4].tile_state.focus_row ;
	wire \mchip.row_sel[7].col_sel[4].tile_state.fsm_state ;
	wire \mchip.row_sel[7].col_sel[4].tile_state.lock_state ;
	wire \mchip.row_sel[7].col_sel[4].tile_state.refresh ;
	wire \mchip.row_sel[7].col_sel[4].tile_state.rst ;
	reg \mchip.row_sel[7].col_sel[4].tile_state.state ;
	reg \mchip.row_sel[7].col_sel[4].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[7].col_sel[4].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[7].col_sel[5].tile.bottom ;
	wire [9:0] \mchip.row_sel[7].col_sel[5].tile.h_idx ;
	wire [9:0] \mchip.row_sel[7].col_sel[5].tile.left ;
	wire [9:0] \mchip.row_sel[7].col_sel[5].tile.right ;
	wire [9:0] \mchip.row_sel[7].col_sel[5].tile.top ;
	wire [9:0] \mchip.row_sel[7].col_sel[5].tile.v_idx ;
	wire \mchip.row_sel[7].col_sel[5].tile_state.clk ;
	wire [2:0] \mchip.row_sel[7].col_sel[5].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[7].col_sel[5].tile_state.focus_row ;
	wire \mchip.row_sel[7].col_sel[5].tile_state.fsm_state ;
	wire \mchip.row_sel[7].col_sel[5].tile_state.lock_state ;
	wire \mchip.row_sel[7].col_sel[5].tile_state.refresh ;
	wire \mchip.row_sel[7].col_sel[5].tile_state.rst ;
	reg \mchip.row_sel[7].col_sel[5].tile_state.state ;
	reg \mchip.row_sel[7].col_sel[5].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[7].col_sel[5].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[7].col_sel[6].tile.bottom ;
	wire [9:0] \mchip.row_sel[7].col_sel[6].tile.h_idx ;
	wire [9:0] \mchip.row_sel[7].col_sel[6].tile.left ;
	wire [9:0] \mchip.row_sel[7].col_sel[6].tile.right ;
	wire [9:0] \mchip.row_sel[7].col_sel[6].tile.top ;
	wire [9:0] \mchip.row_sel[7].col_sel[6].tile.v_idx ;
	wire \mchip.row_sel[7].col_sel[6].tile_state.clk ;
	wire [2:0] \mchip.row_sel[7].col_sel[6].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[7].col_sel[6].tile_state.focus_row ;
	wire \mchip.row_sel[7].col_sel[6].tile_state.fsm_state ;
	wire \mchip.row_sel[7].col_sel[6].tile_state.lock_state ;
	wire [1:0] \mchip.row_sel[7].col_sel[6].tile_state.neighbors_vert ;
	wire \mchip.row_sel[7].col_sel[6].tile_state.refresh ;
	wire \mchip.row_sel[7].col_sel[6].tile_state.rst ;
	reg \mchip.row_sel[7].col_sel[6].tile_state.state ;
	reg \mchip.row_sel[7].col_sel[6].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[7].col_sel[6].tile_state.tile_states ;
	wire [9:0] \mchip.row_sel[7].col_sel[7].tile.bottom ;
	wire [9:0] \mchip.row_sel[7].col_sel[7].tile.h_idx ;
	wire [9:0] \mchip.row_sel[7].col_sel[7].tile.left ;
	wire [9:0] \mchip.row_sel[7].col_sel[7].tile.right ;
	wire [9:0] \mchip.row_sel[7].col_sel[7].tile.top ;
	wire [9:0] \mchip.row_sel[7].col_sel[7].tile.v_idx ;
	wire \mchip.row_sel[7].col_sel[7].tile_state.clk ;
	wire [2:0] \mchip.row_sel[7].col_sel[7].tile_state.focus_col ;
	wire [2:0] \mchip.row_sel[7].col_sel[7].tile_state.focus_row ;
	wire \mchip.row_sel[7].col_sel[7].tile_state.fsm_state ;
	wire \mchip.row_sel[7].col_sel[7].tile_state.lock_state ;
	wire \mchip.row_sel[7].col_sel[7].tile_state.refresh ;
	wire \mchip.row_sel[7].col_sel[7].tile_state.rst ;
	reg \mchip.row_sel[7].col_sel[7].tile_state.state ;
	reg \mchip.row_sel[7].col_sel[7].tile_state.state_locked ;
	wire [63:0] \mchip.row_sel[7].col_sel[7].tile_state.tile_states ;
	wire [63:0] \mchip.tile_states ;
	wire [639:0] \mchip.top ;
	wire [9:0] \mchip.v_idx ;
	wire \mchip.vga.clk ;
	reg [31:0] \mchip.vga.frame_count ;
	reg \mchip.vga.frame_end ;
	reg [9:0] \mchip.vga.h_idx ;
	reg \mchip.vga.hsync ;
	reg \mchip.vga.refresh ;
	wire \mchip.vga.rst ;
	reg [9:0] \mchip.vga.v_idx ;
	reg \mchip.vga.vsync ;
	wire \mchip.vsync ;
	assign _1730_ = \mchip.fsm_state  | ~\mchip.row_sel[1].col_sel[5].tile_state.state ;
	assign _0136_ = \mchip.lock_state  & ~_1730_;
	assign _1731_ = ~\mchip.vga.refresh ;
	assign _1732_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[1].col_sel[5].tile_state.state_locked );
	assign _0050_ = ~(_1732_ | _0136_);
	assign _1733_ = \mchip.fsm_state  | ~\mchip.row_sel[2].col_sel[5].tile_state.state ;
	assign _0152_ = \mchip.lock_state  & ~_1733_;
	assign _1734_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[2].col_sel[5].tile_state.state_locked );
	assign _0042_ = ~(_1734_ | _0152_);
	assign _1735_ = \mchip.fsm_state  | ~\mchip.row_sel[4].col_sel[1].tile_state.state ;
	assign _0176_ = \mchip.lock_state  & ~_1735_;
	assign _1736_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[4].col_sel[1].tile_state.state_locked );
	assign _0030_ = ~(_1736_ | _0176_);
	assign _1737_ = \mchip.fsm_state  | ~\mchip.row_sel[4].col_sel[2].tile_state.state ;
	assign _0178_ = \mchip.lock_state  & ~_1737_;
	assign _1738_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[4].col_sel[2].tile_state.state_locked );
	assign _0029_ = ~(_1738_ | _0178_);
	assign _1739_ = \mchip.fsm_state  | ~\mchip.row_sel[1].col_sel[0].tile_state.state ;
	assign _0126_ = \mchip.lock_state  & ~_1739_;
	assign _1740_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[1].col_sel[0].tile_state.state_locked );
	assign _0055_ = ~(_1740_ | _0126_);
	assign _1741_ = \mchip.fsm_state  | ~\mchip.row_sel[0].col_sel[5].tile_state.state ;
	assign _0120_ = \mchip.lock_state  & ~_1741_;
	assign _1742_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[0].col_sel[5].tile_state.state_locked );
	assign _0058_ = ~(_1742_ | _0120_);
	assign _1743_ = \mchip.fsm_state  | ~\mchip.row_sel[0].col_sel[6].tile_state.state ;
	assign _0122_ = \mchip.lock_state  & ~_1743_;
	assign _1744_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[0].col_sel[6].tile_state.state_locked );
	assign _0057_ = ~(_1744_ | _0122_);
	assign _1745_ = ~(\mchip.vga.h_idx [8] & \mchip.vga.h_idx [7]);
	assign _1746_ = \mchip.vga.h_idx [6] | \mchip.vga.h_idx [5];
	assign _1747_ = \mchip.vga.h_idx [7] | ~\mchip.vga.h_idx [8];
	assign _1748_ = _1746_ & ~_1747_;
	assign _1749_ = _1745_ & ~_1748_;
	assign _1750_ = \mchip.vga.h_idx [9] & ~_1749_;
	assign _1751_ = \mchip.vga.h_idx [9] & \mchip.vga.h_idx [8];
	assign _1752_ = \mchip.vga.h_idx [1] | \mchip.vga.h_idx [4];
	assign _1753_ = \mchip.vga.h_idx [2] | \mchip.vga.h_idx [3];
	assign _1754_ = _1753_ | _1752_;
	assign _1755_ = \mchip.vga.h_idx [6] | \mchip.vga.h_idx [7];
	assign _1756_ = \mchip.vga.h_idx [0] | ~\mchip.vga.h_idx [5];
	assign _1757_ = _1756_ | _1755_;
	assign _1758_ = _1757_ | _1754_;
	assign _1759_ = _1751_ & ~_1758_;
	assign _0252_ = ~(_1759_ | _1750_);
	assign _1760_ = \mchip.fsm_state  | ~\mchip.row_sel[4].col_sel[3].tile_state.state ;
	assign _0180_ = \mchip.lock_state  & ~_1760_;
	assign _1761_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[4].col_sel[3].tile_state.state_locked );
	assign _0028_ = ~(_1761_ | _0180_);
	assign _1762_ = \mchip.fsm_state  | ~\mchip.row_sel[4].col_sel[4].tile_state.state ;
	assign _0182_ = \mchip.lock_state  & ~_1762_;
	assign _1763_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[4].col_sel[4].tile_state.state_locked );
	assign _0027_ = ~(_1763_ | _0182_);
	assign _1764_ = \mchip.fsm_state  | ~\mchip.row_sel[2].col_sel[6].tile_state.state ;
	assign _0154_ = \mchip.lock_state  & ~_1764_;
	assign _1765_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[2].col_sel[6].tile_state.state_locked );
	assign _0041_ = ~(_1765_ | _0154_);
	assign _1766_ = \mchip.fsm_state  | ~\mchip.row_sel[2].col_sel[7].tile_state.state ;
	assign _0156_ = \mchip.lock_state  & ~_1766_;
	assign _1767_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[2].col_sel[7].tile_state.state_locked );
	assign _0040_ = ~(_1767_ | _0156_);
	assign _1768_ = \mchip.fsm_state  | ~\mchip.row_sel[0].col_sel[2].tile_state.state ;
	assign _0114_ = \mchip.lock_state  & ~_1768_;
	assign _1769_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[0].col_sel[2].tile_state.state_locked );
	assign _0061_ = ~(_1769_ | _0114_);
	assign _1770_ = \mchip.fsm_state  | ~\mchip.row_sel[1].col_sel[6].tile_state.state ;
	assign _0138_ = \mchip.lock_state  & ~_1770_;
	assign _1771_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[1].col_sel[6].tile_state.state_locked );
	assign _0049_ = ~(_1771_ | _0138_);
	assign _1772_ = \mchip.fsm_state  | ~\mchip.row_sel[1].col_sel[7].tile_state.state ;
	assign _0140_ = \mchip.lock_state  & ~_1772_;
	assign _1773_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[1].col_sel[7].tile_state.state_locked );
	assign _0048_ = ~(_1773_ | _0140_);
	assign _1774_ = \mchip.fsm_state  | ~\mchip.row_sel[4].col_sel[5].tile_state.state ;
	assign _0184_ = \mchip.lock_state  & ~_1774_;
	assign _1775_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[4].col_sel[5].tile_state.state_locked );
	assign _0026_ = ~(_1775_ | _0184_);
	assign _1776_ = \mchip.fsm_state  | ~\mchip.row_sel[4].col_sel[6].tile_state.state ;
	assign _0186_ = \mchip.lock_state  & ~_1776_;
	assign _1777_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[4].col_sel[6].tile_state.state_locked );
	assign _0025_ = ~(_1777_ | _0186_);
	assign _1778_ = \mchip.fsm_state  | ~\mchip.row_sel[3].col_sel[0].tile_state.state ;
	assign _0158_ = \mchip.lock_state  & ~_1778_;
	assign _1779_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[3].col_sel[0].tile_state.state_locked );
	assign _0039_ = ~(_1779_ | _0158_);
	assign _1780_ = \mchip.fsm_state  | ~\mchip.row_sel[3].col_sel[1].tile_state.state ;
	assign _0160_ = \mchip.lock_state  & ~_1780_;
	assign _1781_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[3].col_sel[1].tile_state.state_locked );
	assign _0038_ = ~(_1781_ | _0160_);
	assign _2115_[0] = ~\mchip.vga.h_idx [0];
	assign _1782_ = \mchip.fsm_state  | ~\mchip.row_sel[4].col_sel[7].tile_state.state ;
	assign _0188_ = \mchip.lock_state  & ~_1782_;
	assign _1783_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[4].col_sel[7].tile_state.state_locked );
	assign _0024_ = ~(_1783_ | _0188_);
	assign _1784_ = \mchip.fsm_state  | ~\mchip.row_sel[1].col_sel[1].tile_state.state ;
	assign _0128_ = \mchip.lock_state  & ~_1784_;
	assign _1785_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[1].col_sel[1].tile_state.state_locked );
	assign _0054_ = ~(_1785_ | _0128_);
	assign _1786_ = \mchip.fsm_state  | ~\mchip.row_sel[1].col_sel[2].tile_state.state ;
	assign _0130_ = \mchip.lock_state  & ~_1786_;
	assign _1787_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[1].col_sel[2].tile_state.state_locked );
	assign _0053_ = ~(_1787_ | _0130_);
	assign _1788_ = \mchip.fsm_state  | ~\mchip.row_sel[5].col_sel[0].tile_state.state ;
	assign _0190_ = \mchip.lock_state  & ~_1788_;
	assign _1789_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[5].col_sel[0].tile_state.state_locked );
	assign _0023_ = ~(_1789_ | _0190_);
	assign _1790_ = \mchip.fsm_state  | ~\mchip.row_sel[5].col_sel[1].tile_state.state ;
	assign _0192_ = \mchip.lock_state  & ~_1790_;
	assign _1791_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[5].col_sel[1].tile_state.state_locked );
	assign _0022_ = ~(_1791_ | _0192_);
	assign _1792_ = \mchip.fsm_state  | ~\mchip.row_sel[3].col_sel[2].tile_state.state ;
	assign _0162_ = \mchip.lock_state  & ~_1792_;
	assign _1793_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[3].col_sel[2].tile_state.state_locked );
	assign _0037_ = ~(_1793_ | _0162_);
	assign _1794_ = \mchip.fsm_state  | ~\mchip.row_sel[2].col_sel[0].tile_state.state ;
	assign _0142_ = \mchip.lock_state  & ~_1794_;
	assign _1795_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[2].col_sel[0].tile_state.state_locked );
	assign _0047_ = ~(_1795_ | _0142_);
	assign _1796_ = \mchip.fsm_state  | ~\mchip.row_sel[2].col_sel[1].tile_state.state ;
	assign _0144_ = \mchip.lock_state  & ~_1796_;
	assign _1797_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[2].col_sel[1].tile_state.state_locked );
	assign _0046_ = ~(_1797_ | _0144_);
	assign _1798_ = \mchip.fsm_state  | ~\mchip.row_sel[5].col_sel[2].tile_state.state ;
	assign _0194_ = \mchip.lock_state  & ~_1798_;
	assign _1799_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[5].col_sel[2].tile_state.state_locked );
	assign _0021_ = ~(_1799_ | _0194_);
	assign _1800_ = \mchip.fsm_state  | ~\mchip.row_sel[5].col_sel[3].tile_state.state ;
	assign _0196_ = \mchip.lock_state  & ~_1800_;
	assign _1801_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[5].col_sel[3].tile_state.state_locked );
	assign _0020_ = ~(_1801_ | _0196_);
	assign _1802_ = \mchip.fsm_state  | ~\mchip.row_sel[0].col_sel[3].tile_state.state ;
	assign _0116_ = \mchip.lock_state  & ~_1802_;
	assign _1803_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[0].col_sel[3].tile_state.state_locked );
	assign _0060_ = ~(_1803_ | _0116_);
	assign _1804_ = \mchip.fsm_state  | ~\mchip.row_sel[0].col_sel[4].tile_state.state ;
	assign _0118_ = \mchip.lock_state  & ~_1804_;
	assign _1805_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[0].col_sel[4].tile_state.state_locked );
	assign _0059_ = ~(_1805_ | _0118_);
	assign _1806_ = \mchip.fsm_state  | ~\mchip.row_sel[0].col_sel[7].tile_state.state ;
	assign _0124_ = \mchip.lock_state  & ~_1806_;
	assign _1807_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[0].col_sel[7].tile_state.state_locked );
	assign _0056_ = ~(_1807_ | _0124_);
	assign _1808_ = \mchip.fsm_state  | ~\mchip.row_sel[3].col_sel[3].tile_state.state ;
	assign _0164_ = \mchip.lock_state  & ~_1808_;
	assign _1809_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[3].col_sel[3].tile_state.state_locked );
	assign _0036_ = ~(_1809_ | _0164_);
	assign _1810_ = \mchip.fsm_state  | ~\mchip.row_sel[3].col_sel[4].tile_state.state ;
	assign _0166_ = \mchip.lock_state  & ~_1810_;
	assign _1811_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[3].col_sel[4].tile_state.state_locked );
	assign _0035_ = ~(_1811_ | _0166_);
	assign _1812_ = \mchip.fsm_state  | ~\mchip.row_sel[5].col_sel[4].tile_state.state ;
	assign _0198_ = \mchip.lock_state  & ~_1812_;
	assign _1813_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[5].col_sel[4].tile_state.state_locked );
	assign _0019_ = ~(_1813_ | _0198_);
	assign _1814_ = \mchip.fsm_state  | ~\mchip.row_sel[2].col_sel[2].tile_state.state ;
	assign _0146_ = \mchip.lock_state  & ~_1814_;
	assign _1815_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[2].col_sel[2].tile_state.state_locked );
	assign _0045_ = ~(_1815_ | _0146_);
	assign _1816_ = \mchip.fsm_state  | ~\mchip.row_sel[5].col_sel[5].tile_state.state ;
	assign _0200_ = \mchip.lock_state  & ~_1816_;
	assign _1817_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[5].col_sel[5].tile_state.state_locked );
	assign _0018_ = ~(_1817_ | _0200_);
	assign _1818_ = \mchip.fsm_state  | ~\mchip.row_sel[5].col_sel[6].tile_state.state ;
	assign _0202_ = \mchip.lock_state  & ~_1818_;
	assign _1819_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[5].col_sel[6].tile_state.state_locked );
	assign _0017_ = ~(_1819_ | _0202_);
	assign _1820_ = \mchip.fsm_state  | ~\mchip.row_sel[0].col_sel[0].tile_state.state ;
	assign _0110_ = \mchip.lock_state  & ~_1820_;
	assign _1821_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[0].col_sel[0].tile_state.state_locked );
	assign _0063_ = ~(_1821_ | _0110_);
	assign _0070_ = \mchip.btn4_sync  & \mchip.vga.frame_end ;
	assign _1822_ = \mchip.fsm_state  | ~\mchip.row_sel[0].col_sel[1].tile_state.state ;
	assign _0112_ = \mchip.lock_state  & ~_1822_;
	assign _1823_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[0].col_sel[1].tile_state.state_locked );
	assign _0062_ = ~(_1823_ | _0112_);
	assign _1824_ = \mchip.fsm_state  | ~\mchip.row_sel[3].col_sel[5].tile_state.state ;
	assign _0168_ = \mchip.lock_state  & ~_1824_;
	assign _1825_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[3].col_sel[5].tile_state.state_locked );
	assign _0034_ = ~(_1825_ | _0168_);
	assign _1826_ = \mchip.fsm_state  | ~\mchip.row_sel[3].col_sel[6].tile_state.state ;
	assign _0170_ = \mchip.lock_state  & ~_1826_;
	assign _1827_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[3].col_sel[6].tile_state.state_locked );
	assign _0033_ = ~(_1827_ | _0170_);
	assign _1828_ = \mchip.fsm_state  | ~\mchip.row_sel[1].col_sel[3].tile_state.state ;
	assign _0132_ = \mchip.lock_state  & ~_1828_;
	assign _1829_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[1].col_sel[3].tile_state.state_locked );
	assign _0052_ = ~(_1829_ | _0132_);
	assign _1830_ = \mchip.fsm_state  | ~\mchip.row_sel[1].col_sel[4].tile_state.state ;
	assign _0134_ = \mchip.lock_state  & ~_1830_;
	assign _1831_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[1].col_sel[4].tile_state.state_locked );
	assign _0051_ = ~(_1831_ | _0134_);
	assign _1832_ = \mchip.fsm_state  | ~\mchip.row_sel[5].col_sel[7].tile_state.state ;
	assign _0204_ = \mchip.lock_state  & ~_1832_;
	assign _1833_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[5].col_sel[7].tile_state.state_locked );
	assign _0016_ = ~(_1833_ | _0204_);
	assign _0103_ = \mchip.btn3_sync  & \mchip.vga.frame_end ;
	assign _1834_ = io_in[2] & ~io_in[3];
	assign _1835_ = _1834_ & ~_0070_;
	assign _1836_ = io_in[3] & ~_0070_;
	assign _1837_ = ~(_1836_ | _1835_);
	assign _0064_ = _1837_ & ~_0103_;
	assign _1838_ = ~(\mchip.focus_col [0] & \mchip.focus_col [1]);
	assign _1839_ = \mchip.focus_col [2] & ~_1838_;
	assign _0065_ = _1839_ & _0103_;
	assign _1840_ = \mchip.fsm_state  | ~\mchip.row_sel[6].col_sel[0].tile_state.state ;
	assign _0206_ = \mchip.lock_state  & ~_1840_;
	assign _1841_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[6].col_sel[0].tile_state.state_locked );
	assign _0015_ = ~(_1841_ | _0206_);
	assign _1842_ = \mchip.fsm_state  | ~\mchip.row_sel[3].col_sel[7].tile_state.state ;
	assign _0172_ = \mchip.lock_state  & ~_1842_;
	assign _1843_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[3].col_sel[7].tile_state.state_locked );
	assign _0032_ = ~(_1843_ | _0172_);
	assign _1844_ = \mchip.fsm_state  | ~\mchip.row_sel[2].col_sel[3].tile_state.state ;
	assign _0148_ = \mchip.lock_state  & ~_1844_;
	assign _1845_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[2].col_sel[3].tile_state.state_locked );
	assign _0044_ = ~(_1845_ | _0148_);
	assign _1846_ = \mchip.fsm_state  | ~\mchip.row_sel[2].col_sel[4].tile_state.state ;
	assign _0150_ = \mchip.lock_state  & ~_1846_;
	assign _1847_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[2].col_sel[4].tile_state.state_locked );
	assign _0043_ = ~(_1847_ | _0150_);
	assign _1848_ = \mchip.fsm_state  | ~\mchip.row_sel[6].col_sel[1].tile_state.state ;
	assign _0208_ = \mchip.lock_state  & ~_1848_;
	assign _1849_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[6].col_sel[1].tile_state.state_locked );
	assign _0014_ = ~(_1849_ | _0208_);
	assign _1850_ = \mchip.fsm_state  | ~\mchip.row_sel[4].col_sel[0].tile_state.state ;
	assign _0174_ = \mchip.lock_state  & ~_1850_;
	assign _1851_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[4].col_sel[0].tile_state.state_locked );
	assign _0031_ = ~(_1851_ | _0174_);
	assign _1852_ = ~(io_in[2] | io_in[3]);
	assign _1853_ = ~(_1852_ | _0103_);
	assign _0066_ = _1853_ & ~_0070_;
	assign _1854_ = \mchip.fsm_state  | ~\mchip.row_sel[6].col_sel[2].tile_state.state ;
	assign _0210_ = \mchip.lock_state  & ~_1854_;
	assign _1855_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[6].col_sel[2].tile_state.state_locked );
	assign _0013_ = ~(_1855_ | _0210_);
	assign _1856_ = \mchip.fsm_state  | ~\mchip.row_sel[6].col_sel[3].tile_state.state ;
	assign _0212_ = \mchip.lock_state  & ~_1856_;
	assign _1857_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[6].col_sel[3].tile_state.state_locked );
	assign _0012_ = ~(_1857_ | _0212_);
	assign _1858_ = \mchip.fsm_state  | ~\mchip.row_sel[6].col_sel[4].tile_state.state ;
	assign _0214_ = \mchip.lock_state  & ~_1858_;
	assign _1859_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[6].col_sel[4].tile_state.state_locked );
	assign _0011_ = ~(_1859_ | _0214_);
	assign _1860_ = \mchip.fsm_state  | ~\mchip.row_sel[6].col_sel[5].tile_state.state ;
	assign _0216_ = \mchip.lock_state  & ~_1860_;
	assign _1861_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[6].col_sel[5].tile_state.state_locked );
	assign _0010_ = ~(_1861_ | _0216_);
	assign _1862_ = \mchip.vga.frame_count [2] & ~\mchip.vga.frame_count [3];
	assign _1863_ = \mchip.vga.frame_count [0] | \mchip.vga.frame_count [1];
	assign _1864_ = _1862_ & ~_1863_;
	assign _1865_ = \mchip.vga.frame_count [7] | ~\mchip.vga.frame_count [6];
	assign _1866_ = \mchip.vga.frame_count [4] | ~\mchip.vga.frame_count [5];
	assign _1867_ = _1866_ | _1865_;
	assign _1868_ = _1864_ & ~_1867_;
	assign _1869_ = \mchip.vga.frame_count [14] | \mchip.vga.frame_count [15];
	assign _1870_ = \mchip.vga.frame_count [12] | \mchip.vga.frame_count [13];
	assign _1871_ = _1870_ | _1869_;
	assign _1872_ = \mchip.vga.frame_count [10] | \mchip.vga.frame_count [11];
	assign _1873_ = \mchip.vga.frame_count [8] | \mchip.vga.frame_count [9];
	assign _1874_ = _1873_ | _1872_;
	assign _1875_ = _1874_ | _1871_;
	assign _1876_ = _1868_ & ~_1875_;
	assign _1877_ = \mchip.vga.frame_count [30] | \mchip.vga.frame_count [31];
	assign _1878_ = \mchip.vga.frame_count [28] | \mchip.vga.frame_count [29];
	assign _1879_ = _1878_ | _1877_;
	assign _1880_ = \mchip.vga.frame_count [26] | \mchip.vga.frame_count [27];
	assign _1881_ = \mchip.vga.frame_count [24] | \mchip.vga.frame_count [25];
	assign _1882_ = _1881_ | _1880_;
	assign _1883_ = _1882_ | _1879_;
	assign _1884_ = \mchip.vga.frame_count [22] | \mchip.vga.frame_count [23];
	assign _1885_ = \mchip.vga.frame_count [20] | \mchip.vga.frame_count [21];
	assign _1886_ = _1885_ | _1884_;
	assign _1887_ = \mchip.vga.frame_count [18] | \mchip.vga.frame_count [19];
	assign _1888_ = \mchip.vga.frame_count [16] | \mchip.vga.frame_count [17];
	assign _1889_ = _1888_ | _1887_;
	assign _1890_ = _1889_ | _1886_;
	assign _1891_ = _1890_ | _1883_;
	assign _0238_ = _1876_ & ~_1891_;
	assign _1892_ = \mchip.vga.h_idx [0] | \mchip.vga.h_idx [1];
	assign _1893_ = \mchip.vga.h_idx [2] | ~\mchip.vga.h_idx [9];
	assign _1894_ = \mchip.vga.h_idx [8] | ~\mchip.vga.h_idx [7];
	assign _1895_ = _1894_ | _1893_;
	assign _1896_ = \mchip.vga.h_idx [4] & ~\mchip.vga.h_idx [3];
	assign _1897_ = _1746_ | ~_1896_;
	assign _1898_ = _1897_ | _1895_;
	assign _1899_ = _1898_ | _1892_;
	assign _1900_ = \mchip.vga.v_idx [8] & ~\mchip.vga.v_idx [9];
	assign _1901_ = ~_1900_;
	assign _1902_ = \mchip.vga.v_idx [5] & ~\mchip.vga.v_idx [4];
	assign _1903_ = \mchip.vga.v_idx [6] & \mchip.vga.v_idx [7];
	assign _1904_ = _1903_ & _1902_;
	assign _1905_ = \mchip.vga.v_idx [3] & ~\mchip.vga.v_idx [2];
	assign _1906_ = \mchip.vga.v_idx [0] | ~\mchip.vga.v_idx [1];
	assign _1907_ = _1905_ & ~_1906_;
	assign _1908_ = ~(_1907_ & _1904_);
	assign _1909_ = _1908_ | _1901_;
	assign _1910_ = _1909_ | _1899_;
	assign _1911_ = _0238_ | io_in[13];
	assign _0067_ = _1911_ | _1910_;
	assign _1912_ = _1750_ & ~_1759_;
	assign _1913_ = _1912_ | io_in[13];
	assign _0068_ = _1913_ | _1759_;
	assign _0069_ = _1910_ | io_in[13];
	assign _1914_ = \mchip.fsm_state  | ~\mchip.row_sel[7].col_sel[7].tile_state.state ;
	assign _0236_ = \mchip.lock_state  & ~_1914_;
	assign _1915_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[7].col_sel[7].tile_state.state_locked );
	assign _0000_ = ~(_1915_ | _0236_);
	assign _1916_ = \mchip.fsm_state  | ~\mchip.row_sel[7].col_sel[6].tile_state.state ;
	assign _0234_ = \mchip.lock_state  & ~_1916_;
	assign _1917_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[7].col_sel[6].tile_state.state_locked );
	assign _0001_ = ~(_1917_ | _0234_);
	assign _1918_ = \mchip.fsm_state  | ~\mchip.row_sel[7].col_sel[5].tile_state.state ;
	assign _0232_ = \mchip.lock_state  & ~_1918_;
	assign _1919_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[7].col_sel[5].tile_state.state_locked );
	assign _0002_ = ~(_1919_ | _0232_);
	assign _1920_ = \mchip.fsm_state  | ~\mchip.row_sel[7].col_sel[4].tile_state.state ;
	assign _0230_ = \mchip.lock_state  & ~_1920_;
	assign _1921_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[7].col_sel[4].tile_state.state_locked );
	assign _0003_ = ~(_1921_ | _0230_);
	assign _1922_ = \mchip.fsm_state  | ~\mchip.row_sel[7].col_sel[3].tile_state.state ;
	assign _0228_ = \mchip.lock_state  & ~_1922_;
	assign _1923_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[7].col_sel[3].tile_state.state_locked );
	assign _0004_ = ~(_1923_ | _0228_);
	assign _1924_ = \mchip.fsm_state  | ~\mchip.row_sel[7].col_sel[2].tile_state.state ;
	assign _0226_ = \mchip.lock_state  & ~_1924_;
	assign _1925_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[7].col_sel[2].tile_state.state_locked );
	assign _0005_ = ~(_1925_ | _0226_);
	assign _1926_ = \mchip.fsm_state  | ~\mchip.row_sel[7].col_sel[1].tile_state.state ;
	assign _0224_ = \mchip.lock_state  & ~_1926_;
	assign _1927_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[7].col_sel[1].tile_state.state_locked );
	assign _0006_ = ~(_1927_ | _0224_);
	assign _1928_ = \mchip.fsm_state  | ~\mchip.row_sel[7].col_sel[0].tile_state.state ;
	assign _0222_ = \mchip.lock_state  & ~_1928_;
	assign _1929_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[7].col_sel[0].tile_state.state_locked );
	assign _0007_ = ~(_1929_ | _0222_);
	assign _1930_ = \mchip.fsm_state  | ~\mchip.row_sel[6].col_sel[7].tile_state.state ;
	assign _0220_ = \mchip.lock_state  & ~_1930_;
	assign _1931_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[6].col_sel[7].tile_state.state_locked );
	assign _0008_ = ~(_1931_ | _0220_);
	assign _1932_ = \mchip.fsm_state  | ~\mchip.row_sel[6].col_sel[6].tile_state.state ;
	assign _0218_ = \mchip.lock_state  & ~_1932_;
	assign _1933_ = (\mchip.fsm_state  ? _1731_ : \mchip.row_sel[6].col_sel[6].tile_state.state_locked );
	assign _0009_ = ~(_1933_ | _0218_);
	assign _1934_ = ~\mchip.vga.frame_count [4];
	assign _1935_ = \mchip.vga.frame_count [2] | \mchip.vga.frame_count [3];
	assign _1936_ = _1935_ | _1863_;
	assign _1937_ = _1934_ & ~_1936_;
	assign _1938_ = \mchip.vga.frame_count [31] & ~_1937_;
	assign _1939_ = _1938_ | \mchip.vga.frame_count [4];
	assign _1940_ = ~(_1939_ | _1936_);
	assign _0239_ = _1940_ & ~_1938_;
	assign _1941_ = \mchip.focus_col [0] | \mchip.focus_col [1];
	assign _1942_ = \mchip.focus_col [2] & ~_1941_;
	assign _1943_ = ~\mchip.focus_row [2];
	assign _1944_ = ~(\mchip.focus_row [1] & \mchip.focus_row [0]);
	assign _1945_ = _1943_ & ~_1944_;
	assign _1946_ = _1945_ & _1942_;
	assign _1947_ = ~(\mchip.row_sel[3].col_sel[4].tile_state.state_locked  | \mchip.fsm_state );
	assign _1948_ = \mchip.row_sel[2].col_sel[4].tile_state.state  ^ \mchip.row_sel[3].col_sel[3].tile_state.state ;
	assign _1949_ = _1948_ ^ \mchip.row_sel[3].col_sel[5].tile_state.state ;
	assign _1950_ = ~(_1949_ & \mchip.row_sel[4].col_sel[4].tile_state.state );
	assign _1951_ = ~(\mchip.row_sel[2].col_sel[4].tile_state.state  & \mchip.row_sel[3].col_sel[3].tile_state.state );
	assign _1952_ = ~\mchip.row_sel[3].col_sel[5].tile_state.state ;
	assign _1953_ = _1948_ & ~_1952_;
	assign _1954_ = _1951_ & ~_1953_;
	assign _1955_ = _1954_ ^ _1950_;
	assign _1956_ = _1949_ ^ \mchip.row_sel[4].col_sel[4].tile_state.state ;
	assign _1957_ = _1956_ | _1955_;
	assign _0167_ = (_1947_ ? _1946_ : _1957_);
	assign _1958_ = \mchip.focus_row [0] | ~\mchip.focus_row [1];
	assign _1959_ = _1943_ & ~_1958_;
	assign _1960_ = _1959_ & _1839_;
	assign _1961_ = ~(\mchip.row_sel[2].col_sel[7].tile_state.state_locked  | \mchip.fsm_state );
	assign _1962_ = ~(\mchip.row_sel[1].col_sel[7].tile_state.state  ^ \mchip.row_sel[2].col_sel[6].tile_state.state );
	assign _1963_ = ~(_1962_ & \mchip.row_sel[3].col_sel[7].tile_state.state );
	assign _1964_ = ~(\mchip.row_sel[1].col_sel[7].tile_state.state  | \mchip.row_sel[2].col_sel[6].tile_state.state );
	assign _1965_ = _1964_ ^ _1963_;
	assign _1966_ = _1962_ ^ \mchip.row_sel[3].col_sel[7].tile_state.state ;
	assign _1967_ = _1966_ | _1965_;
	assign _0157_ = (_1961_ ? _1960_ : _1967_);
	assign _1968_ = \mchip.focus_col [0] | ~\mchip.focus_col [1];
	assign _1969_ = \mchip.focus_col [2] & ~_1968_;
	assign _1970_ = \mchip.focus_row [2] & ~_1958_;
	assign _1971_ = _1970_ & _1969_;
	assign _1972_ = ~(\mchip.row_sel[6].col_sel[6].tile_state.state_locked  | \mchip.fsm_state );
	assign _1973_ = \mchip.row_sel[6].col_sel[7].tile_state.state  | \mchip.row_sel[5].col_sel[6].tile_state.state ;
	assign _1974_ = ~(\mchip.row_sel[6].col_sel[7].tile_state.state  & \mchip.row_sel[5].col_sel[6].tile_state.state );
	assign _1975_ = _1974_ & _1973_;
	assign _1976_ = _1975_ ^ \mchip.row_sel[6].col_sel[5].tile_state.state ;
	assign _1977_ = ~(_1976_ & \mchip.row_sel[7].col_sel[6].tile_state.state );
	assign _1978_ = ~\mchip.row_sel[6].col_sel[5].tile_state.state ;
	assign _1979_ = _1975_ & ~_1978_;
	assign _1980_ = _1974_ & ~_1979_;
	assign _1981_ = _1980_ ^ _1977_;
	assign _1982_ = _1976_ ^ \mchip.row_sel[7].col_sel[6].tile_state.state ;
	assign _1983_ = _1982_ | _1981_;
	assign _0219_ = (_1972_ ? _1971_ : _1983_);
	assign _1984_ = \mchip.focus_row [1] | ~\mchip.focus_row [0];
	assign _1985_ = _1943_ & ~_1984_;
	assign _1986_ = _1985_ & _1839_;
	assign _1987_ = ~(\mchip.row_sel[1].col_sel[7].tile_state.state_locked  | \mchip.fsm_state );
	assign _1988_ = ~\mchip.row_sel[1].col_sel[6].tile_state.state ;
	assign _1989_ = \mchip.row_sel[1].col_sel[6].tile_state.state  | ~\mchip.row_sel[0].col_sel[7].tile_state.state ;
	assign _1990_ = ~(\mchip.row_sel[0].col_sel[7].tile_state.state  ^ \mchip.row_sel[1].col_sel[6].tile_state.state );
	assign _1991_ = _1990_ & \mchip.row_sel[2].col_sel[7].tile_state.state ;
	assign _1992_ = _1989_ & ~_1991_;
	assign _1993_ = _1992_ ^ _1988_;
	assign _1994_ = _1990_ ^ \mchip.row_sel[2].col_sel[7].tile_state.state ;
	assign _1995_ = _1994_ | _1993_;
	assign _0141_ = (_1987_ ? _1986_ : _1995_);
	assign _1996_ = _1945_ & _1839_;
	assign _1997_ = ~(\mchip.row_sel[3].col_sel[7].tile_state.state_locked  | \mchip.fsm_state );
	assign _1998_ = ~(\mchip.row_sel[4].col_sel[7].tile_state.state  ^ \mchip.row_sel[2].col_sel[7].tile_state.state );
	assign _1999_ = ~(_1998_ & \mchip.row_sel[3].col_sel[6].tile_state.state );
	assign _2000_ = ~(\mchip.row_sel[4].col_sel[7].tile_state.state  | \mchip.row_sel[2].col_sel[7].tile_state.state );
	assign _2001_ = _2000_ ^ _1999_;
	assign _2002_ = _1998_ ^ \mchip.row_sel[3].col_sel[6].tile_state.state ;
	assign _2003_ = _2002_ | _2001_;
	assign _0173_ = (_1997_ ? _1996_ : _2003_);
	assign _2004_ = ~\mchip.focus_col [2];
	assign _2005_ = _2004_ & ~_1941_;
	assign _2006_ = _2005_ & _1970_;
	assign _2007_ = ~(\mchip.row_sel[6].col_sel[0].tile_state.state_locked  | \mchip.fsm_state );
	assign _2008_ = ~\mchip.row_sel[6].col_sel[1].tile_state.state ;
	assign _2009_ = \mchip.row_sel[6].col_sel[1].tile_state.state  | ~\mchip.row_sel[5].col_sel[0].tile_state.state ;
	assign _2010_ = ~(\mchip.row_sel[6].col_sel[1].tile_state.state  ^ \mchip.row_sel[5].col_sel[0].tile_state.state );
	assign _2011_ = _2010_ & \mchip.row_sel[7].col_sel[0].tile_state.state ;
	assign _2012_ = _2009_ & ~_2011_;
	assign _2013_ = _2012_ ^ _2008_;
	assign _2014_ = _2010_ ^ \mchip.row_sel[7].col_sel[0].tile_state.state ;
	assign _2015_ = _2014_ | _2013_;
	assign _0207_ = (_2007_ ? _2006_ : _2015_);
	assign _2016_ = \mchip.focus_row [2] & ~_1984_;
	assign _2017_ = _2016_ & _1942_;
	assign _2018_ = ~(\mchip.row_sel[5].col_sel[4].tile_state.state_locked  | \mchip.fsm_state );
	assign _2019_ = \mchip.row_sel[5].col_sel[5].tile_state.state  ^ \mchip.row_sel[4].col_sel[4].tile_state.state ;
	assign _2020_ = _2019_ ^ \mchip.row_sel[5].col_sel[3].tile_state.state ;
	assign _2021_ = ~(_2020_ & \mchip.row_sel[6].col_sel[4].tile_state.state );
	assign _2022_ = ~(\mchip.row_sel[5].col_sel[5].tile_state.state  & \mchip.row_sel[4].col_sel[4].tile_state.state );
	assign _2023_ = ~\mchip.row_sel[5].col_sel[3].tile_state.state ;
	assign _2024_ = _2019_ & ~_2023_;
	assign _2025_ = _2022_ & ~_2024_;
	assign _2026_ = _2025_ ^ _2021_;
	assign _2027_ = _2020_ ^ \mchip.row_sel[6].col_sel[4].tile_state.state ;
	assign _2028_ = _2027_ | _2026_;
	assign _0199_ = (_2018_ ? _2017_ : _2028_);
	assign _2029_ = \mchip.focus_row [1] | \mchip.focus_row [0];
	assign _2030_ = \mchip.focus_row [2] & ~_2029_;
	assign _2031_ = \mchip.focus_col [1] | ~\mchip.focus_col [0];
	assign _2032_ = _2004_ & ~_2031_;
	assign _2033_ = _2032_ & _2030_;
	assign _2034_ = ~(\mchip.row_sel[4].col_sel[1].tile_state.state_locked  | \mchip.fsm_state );
	assign _2035_ = \mchip.row_sel[4].col_sel[0].tile_state.state  ^ \mchip.row_sel[4].col_sel[2].tile_state.state ;
	assign _2036_ = _2035_ ^ \mchip.row_sel[5].col_sel[1].tile_state.state ;
	assign _2037_ = ~(_2036_ & \mchip.row_sel[3].col_sel[1].tile_state.state );
	assign _2038_ = ~(\mchip.row_sel[4].col_sel[0].tile_state.state  & \mchip.row_sel[4].col_sel[2].tile_state.state );
	assign _2039_ = ~\mchip.row_sel[5].col_sel[1].tile_state.state ;
	assign _2040_ = _2035_ & ~_2039_;
	assign _2041_ = _2038_ & ~_2040_;
	assign _2042_ = _2041_ ^ _2037_;
	assign _2043_ = _2036_ ^ \mchip.row_sel[3].col_sel[1].tile_state.state ;
	assign _2044_ = _2043_ | _2042_;
	assign _0177_ = (_2034_ ? _2033_ : _2044_);
	assign _2045_ = _1985_ & _1969_;
	assign _2046_ = ~(\mchip.row_sel[1].col_sel[6].tile_state.state_locked  | \mchip.fsm_state );
	assign _2047_ = ~(\mchip.row_sel[1].col_sel[7].tile_state.state  & \mchip.row_sel[2].col_sel[6].tile_state.state );
	assign _2048_ = _2047_ & ~_1964_;
	assign _2049_ = _2048_ ^ \mchip.row_sel[0].col_sel[6].tile_state.state ;
	assign _2050_ = ~(_2049_ & \mchip.row_sel[1].col_sel[5].tile_state.state );
	assign _2051_ = _2048_ & \mchip.row_sel[0].col_sel[6].tile_state.state ;
	assign _2052_ = _2047_ & ~_2051_;
	assign _2053_ = _2052_ ^ _2050_;
	assign _2054_ = _2049_ ^ \mchip.row_sel[1].col_sel[5].tile_state.state ;
	assign _2055_ = _2054_ | _2053_;
	assign _0139_ = (_2046_ ? _2045_ : _2055_);
	assign _2056_ = _1970_ & _1839_;
	assign _2057_ = ~(\mchip.row_sel[6].col_sel[7].tile_state.state_locked  | \mchip.fsm_state );
	assign _2058_ = ~\mchip.row_sel[6].col_sel[6].tile_state.state ;
	assign _2059_ = \mchip.row_sel[6].col_sel[6].tile_state.state  | ~\mchip.row_sel[5].col_sel[7].tile_state.state ;
	assign _2060_ = ~\mchip.row_sel[7].col_sel[7].tile_state.state ;
	assign _2061_ = ~(\mchip.row_sel[6].col_sel[6].tile_state.state  ^ \mchip.row_sel[5].col_sel[7].tile_state.state );
	assign _2062_ = _2061_ & ~_2060_;
	assign _2063_ = _2059_ & ~_2062_;
	assign _2064_ = _2063_ ^ _2058_;
	assign _2065_ = _2061_ ^ \mchip.row_sel[7].col_sel[7].tile_state.state ;
	assign _2066_ = _2065_ | _2064_;
	assign _0221_ = (_2057_ ? _2056_ : _2066_);
	assign _2067_ = _1969_ & _1959_;
	assign _2068_ = ~(\mchip.row_sel[2].col_sel[6].tile_state.state_locked  | \mchip.fsm_state );
	assign _2069_ = \mchip.row_sel[1].col_sel[6].tile_state.state  ^ \mchip.row_sel[2].col_sel[7].tile_state.state ;
	assign _2070_ = _2069_ ^ \mchip.row_sel[3].col_sel[6].tile_state.state ;
	assign _2071_ = ~(_2070_ & \mchip.row_sel[2].col_sel[5].tile_state.state );
	assign _2072_ = ~(\mchip.row_sel[1].col_sel[6].tile_state.state  & \mchip.row_sel[2].col_sel[7].tile_state.state );
	assign _2073_ = _2069_ & \mchip.row_sel[3].col_sel[6].tile_state.state ;
	assign _2074_ = _2072_ & ~_2073_;
	assign _2075_ = _2074_ ^ _2071_;
	assign _2076_ = _2070_ ^ \mchip.row_sel[2].col_sel[5].tile_state.state ;
	assign _2077_ = _2076_ | _2075_;
	assign _0155_ = (_2068_ ? _2067_ : _2077_);
	assign _2078_ = _2004_ & ~_1838_;
	assign _2079_ = _2078_ & _2030_;
	assign _2080_ = ~(\mchip.row_sel[4].col_sel[3].tile_state.state_locked  | \mchip.fsm_state );
	assign _2081_ = \mchip.row_sel[3].col_sel[3].tile_state.state  ^ \mchip.row_sel[4].col_sel[2].tile_state.state ;
	assign _2082_ = _2081_ ^ \mchip.row_sel[5].col_sel[3].tile_state.state ;
	assign _2083_ = ~(_2082_ & \mchip.row_sel[4].col_sel[4].tile_state.state );
	assign _2084_ = ~(\mchip.row_sel[3].col_sel[3].tile_state.state  & \mchip.row_sel[4].col_sel[2].tile_state.state );
	assign _2085_ = _2081_ & ~_2023_;
	assign _2086_ = _2084_ & ~_2085_;
	assign _2087_ = _2086_ ^ _2083_;
	assign _2088_ = _2082_ ^ \mchip.row_sel[4].col_sel[4].tile_state.state ;
	assign _2089_ = _2088_ | _2087_;
	assign _0181_ = (_2080_ ? _2079_ : _2089_);
	assign _2090_ = _2078_ & _1945_;
	assign _2091_ = ~(\mchip.row_sel[3].col_sel[3].tile_state.state_locked  | \mchip.fsm_state );
	assign _2092_ = \mchip.row_sel[3].col_sel[4].tile_state.state  ^ \mchip.row_sel[4].col_sel[3].tile_state.state ;
	assign _2093_ = _2092_ ^ \mchip.row_sel[2].col_sel[3].tile_state.state ;
	assign _2094_ = ~(_2093_ & \mchip.row_sel[3].col_sel[2].tile_state.state );
	assign _2095_ = ~(\mchip.row_sel[3].col_sel[4].tile_state.state  & \mchip.row_sel[4].col_sel[3].tile_state.state );
	assign _2096_ = ~\mchip.row_sel[2].col_sel[3].tile_state.state ;
	assign _2097_ = _2092_ & ~_2096_;
	assign _2098_ = _2095_ & ~_2097_;
	assign _2099_ = _2098_ ^ _2094_;
	assign _2100_ = _2093_ ^ \mchip.row_sel[3].col_sel[2].tile_state.state ;
	assign _2101_ = _2100_ | _2099_;
	assign _0165_ = (_2091_ ? _2090_ : _2101_);
	assign _2102_ = \mchip.focus_col [2] & ~_2031_;
	assign _2103_ = _2102_ & _1985_;
	assign _2104_ = ~(\mchip.row_sel[1].col_sel[5].tile_state.state_locked  | \mchip.fsm_state );
	assign _2105_ = \mchip.row_sel[1].col_sel[6].tile_state.state  ^ \mchip.row_sel[2].col_sel[5].tile_state.state ;
	assign _2106_ = _2105_ ^ \mchip.row_sel[0].col_sel[5].tile_state.state ;
	assign _2107_ = ~(_2106_ & \mchip.row_sel[1].col_sel[4].tile_state.state );
	assign _2108_ = ~(\mchip.row_sel[1].col_sel[6].tile_state.state  & \mchip.row_sel[2].col_sel[5].tile_state.state );
	assign _2109_ = _2105_ & \mchip.row_sel[0].col_sel[5].tile_state.state ;
	assign _2110_ = _2108_ & ~_2109_;
	assign _2111_ = _2110_ ^ _2107_;
	assign _2112_ = _2106_ ^ \mchip.row_sel[1].col_sel[4].tile_state.state ;
	assign _2113_ = _2112_ | _2111_;
	assign _0137_ = (_2104_ ? _2103_ : _2113_);
	assign _2114_ = _2032_ & _1970_;
	assign _0253_ = ~(\mchip.row_sel[6].col_sel[1].tile_state.state_locked  | \mchip.fsm_state );
	assign _0254_ = \mchip.row_sel[7].col_sel[1].tile_state.state  ^ \mchip.row_sel[6].col_sel[0].tile_state.state ;
	assign _0255_ = _0254_ ^ \mchip.row_sel[5].col_sel[1].tile_state.state ;
	assign _0256_ = ~(_0255_ & \mchip.row_sel[6].col_sel[2].tile_state.state );
	assign _0257_ = ~(\mchip.row_sel[7].col_sel[1].tile_state.state  & \mchip.row_sel[6].col_sel[0].tile_state.state );
	assign _0258_ = _0254_ & ~_2039_;
	assign _0259_ = _0257_ & ~_0258_;
	assign _0260_ = _0259_ ^ _0256_;
	assign _0261_ = _0255_ ^ \mchip.row_sel[6].col_sel[2].tile_state.state ;
	assign _0262_ = _0261_ | _0260_;
	assign _0209_ = (_0253_ ? _2114_ : _0262_);
	assign _0263_ = \mchip.focus_row [2] & ~_1944_;
	assign _0264_ = _0263_ & _2005_;
	assign _0265_ = \mchip.row_sel[7].col_sel[0].tile_state.state_locked  | \mchip.fsm_state ;
	assign _0223_ = (_0265_ ? _0257_ : _0264_);
	assign _0266_ = _2016_ & _2005_;
	assign _0267_ = ~(\mchip.row_sel[5].col_sel[0].tile_state.state_locked  | \mchip.fsm_state );
	assign _0268_ = ~(\mchip.row_sel[6].col_sel[0].tile_state.state  ^ \mchip.row_sel[5].col_sel[1].tile_state.state );
	assign _0269_ = ~(_0268_ & \mchip.row_sel[4].col_sel[0].tile_state.state );
	assign _0270_ = ~(\mchip.row_sel[6].col_sel[0].tile_state.state  | \mchip.row_sel[5].col_sel[1].tile_state.state );
	assign _0271_ = _0270_ ^ _0269_;
	assign _0272_ = _0268_ ^ \mchip.row_sel[4].col_sel[0].tile_state.state ;
	assign _0273_ = _0272_ | _0271_;
	assign _0191_ = (_0267_ ? _0266_ : _0273_);
	assign _0274_ = _2102_ & _1959_;
	assign _0275_ = ~(\mchip.row_sel[2].col_sel[5].tile_state.state_locked  | \mchip.fsm_state );
	assign _0276_ = \mchip.row_sel[2].col_sel[6].tile_state.state  ^ \mchip.row_sel[1].col_sel[5].tile_state.state ;
	assign _0277_ = _0276_ ^ \mchip.row_sel[3].col_sel[5].tile_state.state ;
	assign _0278_ = ~(_0277_ & \mchip.row_sel[2].col_sel[4].tile_state.state );
	assign _0279_ = ~(\mchip.row_sel[2].col_sel[6].tile_state.state  & \mchip.row_sel[1].col_sel[5].tile_state.state );
	assign _0280_ = _0276_ & ~_1952_;
	assign _0281_ = _0279_ & ~_0280_;
	assign _0282_ = _0281_ ^ _0278_;
	assign _0283_ = _0277_ ^ \mchip.row_sel[2].col_sel[4].tile_state.state ;
	assign _0284_ = _0283_ | _0282_;
	assign _0153_ = (_0275_ ? _0274_ : _0284_);
	assign _0285_ = _1985_ & _1942_;
	assign _0286_ = ~(\mchip.row_sel[1].col_sel[4].tile_state.state_locked  | \mchip.fsm_state );
	assign _0287_ = \mchip.row_sel[1].col_sel[3].tile_state.state  ^ \mchip.row_sel[1].col_sel[5].tile_state.state ;
	assign _0288_ = _0287_ ^ \mchip.row_sel[0].col_sel[4].tile_state.state ;
	assign _0289_ = ~(_0288_ & \mchip.row_sel[2].col_sel[4].tile_state.state );
	assign _0290_ = ~(\mchip.row_sel[1].col_sel[3].tile_state.state  & \mchip.row_sel[1].col_sel[5].tile_state.state );
	assign _0291_ = _0287_ & \mchip.row_sel[0].col_sel[4].tile_state.state ;
	assign _0292_ = _0290_ & ~_0291_;
	assign _0293_ = _0292_ ^ _0289_;
	assign _0294_ = _0288_ ^ \mchip.row_sel[2].col_sel[4].tile_state.state ;
	assign _0295_ = _0294_ | _0293_;
	assign _0135_ = (_0286_ ? _0285_ : _0295_);
	assign _0296_ = _1968_ | \mchip.focus_col [2];
	assign _0297_ = _2016_ & ~_0296_;
	assign _0298_ = ~(\mchip.row_sel[5].col_sel[2].tile_state.state_locked  | \mchip.fsm_state );
	assign _0299_ = \mchip.row_sel[6].col_sel[2].tile_state.state  ^ \mchip.row_sel[4].col_sel[2].tile_state.state ;
	assign _0300_ = _0299_ ^ \mchip.row_sel[5].col_sel[1].tile_state.state ;
	assign _0301_ = ~(_0300_ & \mchip.row_sel[5].col_sel[3].tile_state.state );
	assign _0302_ = ~(\mchip.row_sel[6].col_sel[2].tile_state.state  & \mchip.row_sel[4].col_sel[2].tile_state.state );
	assign _0303_ = _0299_ & ~_2039_;
	assign _0304_ = _0302_ & ~_0303_;
	assign _0305_ = _0304_ ^ _0301_;
	assign _0306_ = _0300_ ^ \mchip.row_sel[5].col_sel[3].tile_state.state ;
	assign _0307_ = _0306_ | _0305_;
	assign _0195_ = (_0298_ ? _0297_ : _0307_);
	assign _0308_ = _2102_ & _2016_;
	assign _0309_ = ~(\mchip.row_sel[5].col_sel[5].tile_state.state_locked  | \mchip.fsm_state );
	assign _0310_ = \mchip.row_sel[5].col_sel[6].tile_state.state  ^ \mchip.row_sel[5].col_sel[4].tile_state.state ;
	assign _0311_ = _0310_ ^ \mchip.row_sel[6].col_sel[5].tile_state.state ;
	assign _0312_ = ~(_0311_ & \mchip.row_sel[4].col_sel[5].tile_state.state );
	assign _0313_ = ~(\mchip.row_sel[5].col_sel[6].tile_state.state  & \mchip.row_sel[5].col_sel[4].tile_state.state );
	assign _0314_ = _0310_ & ~_1978_;
	assign _0315_ = _0313_ & ~_0314_;
	assign _0316_ = _0315_ ^ _0312_;
	assign _0317_ = _0311_ ^ \mchip.row_sel[4].col_sel[5].tile_state.state ;
	assign _0318_ = _0317_ | _0316_;
	assign _0201_ = (_0309_ ? _0308_ : _0318_);
	assign _0319_ = _0263_ & _2032_;
	assign _0320_ = ~(\mchip.row_sel[7].col_sel[1].tile_state.state_locked  | \mchip.fsm_state );
	assign _0321_ = \mchip.row_sel[6].col_sel[1].tile_state.state  | ~\mchip.row_sel[7].col_sel[0].tile_state.state ;
	assign _0322_ = ~(\mchip.row_sel[7].col_sel[0].tile_state.state  ^ \mchip.row_sel[6].col_sel[1].tile_state.state );
	assign _0323_ = _0322_ & \mchip.row_sel[7].col_sel[2].tile_state.state ;
	assign _0324_ = _0321_ & ~_0323_;
	assign _0325_ = _0324_ ^ _2008_;
	assign _0326_ = _0322_ ^ \mchip.row_sel[7].col_sel[2].tile_state.state ;
	assign _0327_ = _0326_ | _0325_;
	assign _0225_ = (_0320_ ? _0319_ : _0327_);
	assign _0328_ = _1969_ & _1945_;
	assign _0329_ = ~(\mchip.row_sel[3].col_sel[6].tile_state.state_locked  | \mchip.fsm_state );
	assign _0330_ = \mchip.row_sel[3].col_sel[7].tile_state.state  ^ \mchip.row_sel[2].col_sel[6].tile_state.state ;
	assign _0331_ = _0330_ ^ \mchip.row_sel[4].col_sel[6].tile_state.state ;
	assign _0332_ = ~(_0331_ & \mchip.row_sel[3].col_sel[5].tile_state.state );
	assign _0333_ = ~(\mchip.row_sel[3].col_sel[7].tile_state.state  & \mchip.row_sel[2].col_sel[6].tile_state.state );
	assign _0334_ = ~\mchip.row_sel[4].col_sel[6].tile_state.state ;
	assign _0335_ = _0330_ & ~_0334_;
	assign _0336_ = _0333_ & ~_0335_;
	assign _0337_ = _0336_ ^ _0332_;
	assign _0338_ = _0331_ ^ \mchip.row_sel[3].col_sel[5].tile_state.state ;
	assign _0339_ = _0338_ | _0337_;
	assign _0171_ = (_0329_ ? _0328_ : _0339_);
	assign _0340_ = _2078_ & _1985_;
	assign _0341_ = ~(\mchip.row_sel[1].col_sel[3].tile_state.state_locked  | \mchip.fsm_state );
	assign _0342_ = \mchip.row_sel[1].col_sel[4].tile_state.state  ^ \mchip.row_sel[1].col_sel[2].tile_state.state ;
	assign _0343_ = _0342_ ^ \mchip.row_sel[0].col_sel[3].tile_state.state ;
	assign _0344_ = ~(_0343_ & \mchip.row_sel[2].col_sel[3].tile_state.state );
	assign _0345_ = ~(\mchip.row_sel[1].col_sel[4].tile_state.state  & \mchip.row_sel[1].col_sel[2].tile_state.state );
	assign _0346_ = _0342_ & \mchip.row_sel[0].col_sel[3].tile_state.state ;
	assign _0347_ = _0345_ & ~_0346_;
	assign _0348_ = _0347_ ^ _0344_;
	assign _0349_ = _0343_ ^ \mchip.row_sel[2].col_sel[3].tile_state.state ;
	assign _0350_ = _0349_ | _0348_;
	assign _0133_ = (_0341_ ? _0340_ : _0350_);
	assign _0351_ = _1970_ & ~_0296_;
	assign _0352_ = ~(\mchip.row_sel[6].col_sel[2].tile_state.state_locked  | \mchip.fsm_state );
	assign _0353_ = \mchip.row_sel[6].col_sel[1].tile_state.state  ^ \mchip.row_sel[5].col_sel[2].tile_state.state ;
	assign _0354_ = _0353_ ^ \mchip.row_sel[6].col_sel[3].tile_state.state ;
	assign _0355_ = ~(_0354_ & \mchip.row_sel[7].col_sel[2].tile_state.state );
	assign _0356_ = ~(\mchip.row_sel[6].col_sel[1].tile_state.state  & \mchip.row_sel[5].col_sel[2].tile_state.state );
	assign _0357_ = ~\mchip.row_sel[6].col_sel[3].tile_state.state ;
	assign _0358_ = _0353_ & ~_0357_;
	assign _0359_ = _0356_ & ~_0358_;
	assign _0360_ = _0359_ ^ _0355_;
	assign _0361_ = _0354_ ^ \mchip.row_sel[7].col_sel[2].tile_state.state ;
	assign _0362_ = _0361_ | _0360_;
	assign _0211_ = (_0352_ ? _0351_ : _0362_);
	assign _0363_ = _1959_ & _1942_;
	assign _0364_ = ~(\mchip.row_sel[2].col_sel[4].tile_state.state_locked  | \mchip.fsm_state );
	assign _0365_ = \mchip.row_sel[3].col_sel[4].tile_state.state  ^ \mchip.row_sel[2].col_sel[5].tile_state.state ;
	assign _0366_ = _0365_ ^ \mchip.row_sel[2].col_sel[3].tile_state.state ;
	assign _0367_ = ~(_0366_ & \mchip.row_sel[1].col_sel[4].tile_state.state );
	assign _0368_ = ~(\mchip.row_sel[3].col_sel[4].tile_state.state  & \mchip.row_sel[2].col_sel[5].tile_state.state );
	assign _0369_ = _0365_ & ~_2096_;
	assign _0370_ = _0368_ & ~_0369_;
	assign _0371_ = _0370_ ^ _0367_;
	assign _0372_ = _0366_ ^ \mchip.row_sel[1].col_sel[4].tile_state.state ;
	assign _0373_ = _0372_ | _0371_;
	assign _0151_ = (_0364_ ? _0363_ : _0373_);
	assign _0374_ = _1945_ & ~_0296_;
	assign _0375_ = ~(\mchip.row_sel[3].col_sel[2].tile_state.state_locked  | \mchip.fsm_state );
	assign _0376_ = _2081_ ^ \mchip.row_sel[2].col_sel[2].tile_state.state ;
	assign _0377_ = ~(_0376_ & \mchip.row_sel[3].col_sel[1].tile_state.state );
	assign _0378_ = ~\mchip.row_sel[2].col_sel[2].tile_state.state ;
	assign _0379_ = _2081_ & ~_0378_;
	assign _0380_ = _2084_ & ~_0379_;
	assign _0381_ = _0380_ ^ _0377_;
	assign _0382_ = _0376_ ^ \mchip.row_sel[3].col_sel[1].tile_state.state ;
	assign _0383_ = _0382_ | _0381_;
	assign _0163_ = (_0375_ ? _0374_ : _0383_);
	assign _0384_ = _0263_ & ~_0296_;
	assign _0385_ = ~(\mchip.row_sel[7].col_sel[2].tile_state.state_locked  | \mchip.fsm_state );
	assign _0386_ = ~(\mchip.row_sel[7].col_sel[1].tile_state.state  ^ \mchip.row_sel[7].col_sel[3].tile_state.state );
	assign _0387_ = ~(_0386_ & \mchip.row_sel[6].col_sel[2].tile_state.state );
	assign _0388_ = ~(\mchip.row_sel[7].col_sel[1].tile_state.state  | \mchip.row_sel[7].col_sel[3].tile_state.state );
	assign _0389_ = _0388_ ^ _0387_;
	assign _0390_ = _0386_ ^ \mchip.row_sel[6].col_sel[2].tile_state.state ;
	assign _0391_ = _0390_ | _0389_;
	assign _0227_ = (_0385_ ? _0384_ : _0391_);
	assign _0392_ = _1985_ & ~_0296_;
	assign _0393_ = ~(\mchip.row_sel[1].col_sel[2].tile_state.state_locked  | \mchip.fsm_state );
	assign _0394_ = \mchip.row_sel[1].col_sel[3].tile_state.state  ^ \mchip.row_sel[1].col_sel[1].tile_state.state ;
	assign _0395_ = _0394_ ^ \mchip.row_sel[0].col_sel[2].tile_state.state ;
	assign _0396_ = ~(_0395_ & \mchip.row_sel[2].col_sel[2].tile_state.state );
	assign _0397_ = ~(\mchip.row_sel[1].col_sel[3].tile_state.state  & \mchip.row_sel[1].col_sel[1].tile_state.state );
	assign _0398_ = ~\mchip.row_sel[0].col_sel[2].tile_state.state ;
	assign _0399_ = _0394_ & ~_0398_;
	assign _0400_ = _0397_ & ~_0399_;
	assign _0401_ = _0400_ ^ _0396_;
	assign _0402_ = _0395_ ^ \mchip.row_sel[2].col_sel[2].tile_state.state ;
	assign _0403_ = _0402_ | _0401_;
	assign _0131_ = (_0393_ ? _0392_ : _0403_);
	assign _0404_ = _2030_ & ~_0296_;
	assign _0405_ = ~(\mchip.row_sel[4].col_sel[2].tile_state.state_locked  | \mchip.fsm_state );
	assign _0406_ = \mchip.row_sel[4].col_sel[3].tile_state.state  ^ \mchip.row_sel[4].col_sel[1].tile_state.state ;
	assign _0407_ = _0406_ ^ \mchip.row_sel[3].col_sel[2].tile_state.state ;
	assign _0408_ = ~(_0407_ & \mchip.row_sel[5].col_sel[2].tile_state.state );
	assign _0409_ = ~(\mchip.row_sel[4].col_sel[3].tile_state.state  & \mchip.row_sel[4].col_sel[1].tile_state.state );
	assign _0410_ = _0406_ & \mchip.row_sel[3].col_sel[2].tile_state.state ;
	assign _0411_ = _0409_ & ~_0410_;
	assign _0412_ = _0411_ ^ _0408_;
	assign _0413_ = _0407_ ^ \mchip.row_sel[5].col_sel[2].tile_state.state ;
	assign _0414_ = _0413_ | _0412_;
	assign _0179_ = (_0405_ ? _0404_ : _0414_);
	assign _0415_ = _2030_ & _1839_;
	assign _0416_ = ~(\mchip.row_sel[4].col_sel[7].tile_state.state_locked  | \mchip.fsm_state );
	assign _0417_ = ~(\mchip.row_sel[3].col_sel[7].tile_state.state  ^ \mchip.row_sel[4].col_sel[6].tile_state.state );
	assign _0418_ = ~(_0417_ & \mchip.row_sel[5].col_sel[7].tile_state.state );
	assign _0419_ = ~(\mchip.row_sel[3].col_sel[7].tile_state.state  | \mchip.row_sel[4].col_sel[6].tile_state.state );
	assign _0420_ = _0419_ ^ _0418_;
	assign _0421_ = _0417_ ^ \mchip.row_sel[5].col_sel[7].tile_state.state ;
	assign _0422_ = _0421_ | _0420_;
	assign _0189_ = (_0416_ ? _0415_ : _0422_);
	assign _0423_ = _2030_ & _2005_;
	assign _0424_ = ~(\mchip.row_sel[4].col_sel[0].tile_state.state_locked  | \mchip.fsm_state );
	assign _0425_ = ~(\mchip.row_sel[3].col_sel[0].tile_state.state  ^ \mchip.row_sel[4].col_sel[1].tile_state.state );
	assign _0426_ = ~(_0425_ & \mchip.row_sel[5].col_sel[0].tile_state.state );
	assign _0427_ = ~(\mchip.row_sel[3].col_sel[0].tile_state.state  | \mchip.row_sel[4].col_sel[1].tile_state.state );
	assign _0428_ = _0427_ ^ _0426_;
	assign _0429_ = _0425_ ^ \mchip.row_sel[5].col_sel[0].tile_state.state ;
	assign _0430_ = _0429_ | _0428_;
	assign _0175_ = (_0424_ ? _0423_ : _0430_);
	assign _0431_ = _2078_ & _1959_;
	assign _0432_ = ~(\mchip.row_sel[2].col_sel[3].tile_state.state_locked  | \mchip.fsm_state );
	assign _0433_ = \mchip.row_sel[1].col_sel[3].tile_state.state  ^ \mchip.row_sel[3].col_sel[3].tile_state.state ;
	assign _0434_ = _0433_ ^ \mchip.row_sel[2].col_sel[2].tile_state.state ;
	assign _0435_ = ~(_0434_ & \mchip.row_sel[2].col_sel[4].tile_state.state );
	assign _0436_ = ~(\mchip.row_sel[1].col_sel[3].tile_state.state  & \mchip.row_sel[3].col_sel[3].tile_state.state );
	assign _0437_ = _0433_ & ~_0378_;
	assign _0438_ = _0436_ & ~_0437_;
	assign _0439_ = _0438_ ^ _0435_;
	assign _0440_ = _0434_ ^ \mchip.row_sel[2].col_sel[4].tile_state.state ;
	assign _0441_ = _0440_ | _0439_;
	assign _0149_ = (_0432_ ? _0431_ : _0441_);
	assign _0442_ = _2032_ & _1985_;
	assign _0443_ = ~(\mchip.row_sel[1].col_sel[1].tile_state.state_locked  | \mchip.fsm_state );
	assign _0444_ = \mchip.row_sel[1].col_sel[2].tile_state.state  ^ \mchip.row_sel[1].col_sel[0].tile_state.state ;
	assign _0445_ = _0444_ ^ \mchip.row_sel[0].col_sel[1].tile_state.state ;
	assign _0446_ = ~(_0445_ & \mchip.row_sel[2].col_sel[1].tile_state.state );
	assign _0447_ = ~(\mchip.row_sel[1].col_sel[2].tile_state.state  & \mchip.row_sel[1].col_sel[0].tile_state.state );
	assign _0448_ = _0444_ & \mchip.row_sel[0].col_sel[1].tile_state.state ;
	assign _0449_ = _0447_ & ~_0448_;
	assign _0450_ = _0449_ ^ _0446_;
	assign _0451_ = _0445_ ^ \mchip.row_sel[2].col_sel[1].tile_state.state ;
	assign _0452_ = _0451_ | _0450_;
	assign _0129_ = (_0443_ ? _0442_ : _0452_);
	assign _0453_ = _0263_ & _2078_;
	assign _0454_ = ~(\mchip.row_sel[7].col_sel[3].tile_state.state_locked  | \mchip.fsm_state );
	assign _0455_ = ~(\mchip.row_sel[7].col_sel[2].tile_state.state  ^ \mchip.row_sel[7].col_sel[4].tile_state.state );
	assign _0456_ = ~(_0455_ & \mchip.row_sel[6].col_sel[3].tile_state.state );
	assign _0457_ = ~(\mchip.row_sel[7].col_sel[2].tile_state.state  | \mchip.row_sel[7].col_sel[4].tile_state.state );
	assign _0458_ = _0457_ ^ _0456_;
	assign _0459_ = _0455_ ^ \mchip.row_sel[6].col_sel[3].tile_state.state ;
	assign _0460_ = _0459_ | _0458_;
	assign _0229_ = (_0454_ ? _0453_ : _0460_);
	assign _0461_ = _2078_ & _1970_;
	assign _0462_ = ~(\mchip.row_sel[6].col_sel[3].tile_state.state_locked  | \mchip.fsm_state );
	assign _0463_ = \mchip.row_sel[7].col_sel[3].tile_state.state  ^ \mchip.row_sel[6].col_sel[2].tile_state.state ;
	assign _0464_ = _0463_ ^ \mchip.row_sel[5].col_sel[3].tile_state.state ;
	assign _0465_ = ~(_0464_ & \mchip.row_sel[6].col_sel[4].tile_state.state );
	assign _0466_ = ~(\mchip.row_sel[7].col_sel[3].tile_state.state  & \mchip.row_sel[6].col_sel[2].tile_state.state );
	assign _0467_ = _0463_ & ~_2023_;
	assign _0468_ = _0466_ & ~_0467_;
	assign _0469_ = _0468_ ^ _0465_;
	assign _0470_ = _0464_ ^ \mchip.row_sel[6].col_sel[4].tile_state.state ;
	assign _0471_ = _0470_ | _0469_;
	assign _0213_ = (_0462_ ? _0461_ : _0471_);
	assign _0472_ = _2016_ & _1969_;
	assign _0473_ = ~(\mchip.row_sel[5].col_sel[6].tile_state.state_locked  | \mchip.fsm_state );
	assign _0474_ = \mchip.row_sel[6].col_sel[6].tile_state.state  ^ \mchip.row_sel[5].col_sel[5].tile_state.state ;
	assign _0475_ = _0474_ ^ \mchip.row_sel[4].col_sel[6].tile_state.state ;
	assign _0476_ = ~(_0475_ & \mchip.row_sel[5].col_sel[7].tile_state.state );
	assign _0477_ = ~(\mchip.row_sel[6].col_sel[6].tile_state.state  & \mchip.row_sel[5].col_sel[5].tile_state.state );
	assign _0478_ = _0474_ & ~_0334_;
	assign _0479_ = _0477_ & ~_0478_;
	assign _0480_ = _0479_ ^ _0476_;
	assign _0481_ = _0475_ ^ \mchip.row_sel[5].col_sel[7].tile_state.state ;
	assign _0482_ = _0481_ | _0480_;
	assign _0203_ = (_0473_ ? _0472_ : _0482_);
	assign _0483_ = _2032_ & _1945_;
	assign _0484_ = ~(\mchip.row_sel[3].col_sel[1].tile_state.state_locked  | \mchip.fsm_state );
	assign _0485_ = \mchip.row_sel[3].col_sel[2].tile_state.state  ^ \mchip.row_sel[4].col_sel[1].tile_state.state ;
	assign _0486_ = _0485_ ^ \mchip.row_sel[3].col_sel[0].tile_state.state ;
	assign _0487_ = ~(_0486_ & \mchip.row_sel[2].col_sel[1].tile_state.state );
	assign _0488_ = ~(\mchip.row_sel[3].col_sel[2].tile_state.state  & \mchip.row_sel[4].col_sel[1].tile_state.state );
	assign _0489_ = _0485_ & \mchip.row_sel[3].col_sel[0].tile_state.state ;
	assign _0490_ = _0488_ & ~_0489_;
	assign _0491_ = _0490_ ^ _0487_;
	assign _0492_ = _0486_ ^ \mchip.row_sel[2].col_sel[1].tile_state.state ;
	assign _0493_ = _0492_ | _0491_;
	assign _0161_ = (_0484_ ? _0483_ : _0493_);
	assign _0494_ = _2005_ & _1985_;
	assign _0495_ = ~(\mchip.row_sel[1].col_sel[0].tile_state.state_locked  | \mchip.fsm_state );
	assign _0496_ = ~\mchip.row_sel[1].col_sel[1].tile_state.state ;
	assign _0497_ = \mchip.row_sel[1].col_sel[1].tile_state.state  | ~\mchip.row_sel[0].col_sel[0].tile_state.state ;
	assign _0498_ = ~\mchip.row_sel[2].col_sel[0].tile_state.state ;
	assign _0499_ = ~(\mchip.row_sel[0].col_sel[0].tile_state.state  ^ \mchip.row_sel[1].col_sel[1].tile_state.state );
	assign _0500_ = _0499_ & ~_0498_;
	assign _0501_ = _0497_ & ~_0500_;
	assign _0502_ = _0501_ ^ _0496_;
	assign _0503_ = _0499_ ^ \mchip.row_sel[2].col_sel[0].tile_state.state ;
	assign _0504_ = _0503_ | _0502_;
	assign _0127_ = (_0495_ ? _0494_ : _0504_);
	assign _0505_ = _2030_ & _1942_;
	assign _0506_ = ~(\mchip.row_sel[4].col_sel[4].tile_state.state_locked  | \mchip.fsm_state );
	assign _0507_ = \mchip.row_sel[5].col_sel[4].tile_state.state  ^ \mchip.row_sel[3].col_sel[4].tile_state.state ;
	assign _0508_ = _0507_ ^ \mchip.row_sel[4].col_sel[5].tile_state.state ;
	assign _0509_ = ~(_0508_ & \mchip.row_sel[4].col_sel[3].tile_state.state );
	assign _0510_ = ~(\mchip.row_sel[5].col_sel[4].tile_state.state  & \mchip.row_sel[3].col_sel[4].tile_state.state );
	assign _0511_ = ~\mchip.row_sel[4].col_sel[5].tile_state.state ;
	assign _0512_ = _0507_ & ~_0511_;
	assign _0513_ = _0510_ & ~_0512_;
	assign _0514_ = _0513_ ^ _0509_;
	assign _0515_ = _0508_ ^ \mchip.row_sel[4].col_sel[3].tile_state.state ;
	assign _0516_ = _0515_ | _0514_;
	assign _0183_ = (_0506_ ? _0505_ : _0516_);
	assign _0517_ = _0263_ & _1942_;
	assign _0518_ = ~(\mchip.row_sel[7].col_sel[4].tile_state.state_locked  | \mchip.fsm_state );
	assign _0519_ = ~(\mchip.row_sel[7].col_sel[3].tile_state.state  ^ \mchip.row_sel[7].col_sel[5].tile_state.state );
	assign _0520_ = ~(_0519_ & \mchip.row_sel[6].col_sel[4].tile_state.state );
	assign _0521_ = ~(\mchip.row_sel[7].col_sel[3].tile_state.state  | \mchip.row_sel[7].col_sel[5].tile_state.state );
	assign _0522_ = _0521_ ^ _0520_;
	assign _0523_ = _0519_ ^ \mchip.row_sel[6].col_sel[4].tile_state.state ;
	assign _0524_ = _0523_ | _0522_;
	assign _0231_ = (_0518_ ? _0517_ : _0524_);
	assign _0525_ = _1959_ & ~_0296_;
	assign _0526_ = ~(\mchip.row_sel[2].col_sel[2].tile_state.state_locked  | \mchip.fsm_state );
	assign _0527_ = \mchip.row_sel[3].col_sel[2].tile_state.state  ^ \mchip.row_sel[1].col_sel[2].tile_state.state ;
	assign _0528_ = _0527_ ^ \mchip.row_sel[2].col_sel[1].tile_state.state ;
	assign _0529_ = ~(_0528_ & \mchip.row_sel[2].col_sel[3].tile_state.state );
	assign _0530_ = ~(\mchip.row_sel[3].col_sel[2].tile_state.state  & \mchip.row_sel[1].col_sel[2].tile_state.state );
	assign _0531_ = _0527_ & \mchip.row_sel[2].col_sel[1].tile_state.state ;
	assign _0532_ = _0530_ & ~_0531_;
	assign _0533_ = _0532_ ^ _0529_;
	assign _0534_ = _0528_ ^ \mchip.row_sel[2].col_sel[3].tile_state.state ;
	assign _0535_ = _0534_ | _0533_;
	assign _0147_ = (_0526_ ? _0525_ : _0535_);
	assign _0536_ = _2102_ & _1945_;
	assign _0537_ = ~(\mchip.row_sel[3].col_sel[5].tile_state.state_locked  | \mchip.fsm_state );
	assign _0538_ = _0365_ ^ \mchip.row_sel[4].col_sel[5].tile_state.state ;
	assign _0539_ = ~(_0538_ & \mchip.row_sel[3].col_sel[6].tile_state.state );
	assign _0540_ = _0365_ & ~_0511_;
	assign _0541_ = _0368_ & ~_0540_;
	assign _0542_ = _0541_ ^ _0539_;
	assign _0543_ = _0538_ ^ \mchip.row_sel[3].col_sel[6].tile_state.state ;
	assign _0544_ = _0543_ | _0542_;
	assign _0169_ = (_0537_ ? _0536_ : _0544_);
	assign _0545_ = _2029_ | \mchip.focus_row [2];
	assign _0546_ = _1839_ & ~_0545_;
	assign _0547_ = ~(\mchip.row_sel[0].col_sel[7].tile_state.state_locked  | \mchip.fsm_state );
	assign _0548_ = ~(\mchip.row_sel[1].col_sel[7].tile_state.state  & \mchip.row_sel[0].col_sel[6].tile_state.state );
	assign _0125_ = (_0547_ ? _0546_ : _0548_);
	assign _0549_ = _1970_ & _1942_;
	assign _0550_ = ~(\mchip.row_sel[6].col_sel[4].tile_state.state_locked  | \mchip.fsm_state );
	assign _0551_ = \mchip.row_sel[6].col_sel[3].tile_state.state  ^ \mchip.row_sel[5].col_sel[4].tile_state.state ;
	assign _0552_ = _0551_ ^ \mchip.row_sel[6].col_sel[5].tile_state.state ;
	assign _0553_ = ~(_0552_ & \mchip.row_sel[7].col_sel[4].tile_state.state );
	assign _0554_ = ~(\mchip.row_sel[6].col_sel[3].tile_state.state  & \mchip.row_sel[5].col_sel[4].tile_state.state );
	assign _0555_ = _0551_ & ~_1978_;
	assign _0556_ = _0554_ & ~_0555_;
	assign _0557_ = _0556_ ^ _0553_;
	assign _0558_ = _0552_ ^ \mchip.row_sel[7].col_sel[4].tile_state.state ;
	assign _0559_ = _0558_ | _0557_;
	assign _0215_ = (_0550_ ? _0549_ : _0559_);
	assign _0560_ = _2078_ & _2016_;
	assign _0561_ = ~(\mchip.row_sel[5].col_sel[3].tile_state.state_locked  | \mchip.fsm_state );
	assign _0562_ = \mchip.row_sel[5].col_sel[4].tile_state.state  ^ \mchip.row_sel[4].col_sel[3].tile_state.state ;
	assign _0563_ = _0562_ ^ \mchip.row_sel[6].col_sel[3].tile_state.state ;
	assign _0564_ = ~(_0563_ & \mchip.row_sel[5].col_sel[2].tile_state.state );
	assign _0565_ = ~(\mchip.row_sel[5].col_sel[4].tile_state.state  & \mchip.row_sel[4].col_sel[3].tile_state.state );
	assign _0566_ = _0562_ & ~_0357_;
	assign _0567_ = _0565_ & ~_0566_;
	assign _0568_ = _0567_ ^ _0564_;
	assign _0569_ = _0563_ ^ \mchip.row_sel[5].col_sel[2].tile_state.state ;
	assign _0570_ = _0569_ | _0568_;
	assign _0197_ = (_0561_ ? _0560_ : _0570_);
	assign _0571_ = _0263_ & _2102_;
	assign _0572_ = ~(\mchip.row_sel[7].col_sel[5].tile_state.state_locked  | \mchip.fsm_state );
	assign _0573_ = ~(\mchip.row_sel[7].col_sel[4].tile_state.state  ^ \mchip.row_sel[6].col_sel[5].tile_state.state );
	assign _0574_ = ~(_0573_ & \mchip.row_sel[7].col_sel[6].tile_state.state );
	assign _0575_ = ~(\mchip.row_sel[7].col_sel[4].tile_state.state  | \mchip.row_sel[6].col_sel[5].tile_state.state );
	assign _0576_ = _0575_ ^ _0574_;
	assign _0577_ = _0573_ ^ \mchip.row_sel[7].col_sel[6].tile_state.state ;
	assign _0578_ = _0577_ | _0576_;
	assign _0233_ = (_0572_ ? _0571_ : _0578_);
	assign _0579_ = _2102_ & _2030_;
	assign _0580_ = ~(\mchip.row_sel[4].col_sel[5].tile_state.state_locked  | \mchip.fsm_state );
	assign _0581_ = _2019_ ^ \mchip.row_sel[4].col_sel[6].tile_state.state ;
	assign _0582_ = ~(_0581_ & \mchip.row_sel[3].col_sel[5].tile_state.state );
	assign _0583_ = _2019_ & ~_0334_;
	assign _0584_ = _2022_ & ~_0583_;
	assign _0585_ = _0584_ ^ _0582_;
	assign _0586_ = _0581_ ^ \mchip.row_sel[3].col_sel[5].tile_state.state ;
	assign _0587_ = _0586_ | _0585_;
	assign _0185_ = (_0580_ ? _0579_ : _0587_);
	assign _0588_ = _1969_ & ~_0545_;
	assign _0589_ = ~(\mchip.row_sel[0].col_sel[6].tile_state.state_locked  | \mchip.fsm_state );
	assign _0590_ = \mchip.row_sel[1].col_sel[6].tile_state.state  | ~\mchip.row_sel[0].col_sel[5].tile_state.state ;
	assign _0591_ = ~(\mchip.row_sel[1].col_sel[6].tile_state.state  ^ \mchip.row_sel[0].col_sel[5].tile_state.state );
	assign _0592_ = _0591_ & \mchip.row_sel[0].col_sel[7].tile_state.state ;
	assign _0593_ = _0590_ & ~_0592_;
	assign _0594_ = _0593_ ^ _1988_;
	assign _0595_ = _0591_ ^ \mchip.row_sel[0].col_sel[7].tile_state.state ;
	assign _0596_ = _0595_ | _0594_;
	assign _0123_ = (_0589_ ? _0588_ : _0596_);
	assign _0597_ = _2032_ & _1959_;
	assign _0598_ = ~(\mchip.row_sel[2].col_sel[1].tile_state.state_locked  | \mchip.fsm_state );
	assign _0599_ = \mchip.row_sel[1].col_sel[1].tile_state.state  ^ \mchip.row_sel[3].col_sel[1].tile_state.state ;
	assign _0600_ = _0599_ ^ \mchip.row_sel[2].col_sel[0].tile_state.state ;
	assign _0601_ = ~(_0600_ & \mchip.row_sel[2].col_sel[2].tile_state.state );
	assign _0602_ = ~(\mchip.row_sel[1].col_sel[1].tile_state.state  & \mchip.row_sel[3].col_sel[1].tile_state.state );
	assign _0603_ = _0599_ & ~_0498_;
	assign _0604_ = _0602_ & ~_0603_;
	assign _0605_ = _0604_ ^ _0601_;
	assign _0606_ = _0600_ ^ \mchip.row_sel[2].col_sel[2].tile_state.state ;
	assign _0607_ = _0606_ | _0605_;
	assign _0145_ = (_0598_ ? _0597_ : _0607_);
	assign _0608_ = _2005_ & _1945_;
	assign _0609_ = ~(\mchip.row_sel[3].col_sel[0].tile_state.state_locked  | \mchip.fsm_state );
	assign _0610_ = ~(\mchip.row_sel[4].col_sel[0].tile_state.state  ^ \mchip.row_sel[2].col_sel[0].tile_state.state );
	assign _0611_ = ~(_0610_ & \mchip.row_sel[3].col_sel[1].tile_state.state );
	assign _0612_ = ~(\mchip.row_sel[4].col_sel[0].tile_state.state  | \mchip.row_sel[2].col_sel[0].tile_state.state );
	assign _0613_ = _0612_ ^ _0611_;
	assign _0614_ = _0610_ ^ \mchip.row_sel[3].col_sel[1].tile_state.state ;
	assign _0615_ = _0614_ | _0613_;
	assign _0159_ = (_0609_ ? _0608_ : _0615_);
	assign _0616_ = _2016_ & _1839_;
	assign _0617_ = ~(\mchip.row_sel[5].col_sel[7].tile_state.state_locked  | \mchip.fsm_state );
	assign _0618_ = ~(\mchip.row_sel[6].col_sel[7].tile_state.state  ^ \mchip.row_sel[5].col_sel[6].tile_state.state );
	assign _0619_ = _0618_ & \mchip.row_sel[4].col_sel[7].tile_state.state ;
	assign _0620_ = _0619_ ^ _1973_;
	assign _0621_ = _0618_ ^ \mchip.row_sel[4].col_sel[7].tile_state.state ;
	assign _0622_ = _0621_ | _0620_;
	assign _0205_ = (_0617_ ? _0616_ : _0622_);
	assign _0623_ = _0263_ & _1969_;
	assign _0624_ = ~(\mchip.row_sel[7].col_sel[6].tile_state.state_locked  | \mchip.fsm_state );
	assign _0625_ = \mchip.row_sel[6].col_sel[6].tile_state.state  | ~\mchip.row_sel[7].col_sel[5].tile_state.state ;
	assign _0626_ = ~(\mchip.row_sel[6].col_sel[6].tile_state.state  ^ \mchip.row_sel[7].col_sel[5].tile_state.state );
	assign _0627_ = _0626_ & ~_2060_;
	assign _0628_ = _0625_ & ~_0627_;
	assign _0629_ = _0628_ ^ _2058_;
	assign _0630_ = _0626_ ^ \mchip.row_sel[7].col_sel[7].tile_state.state ;
	assign _0631_ = _0630_ | _0629_;
	assign _0235_ = (_0624_ ? _0623_ : _0631_);
	assign _0632_ = _2102_ & ~_0545_;
	assign _0633_ = ~(\mchip.row_sel[0].col_sel[5].tile_state.state_locked  | \mchip.fsm_state );
	assign _0634_ = ~(\mchip.row_sel[0].col_sel[4].tile_state.state  ^ \mchip.row_sel[1].col_sel[5].tile_state.state );
	assign _0635_ = ~(_0634_ & \mchip.row_sel[0].col_sel[6].tile_state.state );
	assign _0636_ = ~(\mchip.row_sel[0].col_sel[4].tile_state.state  | \mchip.row_sel[1].col_sel[5].tile_state.state );
	assign _0637_ = _0636_ ^ _0635_;
	assign _0638_ = _0634_ ^ \mchip.row_sel[0].col_sel[6].tile_state.state ;
	assign _0639_ = _0638_ | _0637_;
	assign _0121_ = (_0633_ ? _0632_ : _0639_);
	assign _0640_ = _2102_ & _1970_;
	assign _0641_ = ~(\mchip.row_sel[6].col_sel[5].tile_state.state_locked  | \mchip.fsm_state );
	assign _0642_ = _0474_ ^ \mchip.row_sel[7].col_sel[5].tile_state.state ;
	assign _0643_ = ~(_0642_ & \mchip.row_sel[6].col_sel[4].tile_state.state );
	assign _0644_ = _0474_ & \mchip.row_sel[7].col_sel[5].tile_state.state ;
	assign _0645_ = _0477_ & ~_0644_;
	assign _0646_ = _0645_ ^ _0643_;
	assign _0647_ = _0642_ ^ \mchip.row_sel[6].col_sel[4].tile_state.state ;
	assign _0648_ = _0647_ | _0646_;
	assign _0217_ = (_0641_ ? _0640_ : _0648_);
	assign _0649_ = _2032_ & _2016_;
	assign _0650_ = ~(\mchip.row_sel[5].col_sel[1].tile_state.state_locked  | \mchip.fsm_state );
	assign _0651_ = \mchip.row_sel[6].col_sel[1].tile_state.state  ^ \mchip.row_sel[4].col_sel[1].tile_state.state ;
	assign _0652_ = _0651_ ^ \mchip.row_sel[5].col_sel[2].tile_state.state ;
	assign _0653_ = ~(_0652_ & \mchip.row_sel[5].col_sel[0].tile_state.state );
	assign _0654_ = ~(\mchip.row_sel[6].col_sel[1].tile_state.state  & \mchip.row_sel[4].col_sel[1].tile_state.state );
	assign _0655_ = _0651_ & \mchip.row_sel[5].col_sel[2].tile_state.state ;
	assign _0656_ = _0654_ & ~_0655_;
	assign _0657_ = _0656_ ^ _0653_;
	assign _0658_ = _0652_ ^ \mchip.row_sel[5].col_sel[0].tile_state.state ;
	assign _0659_ = _0658_ | _0657_;
	assign _0193_ = (_0650_ ? _0649_ : _0659_);
	assign _0660_ = _2005_ & _1959_;
	assign _0661_ = ~(\mchip.row_sel[2].col_sel[0].tile_state.state_locked  | \mchip.fsm_state );
	assign _0662_ = ~(\mchip.row_sel[3].col_sel[0].tile_state.state  ^ \mchip.row_sel[1].col_sel[0].tile_state.state );
	assign _0663_ = ~(_0662_ & \mchip.row_sel[2].col_sel[1].tile_state.state );
	assign _0664_ = ~(\mchip.row_sel[3].col_sel[0].tile_state.state  | \mchip.row_sel[1].col_sel[0].tile_state.state );
	assign _0665_ = _0664_ ^ _0663_;
	assign _0666_ = _0662_ ^ \mchip.row_sel[2].col_sel[1].tile_state.state ;
	assign _0667_ = _0666_ | _0665_;
	assign _0143_ = (_0661_ ? _0660_ : _0667_);
	assign _0668_ = _2030_ & _1969_;
	assign _0669_ = ~(\mchip.row_sel[4].col_sel[6].tile_state.state_locked  | \mchip.fsm_state );
	assign _0670_ = \mchip.row_sel[3].col_sel[6].tile_state.state  ^ \mchip.row_sel[4].col_sel[7].tile_state.state ;
	assign _0671_ = _0670_ ^ \mchip.row_sel[4].col_sel[5].tile_state.state ;
	assign _0672_ = ~(_0671_ & \mchip.row_sel[5].col_sel[6].tile_state.state );
	assign _0673_ = ~(\mchip.row_sel[3].col_sel[6].tile_state.state  & \mchip.row_sel[4].col_sel[7].tile_state.state );
	assign _0674_ = _0670_ & ~_0511_;
	assign _0675_ = _0673_ & ~_0674_;
	assign _0676_ = _0675_ ^ _0672_;
	assign _0677_ = _0671_ ^ \mchip.row_sel[5].col_sel[6].tile_state.state ;
	assign _0678_ = _0677_ | _0676_;
	assign _0187_ = (_0669_ ? _0668_ : _0678_);
	assign _0679_ = _1942_ & ~_0545_;
	assign _0680_ = ~(\mchip.row_sel[0].col_sel[4].tile_state.state_locked  | \mchip.fsm_state );
	assign _0681_ = ~(\mchip.row_sel[1].col_sel[4].tile_state.state  ^ \mchip.row_sel[0].col_sel[3].tile_state.state );
	assign _0682_ = ~(_0681_ & \mchip.row_sel[0].col_sel[5].tile_state.state );
	assign _0683_ = ~(\mchip.row_sel[1].col_sel[4].tile_state.state  | \mchip.row_sel[0].col_sel[3].tile_state.state );
	assign _0684_ = _0683_ ^ _0682_;
	assign _0685_ = _0681_ ^ \mchip.row_sel[0].col_sel[5].tile_state.state ;
	assign _0686_ = _0685_ | _0684_;
	assign _0119_ = (_0680_ ? _0679_ : _0686_);
	assign _0687_ = ~(\mchip.row_sel[6].col_sel[7].tile_state.state  & \mchip.row_sel[7].col_sel[6].tile_state.state );
	assign _0688_ = \mchip.row_sel[7].col_sel[7].tile_state.state_locked  | \mchip.fsm_state ;
	assign _0689_ = _0263_ & _1839_;
	assign _0237_ = (_0688_ ? _0687_ : _0689_);
	assign _0690_ = _2078_ & ~_0545_;
	assign _0691_ = ~(\mchip.row_sel[0].col_sel[3].tile_state.state_locked  | \mchip.fsm_state );
	assign _0692_ = ~(\mchip.row_sel[1].col_sel[3].tile_state.state  ^ \mchip.row_sel[0].col_sel[2].tile_state.state );
	assign _0693_ = ~(_0692_ & \mchip.row_sel[0].col_sel[4].tile_state.state );
	assign _0694_ = ~(\mchip.row_sel[1].col_sel[3].tile_state.state  | \mchip.row_sel[0].col_sel[2].tile_state.state );
	assign _0695_ = _0694_ ^ _0693_;
	assign _0696_ = _0692_ ^ \mchip.row_sel[0].col_sel[4].tile_state.state ;
	assign _0697_ = _0696_ | _0695_;
	assign _0117_ = (_0691_ ? _0690_ : _0697_);
	assign _0698_ = ~(_0545_ | _0296_);
	assign _0699_ = ~(\mchip.row_sel[0].col_sel[2].tile_state.state_locked  | \mchip.fsm_state );
	assign _0700_ = ~(\mchip.row_sel[0].col_sel[1].tile_state.state  ^ \mchip.row_sel[1].col_sel[2].tile_state.state );
	assign _0701_ = ~(_0700_ & \mchip.row_sel[0].col_sel[3].tile_state.state );
	assign _0702_ = ~(\mchip.row_sel[0].col_sel[1].tile_state.state  | \mchip.row_sel[1].col_sel[2].tile_state.state );
	assign _0703_ = _0702_ ^ _0701_;
	assign _0704_ = _0700_ ^ \mchip.row_sel[0].col_sel[3].tile_state.state ;
	assign _0705_ = _0704_ | _0703_;
	assign _0115_ = (_0699_ ? _0698_ : _0705_);
	assign _0706_ = _2032_ & ~_0545_;
	assign _0707_ = ~(\mchip.row_sel[0].col_sel[1].tile_state.state_locked  | \mchip.fsm_state );
	assign _0708_ = _0499_ & ~_0398_;
	assign _0709_ = _0497_ & ~_0708_;
	assign _0710_ = _0709_ ^ _0496_;
	assign _0711_ = _0499_ ^ \mchip.row_sel[0].col_sel[2].tile_state.state ;
	assign _0712_ = _0711_ | _0710_;
	assign _0113_ = (_0707_ ? _0706_ : _0712_);
	assign _0713_ = _2005_ & ~_0545_;
	assign _0714_ = ~(\mchip.row_sel[0].col_sel[0].tile_state.state_locked  | \mchip.fsm_state );
	assign _0715_ = ~(\mchip.row_sel[0].col_sel[1].tile_state.state  & \mchip.row_sel[1].col_sel[0].tile_state.state );
	assign _0111_ = (_0714_ ? _0713_ : _0715_);
	assign _0716_ = \mchip.vga.v_idx [1] | ~\mchip.vga.v_idx [0];
	assign _0717_ = \mchip.vga.v_idx [2] & \mchip.vga.v_idx [3];
	assign _0718_ = _0716_ | ~_0717_;
	assign _0719_ = \mchip.vga.v_idx [6] | \mchip.vga.v_idx [7];
	assign _0720_ = ~(\mchip.vga.v_idx [4] | \mchip.vga.v_idx [5]);
	assign _0721_ = _0719_ | ~_0720_;
	assign _0722_ = ~(_0721_ | _0718_);
	assign _0723_ = \mchip.vga.v_idx [9] & ~\mchip.vga.v_idx [8];
	assign _0724_ = ~(_0723_ & _0722_);
	assign _0725_ = _0720_ & ~_0719_;
	assign _0726_ = ~(\mchip.vga.v_idx [1] | \mchip.vga.v_idx [0]);
	assign _0727_ = _0717_ & ~_0726_;
	assign _0728_ = _0727_ & ~_0721_;
	assign _0729_ = _0725_ & ~_0728_;
	assign _0730_ = _0723_ & ~_0729_;
	assign _0731_ = \mchip.vga.v_idx [9] & \mchip.vga.v_idx [8];
	assign _0732_ = _0731_ | _0730_;
	assign _0733_ = _0724_ & ~_0732_;
	assign _0734_ = ~(_0733_ ^ \mchip.vga.frame_count [0]);
	assign _0735_ = (_0252_ ? \mchip.vga.frame_count [0] : _0734_);
	assign _0736_ = _0735_ & ~_0238_;
	assign _0071_ = (_1910_ ? _0735_ : _0736_);
	assign _0737_ = \mchip.vga.frame_count [0] & \mchip.vga.frame_count [1];
	assign _0738_ = _1863_ & ~_0737_;
	assign _0739_ = (_0733_ ? \mchip.vga.frame_count [1] : _0738_);
	assign _0740_ = (_0252_ ? \mchip.vga.frame_count [1] : _0739_);
	assign _0741_ = _0740_ & ~_0238_;
	assign _0082_ = (_1910_ ? _0740_ : _0741_);
	assign _0742_ = _0737_ ^ \mchip.vga.frame_count [2];
	assign _0743_ = (_0733_ ? \mchip.vga.frame_count [2] : _0742_);
	assign _0744_ = (_0252_ ? \mchip.vga.frame_count [2] : _0743_);
	assign _0745_ = _0744_ & ~_0238_;
	assign _0093_ = (_1910_ ? _0744_ : _0745_);
	assign _0746_ = _0737_ & \mchip.vga.frame_count [2];
	assign _0747_ = _0746_ ^ \mchip.vga.frame_count [3];
	assign _0748_ = (_0733_ ? \mchip.vga.frame_count [3] : _0747_);
	assign _0749_ = (_0252_ ? \mchip.vga.frame_count [3] : _0748_);
	assign _0750_ = _0749_ & ~_0238_;
	assign _0096_ = (_1910_ ? _0749_ : _0750_);
	assign _0751_ = ~(\mchip.vga.frame_count [2] & \mchip.vga.frame_count [3]);
	assign _0752_ = _0737_ & ~_0751_;
	assign _0753_ = _0752_ ^ \mchip.vga.frame_count [4];
	assign _0754_ = (_0733_ ? \mchip.vga.frame_count [4] : _0753_);
	assign _0755_ = (_0252_ ? \mchip.vga.frame_count [4] : _0754_);
	assign _0756_ = _0755_ & ~_0238_;
	assign _0097_ = (_1910_ ? _0755_ : _0756_);
	assign _0757_ = _0752_ & ~_1934_;
	assign _0758_ = _0757_ ^ \mchip.vga.frame_count [5];
	assign _0759_ = (_0733_ ? \mchip.vga.frame_count [5] : _0758_);
	assign _0760_ = (_0252_ ? \mchip.vga.frame_count [5] : _0759_);
	assign _0761_ = _0760_ & ~_0238_;
	assign _0098_ = (_1910_ ? _0760_ : _0761_);
	assign _0762_ = ~(\mchip.vga.frame_count [5] & \mchip.vga.frame_count [4]);
	assign _0763_ = _0752_ & ~_0762_;
	assign _0764_ = _0763_ ^ \mchip.vga.frame_count [6];
	assign _0765_ = (_0733_ ? \mchip.vga.frame_count [6] : _0764_);
	assign _0766_ = (_0252_ ? \mchip.vga.frame_count [6] : _0765_);
	assign _0767_ = _0766_ & ~_0238_;
	assign _0099_ = (_1910_ ? _0766_ : _0767_);
	assign _0768_ = _0763_ & \mchip.vga.frame_count [6];
	assign _0769_ = _0768_ ^ \mchip.vga.frame_count [7];
	assign _0770_ = (_0733_ ? \mchip.vga.frame_count [7] : _0769_);
	assign _0771_ = (_0252_ ? \mchip.vga.frame_count [7] : _0770_);
	assign _0772_ = _0771_ & ~_0238_;
	assign _0100_ = (_1910_ ? _0771_ : _0772_);
	assign _0773_ = ~(\mchip.vga.frame_count [6] & \mchip.vga.frame_count [7]);
	assign _0774_ = _0773_ | _0762_;
	assign _0775_ = _0752_ & ~_0774_;
	assign _0776_ = _0775_ ^ \mchip.vga.frame_count [8];
	assign _0777_ = (_0733_ ? \mchip.vga.frame_count [8] : _0776_);
	assign _0778_ = (_0252_ ? \mchip.vga.frame_count [8] : _0777_);
	assign _0779_ = _0778_ & ~_0238_;
	assign _0101_ = (_1910_ ? _0778_ : _0779_);
	assign _0780_ = _0775_ & \mchip.vga.frame_count [8];
	assign _0781_ = _0780_ ^ \mchip.vga.frame_count [9];
	assign _0782_ = (_0733_ ? \mchip.vga.frame_count [9] : _0781_);
	assign _0783_ = (_0252_ ? \mchip.vga.frame_count [9] : _0782_);
	assign _0784_ = _0783_ & ~_0238_;
	assign _0102_ = (_1910_ ? _0783_ : _0784_);
	assign _0785_ = ~(\mchip.vga.frame_count [8] & \mchip.vga.frame_count [9]);
	assign _0786_ = _0775_ & ~_0785_;
	assign _0787_ = _0786_ ^ \mchip.vga.frame_count [10];
	assign _0788_ = (_0733_ ? \mchip.vga.frame_count [10] : _0787_);
	assign _0789_ = (_0252_ ? \mchip.vga.frame_count [10] : _0788_);
	assign _0790_ = _0789_ & ~_0238_;
	assign _0072_ = (_1910_ ? _0789_ : _0790_);
	assign _0791_ = _0786_ & \mchip.vga.frame_count [10];
	assign _0792_ = _0791_ ^ \mchip.vga.frame_count [11];
	assign _0793_ = (_0733_ ? \mchip.vga.frame_count [11] : _0792_);
	assign _0794_ = (_0252_ ? \mchip.vga.frame_count [11] : _0793_);
	assign _0795_ = _0794_ & ~_0238_;
	assign _0073_ = (_1910_ ? _0794_ : _0795_);
	assign _0796_ = ~(\mchip.vga.frame_count [10] & \mchip.vga.frame_count [11]);
	assign _0797_ = _0796_ | _0785_;
	assign _0798_ = _0775_ & ~_0797_;
	assign _0799_ = _0798_ ^ \mchip.vga.frame_count [12];
	assign _0800_ = (_0733_ ? \mchip.vga.frame_count [12] : _0799_);
	assign _0801_ = (_0252_ ? \mchip.vga.frame_count [12] : _0800_);
	assign _0802_ = _0801_ & ~_0238_;
	assign _0074_ = (_1910_ ? _0801_ : _0802_);
	assign _0803_ = _0798_ & \mchip.vga.frame_count [12];
	assign _0804_ = _0803_ ^ \mchip.vga.frame_count [13];
	assign _0805_ = (_0733_ ? \mchip.vga.frame_count [13] : _0804_);
	assign _0806_ = (_0252_ ? \mchip.vga.frame_count [13] : _0805_);
	assign _0807_ = _0806_ & ~_0238_;
	assign _0075_ = (_1910_ ? _0806_ : _0807_);
	assign _0808_ = ~(\mchip.vga.frame_count [12] & \mchip.vga.frame_count [13]);
	assign _0809_ = _0798_ & ~_0808_;
	assign _0810_ = _0809_ ^ \mchip.vga.frame_count [14];
	assign _0811_ = (_0733_ ? \mchip.vga.frame_count [14] : _0810_);
	assign _0812_ = (_0252_ ? \mchip.vga.frame_count [14] : _0811_);
	assign _0813_ = _0812_ & ~_0238_;
	assign _0076_ = (_1910_ ? _0812_ : _0813_);
	assign _0814_ = _0809_ & \mchip.vga.frame_count [14];
	assign _0815_ = _0814_ ^ \mchip.vga.frame_count [15];
	assign _0816_ = (_0733_ ? \mchip.vga.frame_count [15] : _0815_);
	assign _0817_ = (_0252_ ? \mchip.vga.frame_count [15] : _0816_);
	assign _0818_ = _0817_ & ~_0238_;
	assign _0077_ = (_1910_ ? _0817_ : _0818_);
	assign _0819_ = ~(\mchip.vga.frame_count [14] & \mchip.vga.frame_count [15]);
	assign _0820_ = _0819_ | _0808_;
	assign _0821_ = _0820_ | _0797_;
	assign _0822_ = _0775_ & ~_0821_;
	assign _0823_ = _0822_ ^ \mchip.vga.frame_count [16];
	assign _0824_ = (_0733_ ? \mchip.vga.frame_count [16] : _0823_);
	assign _0825_ = (_0252_ ? \mchip.vga.frame_count [16] : _0824_);
	assign _0826_ = _0825_ & ~_0238_;
	assign _0078_ = (_1910_ ? _0825_ : _0826_);
	assign _0827_ = _0822_ & \mchip.vga.frame_count [16];
	assign _0828_ = _0827_ ^ \mchip.vga.frame_count [17];
	assign _0829_ = (_0733_ ? \mchip.vga.frame_count [17] : _0828_);
	assign _0830_ = (_0252_ ? \mchip.vga.frame_count [17] : _0829_);
	assign _0831_ = _0830_ & ~_0238_;
	assign _0079_ = (_1910_ ? _0830_ : _0831_);
	assign _0832_ = ~(\mchip.vga.frame_count [16] & \mchip.vga.frame_count [17]);
	assign _0833_ = _0822_ & ~_0832_;
	assign _0834_ = _0833_ ^ \mchip.vga.frame_count [18];
	assign _0835_ = (_0733_ ? \mchip.vga.frame_count [18] : _0834_);
	assign _0836_ = (_0252_ ? \mchip.vga.frame_count [18] : _0835_);
	assign _0837_ = _0836_ & ~_0238_;
	assign _0080_ = (_1910_ ? _0836_ : _0837_);
	assign _0838_ = _0833_ & \mchip.vga.frame_count [18];
	assign _0839_ = _0838_ ^ \mchip.vga.frame_count [19];
	assign _0840_ = (_0733_ ? \mchip.vga.frame_count [19] : _0839_);
	assign _0841_ = (_0252_ ? \mchip.vga.frame_count [19] : _0840_);
	assign _0842_ = _0841_ & ~_0238_;
	assign _0081_ = (_1910_ ? _0841_ : _0842_);
	assign _0843_ = ~(\mchip.vga.frame_count [18] & \mchip.vga.frame_count [19]);
	assign _0844_ = _0843_ | _0832_;
	assign _0845_ = _0822_ & ~_0844_;
	assign _0846_ = _0845_ ^ \mchip.vga.frame_count [20];
	assign _0847_ = (_0733_ ? \mchip.vga.frame_count [20] : _0846_);
	assign _0848_ = (_0252_ ? \mchip.vga.frame_count [20] : _0847_);
	assign _0849_ = _0848_ & ~_0238_;
	assign _0083_ = (_1910_ ? _0848_ : _0849_);
	assign _0850_ = _0845_ & \mchip.vga.frame_count [20];
	assign _0851_ = _0850_ ^ \mchip.vga.frame_count [21];
	assign _0852_ = (_0733_ ? \mchip.vga.frame_count [21] : _0851_);
	assign _0853_ = (_0252_ ? \mchip.vga.frame_count [21] : _0852_);
	assign _0854_ = _0853_ & ~_0238_;
	assign _0084_ = (_1910_ ? _0853_ : _0854_);
	assign _0855_ = ~(\mchip.vga.frame_count [20] & \mchip.vga.frame_count [21]);
	assign _0856_ = _0845_ & ~_0855_;
	assign _0857_ = _0856_ ^ \mchip.vga.frame_count [22];
	assign _0858_ = (_0733_ ? \mchip.vga.frame_count [22] : _0857_);
	assign _0859_ = (_0252_ ? \mchip.vga.frame_count [22] : _0858_);
	assign _0860_ = _0859_ & ~_0238_;
	assign _0085_ = (_1910_ ? _0859_ : _0860_);
	assign _0861_ = _0856_ & \mchip.vga.frame_count [22];
	assign _0862_ = _0861_ ^ \mchip.vga.frame_count [23];
	assign _0863_ = (_0733_ ? \mchip.vga.frame_count [23] : _0862_);
	assign _0864_ = (_0252_ ? \mchip.vga.frame_count [23] : _0863_);
	assign _0865_ = _0864_ & ~_0238_;
	assign _0086_ = (_1910_ ? _0864_ : _0865_);
	assign _0866_ = ~(\mchip.vga.frame_count [22] & \mchip.vga.frame_count [23]);
	assign _0867_ = _0866_ | _0855_;
	assign _0868_ = _0867_ | _0844_;
	assign _0869_ = _0822_ & ~_0868_;
	assign _0870_ = _0869_ ^ \mchip.vga.frame_count [24];
	assign _0871_ = (_0733_ ? \mchip.vga.frame_count [24] : _0870_);
	assign _0872_ = (_0252_ ? \mchip.vga.frame_count [24] : _0871_);
	assign _0873_ = _0872_ & ~_0238_;
	assign _0087_ = (_1910_ ? _0872_ : _0873_);
	assign _0874_ = _0869_ & \mchip.vga.frame_count [24];
	assign _0875_ = _0874_ ^ \mchip.vga.frame_count [25];
	assign _0876_ = (_0733_ ? \mchip.vga.frame_count [25] : _0875_);
	assign _0877_ = (_0252_ ? \mchip.vga.frame_count [25] : _0876_);
	assign _0878_ = _0877_ & ~_0238_;
	assign _0088_ = (_1910_ ? _0877_ : _0878_);
	assign _0879_ = ~(\mchip.vga.frame_count [24] & \mchip.vga.frame_count [25]);
	assign _0880_ = _0869_ & ~_0879_;
	assign _0881_ = _0880_ ^ \mchip.vga.frame_count [26];
	assign _0882_ = (_0733_ ? \mchip.vga.frame_count [26] : _0881_);
	assign _0883_ = (_0252_ ? \mchip.vga.frame_count [26] : _0882_);
	assign _0884_ = _0883_ & ~_0238_;
	assign _0089_ = (_1910_ ? _0883_ : _0884_);
	assign _0885_ = _0880_ & \mchip.vga.frame_count [26];
	assign _0886_ = _0885_ ^ \mchip.vga.frame_count [27];
	assign _0887_ = (_0733_ ? \mchip.vga.frame_count [27] : _0886_);
	assign _0888_ = (_0252_ ? \mchip.vga.frame_count [27] : _0887_);
	assign _0889_ = _0888_ & ~_0238_;
	assign _0090_ = (_1910_ ? _0888_ : _0889_);
	assign _0890_ = ~(\mchip.vga.frame_count [26] & \mchip.vga.frame_count [27]);
	assign _0891_ = _0890_ | _0879_;
	assign _0892_ = _0869_ & ~_0891_;
	assign _0893_ = _0892_ ^ \mchip.vga.frame_count [28];
	assign _0894_ = (_0733_ ? \mchip.vga.frame_count [28] : _0893_);
	assign _0895_ = (_0252_ ? \mchip.vga.frame_count [28] : _0894_);
	assign _0896_ = _0895_ & ~_0238_;
	assign _0091_ = (_1910_ ? _0895_ : _0896_);
	assign _0897_ = _0892_ & \mchip.vga.frame_count [28];
	assign _0898_ = _0897_ ^ \mchip.vga.frame_count [29];
	assign _0899_ = (_0733_ ? \mchip.vga.frame_count [29] : _0898_);
	assign _0900_ = (_0252_ ? \mchip.vga.frame_count [29] : _0899_);
	assign _0901_ = _0900_ & ~_0238_;
	assign _0092_ = (_1910_ ? _0900_ : _0901_);
	assign _0902_ = ~(\mchip.vga.frame_count [28] & \mchip.vga.frame_count [29]);
	assign _0903_ = _0892_ & ~_0902_;
	assign _0904_ = _0903_ ^ \mchip.vga.frame_count [30];
	assign _0905_ = (_0733_ ? \mchip.vga.frame_count [30] : _0904_);
	assign _0906_ = (_0252_ ? \mchip.vga.frame_count [30] : _0905_);
	assign _0907_ = _0906_ & ~_0238_;
	assign _0094_ = (_1910_ ? _0906_ : _0907_);
	assign _0908_ = _0903_ & \mchip.vga.frame_count [30];
	assign _0909_ = _0908_ ^ \mchip.vga.frame_count [31];
	assign _0910_ = (_0733_ ? \mchip.vga.frame_count [31] : _0909_);
	assign _0911_ = (_0252_ ? \mchip.vga.frame_count [31] : _0910_);
	assign _0912_ = _0911_ & ~_0238_;
	assign _0095_ = (_1910_ ? _0911_ : _0912_);
	assign _0241_ = _0733_ & ~\mchip.vga.v_idx [0];
	assign _0913_ = _0716_ & _1906_;
	assign _0242_ = _0733_ & ~_0913_;
	assign _0914_ = \mchip.vga.v_idx [1] & \mchip.vga.v_idx [0];
	assign _0915_ = ~(_0914_ ^ \mchip.vga.v_idx [2]);
	assign _0243_ = _0733_ & ~_0915_;
	assign _0916_ = _0914_ & \mchip.vga.v_idx [2];
	assign _0917_ = ~(_0916_ ^ \mchip.vga.v_idx [3]);
	assign _0244_ = _0733_ & ~_0917_;
	assign _0918_ = ~(_0914_ & _0717_);
	assign _0919_ = _0918_ ^ \mchip.vga.v_idx [4];
	assign _0245_ = _0733_ & ~_0919_;
	assign _0920_ = ~\mchip.vga.v_idx [5];
	assign _0921_ = \mchip.vga.v_idx [4] & ~_0918_;
	assign _0922_ = _0921_ ^ _0920_;
	assign _0246_ = _0733_ & ~_0922_;
	assign _0923_ = ~\mchip.vga.v_idx [6];
	assign _0924_ = ~(\mchip.vga.v_idx [4] & \mchip.vga.v_idx [5]);
	assign _0925_ = ~(_0924_ | _0918_);
	assign _0926_ = _0925_ ^ _0923_;
	assign _0247_ = _0733_ & ~_0926_;
	assign _0927_ = ~(_0925_ & \mchip.vga.v_idx [6]);
	assign _0928_ = _0927_ ^ \mchip.vga.v_idx [7];
	assign _0248_ = _0733_ & ~_0928_;
	assign _0929_ = _1903_ & ~_0924_;
	assign _0930_ = _0929_ & ~_0918_;
	assign _0931_ = ~(_0930_ ^ \mchip.vga.v_idx [8]);
	assign _0249_ = _0733_ & ~_0931_;
	assign _0932_ = ~(_0930_ & \mchip.vga.v_idx [8]);
	assign _0933_ = _0932_ ^ \mchip.vga.v_idx [9];
	assign _0250_ = _0733_ & ~_0933_;
	assign _0104_ = ~(_1839_ | \mchip.focus_col [0]);
	assign _0105_ = \mchip.focus_col [0] ^ \mchip.focus_col [1];
	assign _0106_ = _1838_ ^ _2004_;
	assign _0107_ = ~(_0689_ | \mchip.focus_row [0]);
	assign _0108_ = ~(_1984_ & _1958_);
	assign _0934_ = _1944_ ^ _1943_;
	assign _0109_ = _0934_ & ~_0689_;
	assign _0935_ = \mchip.vga.h_idx [6] & \mchip.vga.h_idx [7];
	assign _0936_ = ~(\mchip.vga.h_idx [5] & \mchip.vga.h_idx [4]);
	assign _0937_ = _0935_ & ~_0936_;
	assign _0938_ = \mchip.vga.h_idx [9] & ~\mchip.vga.h_idx [8];
	assign _0939_ = _0938_ & _0937_;
	assign _0940_ = _0939_ | _1751_;
	assign _0941_ = \mchip.vga.h_idx [5] | \mchip.vga.h_idx [4];
	assign _0942_ = \mchip.vga.h_idx [6] | ~\mchip.vga.h_idx [7];
	assign _0943_ = _0942_ | ~_0941_;
	assign _0944_ = _0943_ & ~_0935_;
	assign _0945_ = _0938_ & ~_0944_;
	assign _0946_ = _0945_ | _1751_;
	assign _0947_ = _1899_ & ~_0946_;
	assign _0240_ = _0947_ | _0940_;
	assign _0948_ = _0726_ & _0717_;
	assign _0949_ = ~(_0948_ & _1904_);
	assign _0950_ = _1900_ & ~_0949_;
	assign _0951_ = ~(\mchip.vga.v_idx [9] | \mchip.vga.v_idx [8]);
	assign _0952_ = ~_0951_;
	assign _0953_ = _1903_ & ~_0920_;
	assign _0954_ = _0726_ | ~_0717_;
	assign _0955_ = _0954_ & _1904_;
	assign _0956_ = _0953_ & ~_0955_;
	assign _0957_ = _1900_ & ~_0956_;
	assign _0958_ = _0952_ & ~_0957_;
	assign _0959_ = _0958_ | _0950_;
	assign _0960_ = _1905_ & ~_0914_;
	assign _0961_ = \mchip.vga.v_idx [3] & ~_0960_;
	assign _0962_ = _1904_ & ~_0961_;
	assign _0963_ = _0953_ & ~_0962_;
	assign _0964_ = _1900_ & ~_0963_;
	assign _0965_ = _0952_ & ~_0964_;
	assign _0966_ = _1909_ & ~_0965_;
	assign _0251_ = _0966_ | _0959_;
	assign _2116_[1] = \mchip.vga.h_idx [0] ^ \mchip.vga.h_idx [1];
	assign _0967_ = \mchip.vga.h_idx [0] & \mchip.vga.h_idx [1];
	assign _2116_[2] = _0967_ ^ \mchip.vga.h_idx [2];
	assign _0968_ = ~(\mchip.vga.h_idx [0] & \mchip.vga.h_idx [1]);
	assign _0969_ = \mchip.vga.h_idx [2] & ~_0968_;
	assign _2116_[3] = _0969_ ^ \mchip.vga.h_idx [3];
	assign _0970_ = ~(\mchip.vga.h_idx [2] & \mchip.vga.h_idx [3]);
	assign _0971_ = _0967_ & ~_0970_;
	assign _2116_[4] = _0971_ ^ \mchip.vga.h_idx [4];
	assign _0972_ = _0971_ & \mchip.vga.h_idx [4];
	assign _2116_[5] = _0972_ ^ \mchip.vga.h_idx [5];
	assign _0973_ = _0971_ & ~_0936_;
	assign _2116_[6] = _0973_ ^ \mchip.vga.h_idx [6];
	assign _0974_ = ~\mchip.vga.h_idx [6];
	assign _0975_ = _0973_ & ~_0974_;
	assign _2116_[7] = _0975_ ^ \mchip.vga.h_idx [7];
	assign _0976_ = _0971_ & _0937_;
	assign _2116_[8] = _0976_ ^ \mchip.vga.h_idx [8];
	assign _0977_ = _0976_ & \mchip.vga.h_idx [8];
	assign _2116_[9] = _0977_ ^ \mchip.vga.h_idx [9];
	assign _0978_ = \mchip.vga.v_idx [2] | \mchip.vga.v_idx [3];
	assign _0979_ = _0978_ | ~_0726_;
	assign _0980_ = _1904_ & ~_0979_;
	assign _0981_ = _0953_ & ~_0980_;
	assign _0982_ = _1900_ & ~_0981_;
	assign _0983_ = _0982_ | _0951_;
	assign _0984_ = _0980_ & ~_1901_;
	assign _0985_ = _0983_ & ~_0984_;
	assign _0986_ = ~(\mchip.vga.h_idx [8] | \mchip.vga.h_idx [7]);
	assign _0987_ = \mchip.vga.h_idx [9] & ~_0986_;
	assign _0988_ = _0985_ & ~_0987_;
	assign _0989_ = \mchip.vga.v_idx [7] | ~\mchip.vga.v_idx [6];
	assign _0990_ = _0720_ & ~_0989_;
	assign _0991_ = _0719_ & ~_0990_;
	assign _0992_ = \mchip.vga.v_idx [4] & ~\mchip.vga.v_idx [5];
	assign _0993_ = _0992_ & ~_0989_;
	assign _0994_ = _0914_ & _0717_;
	assign _0995_ = _0993_ & ~_0994_;
	assign _0996_ = _0991_ & ~_0995_;
	assign _0997_ = _1900_ & ~_0996_;
	assign _0998_ = _0997_ | _0951_;
	assign _0999_ = \mchip.vga.h_idx [8] & ~\mchip.vga.h_idx [9];
	assign _1000_ = ~_0999_;
	assign _1001_ = \mchip.vga.h_idx [6] & ~\mchip.vga.h_idx [7];
	assign _1002_ = _1001_ & ~_0941_;
	assign _1003_ = _1755_ & ~_1002_;
	assign _1004_ = \mchip.vga.h_idx [5] | ~\mchip.vga.h_idx [4];
	assign _1005_ = _1001_ & ~_1004_;
	assign _1006_ = _1005_ & ~_0971_;
	assign _1007_ = _1003_ & ~_1006_;
	assign _1008_ = ~(_1007_ | _1000_);
	assign _1009_ = ~(\mchip.vga.h_idx [9] | \mchip.vga.h_idx [8]);
	assign _1010_ = _1009_ | _1008_;
	assign _1011_ = _0999_ & ~_0968_;
	assign _1012_ = ~(_0942_ | _0941_);
	assign _1013_ = _1012_ & _1011_;
	assign _1014_ = _1013_ & ~_0970_;
	assign _1015_ = ~_1009_;
	assign _1016_ = \mchip.vga.h_idx [7] & ~_1012_;
	assign _1017_ = _0999_ & ~_1016_;
	assign _1018_ = _1015_ & ~_1017_;
	assign _1019_ = _1018_ | _1014_;
	assign _1020_ = _1019_ | _1010_;
	assign _1021_ = ~(_1020_ | _0998_);
	assign _1022_ = \mchip.vga.v_idx [6] | ~\mchip.vga.v_idx [7];
	assign _1023_ = _0720_ & ~_1022_;
	assign _1024_ = _0918_ | ~_1023_;
	assign _1025_ = _1900_ & ~_1024_;
	assign _1026_ = \mchip.vga.v_idx [7] & ~_1023_;
	assign _1027_ = _1900_ & ~_1026_;
	assign _1028_ = _0952_ & ~_1027_;
	assign _1029_ = _1028_ | _1025_;
	assign _1030_ = _1029_ | ~_1021_;
	assign _1031_ = _0719_ | \mchip.vga.v_idx [5];
	assign _1032_ = _0719_ | ~_1902_;
	assign _1033_ = _0954_ & ~_1032_;
	assign _1034_ = _1031_ & ~_1033_;
	assign _1035_ = _1900_ & ~_1034_;
	assign _1036_ = _1035_ | _0951_;
	assign _1037_ = ~(_1036_ | _1020_);
	assign _1038_ = \mchip.vga.v_idx [9] | ~\mchip.vga.v_idx [0];
	assign _1039_ = \mchip.vga.v_idx [1] | ~\mchip.vga.v_idx [2];
	assign _1040_ = \mchip.vga.v_idx [4] & \mchip.vga.v_idx [3];
	assign _1041_ = _1040_ & ~_1039_;
	assign _1042_ = \mchip.vga.v_idx [7] | ~\mchip.vga.v_idx [8];
	assign _1043_ = \mchip.vga.v_idx [5] | ~\mchip.vga.v_idx [6];
	assign _1044_ = ~(_1043_ | _1042_);
	assign _1045_ = ~(_1044_ & _1041_);
	assign _1046_ = ~(_1045_ | _1038_);
	assign _1047_ = _0923_ & ~_1042_;
	assign _1048_ = \mchip.vga.v_idx [8] & ~_1047_;
	assign _1049_ = ~(\mchip.vga.v_idx [2] & \mchip.vga.v_idx [1]);
	assign _1050_ = _1040_ & ~_1049_;
	assign _1051_ = _1044_ & ~_1050_;
	assign _1052_ = _1048_ & ~_1051_;
	assign _1053_ = _1052_ | \mchip.vga.v_idx [9];
	assign _1054_ = _1053_ | _1046_;
	assign _1055_ = _1054_ | ~_1037_;
	assign _1056_ = _1755_ | \mchip.vga.h_idx [5];
	assign _1057_ = \mchip.vga.h_idx [4] | ~\mchip.vga.h_idx [5];
	assign _1058_ = ~(_1057_ | _1755_);
	assign _1059_ = _1892_ & ~_0970_;
	assign _1060_ = _1058_ & ~_1059_;
	assign _1061_ = _1056_ & ~_1060_;
	assign _1062_ = _0999_ & ~_1061_;
	assign _1063_ = _1062_ | _1009_;
	assign _1064_ = \mchip.vga.h_idx [0] & ~\mchip.vga.h_idx [9];
	assign _1065_ = ~(\mchip.vga.h_idx [4] & \mchip.vga.h_idx [3]);
	assign _1066_ = \mchip.vga.h_idx [1] | ~\mchip.vga.h_idx [2];
	assign _1067_ = ~(_1066_ | _1065_);
	assign _1068_ = \mchip.vga.h_idx [5] | ~\mchip.vga.h_idx [6];
	assign _1069_ = ~(_1068_ | _1747_);
	assign _1070_ = ~(_1069_ & _1067_);
	assign _1071_ = _1064_ & ~_1070_;
	assign _1072_ = _0974_ & ~_1747_;
	assign _1073_ = \mchip.vga.h_idx [8] & ~_1072_;
	assign _1074_ = \mchip.vga.h_idx [1] & \mchip.vga.h_idx [2];
	assign _1075_ = _1074_ & ~_1065_;
	assign _1076_ = _1069_ & ~_1075_;
	assign _1077_ = _1073_ & ~_1076_;
	assign _1078_ = _1077_ | \mchip.vga.h_idx [9];
	assign _1079_ = _1078_ | _1071_;
	assign _1080_ = _1079_ | _1063_;
	assign _1081_ = _1080_ | _0998_;
	assign _1082_ = ~(_1081_ | _1029_);
	assign _1083_ = _1082_ ^ _1030_;
	assign _1084_ = \mchip.vga.h_idx [2] | ~\mchip.vga.h_idx [3];
	assign _1085_ = _0968_ & ~_1084_;
	assign _1086_ = \mchip.vga.h_idx [3] & ~_1085_;
	assign _1087_ = _0937_ & ~_1086_;
	assign _1088_ = _0937_ & ~_1087_;
	assign _1089_ = _1009_ & ~_1088_;
	assign _1090_ = ~(_1084_ | _1057_);
	assign _1091_ = _0999_ & ~_1755_;
	assign _1092_ = ~(_1091_ & _1090_);
	assign _1093_ = _0967_ & ~_1092_;
	assign _1094_ = _0970_ & ~_1057_;
	assign _1095_ = \mchip.vga.h_idx [5] & ~_1094_;
	assign _1096_ = _1091_ & ~_1095_;
	assign _1097_ = _1015_ & ~_1096_;
	assign _1098_ = _1097_ | _1093_;
	assign _1099_ = _1098_ | _1089_;
	assign _1100_ = _1099_ | _0998_;
	assign _1101_ = _1100_ | _1029_;
	assign _1102_ = _0935_ & ~_0941_;
	assign _1103_ = ~(\mchip.vga.h_idx [0] | \mchip.vga.h_idx [1]);
	assign _1104_ = _1103_ & ~_1084_;
	assign _1105_ = \mchip.vga.h_idx [3] & ~_1104_;
	assign _1106_ = _1102_ & ~_1105_;
	assign _1107_ = _0935_ & ~_1106_;
	assign _1108_ = _1009_ & ~_1107_;
	assign _1109_ = \mchip.vga.h_idx [1] | \mchip.vga.h_idx [2];
	assign _1110_ = ~(_1109_ | _1065_);
	assign _1111_ = \mchip.vga.h_idx [7] & ~\mchip.vga.h_idx [8];
	assign _1112_ = ~(\mchip.vga.h_idx [6] & \mchip.vga.h_idx [5]);
	assign _1113_ = _1111_ & ~_1112_;
	assign _1114_ = ~(_1113_ & _1110_);
	assign _1115_ = _1064_ & ~_1114_;
	assign _1116_ = ~_0986_;
	assign _1117_ = _1112_ & ~_1894_;
	assign _1118_ = _1116_ & ~_1117_;
	assign _1119_ = _1109_ & ~_1065_;
	assign _1120_ = _1113_ & ~_1119_;
	assign _1121_ = _1118_ & ~_1120_;
	assign _1122_ = _1121_ | \mchip.vga.h_idx [9];
	assign _1123_ = _1122_ | _1115_;
	assign _1124_ = _1123_ | _1108_;
	assign _1125_ = _1124_ | _0998_;
	assign _1126_ = ~(_1125_ | _1029_);
	assign _1127_ = _1126_ ^ _1101_;
	assign _1128_ = ~(_1127_ ^ _1083_);
	assign _1129_ = \mchip.vga.h_idx [3] | ~\mchip.vga.h_idx [2];
	assign _1130_ = _1129_ | _0967_;
	assign _1131_ = ~(_1130_ & _1753_);
	assign _1132_ = _1004_ | _0942_;
	assign _1133_ = _1131_ & ~_1132_;
	assign _1134_ = _1016_ & ~_1133_;
	assign _1135_ = _1009_ & ~_1134_;
	assign _1136_ = \mchip.vga.h_idx [4] | \mchip.vga.h_idx [3];
	assign _1137_ = ~(_1136_ | _1068_);
	assign _1138_ = _1064_ & ~_1894_;
	assign _1139_ = ~(_1138_ & _1137_);
	assign _1140_ = _1074_ & ~_1139_;
	assign _1141_ = \mchip.vga.h_idx [6] & ~_1137_;
	assign _1142_ = _1111_ & ~_1141_;
	assign _1143_ = _1116_ & ~_1142_;
	assign _1144_ = _1143_ | \mchip.vga.h_idx [9];
	assign _1145_ = _1144_ | _1140_;
	assign _1146_ = _1145_ | _1135_;
	assign _1147_ = _1146_ | _0998_;
	assign _1148_ = ~(_1147_ | _1029_);
	assign _1149_ = _1001_ & ~\mchip.vga.h_idx [5];
	assign _1150_ = _1755_ & ~_1149_;
	assign _1151_ = _1001_ & ~_1057_;
	assign _1152_ = _1103_ & ~_1129_;
	assign _1153_ = _1753_ & ~_1152_;
	assign _1154_ = _1151_ & ~_1153_;
	assign _1155_ = _1150_ & ~_1154_;
	assign _1156_ = _1009_ & ~_1155_;
	assign _1157_ = _1111_ & ~_1746_;
	assign _1158_ = _1896_ & ~_1066_;
	assign _1159_ = ~(_1158_ & _1157_);
	assign _1160_ = _1064_ & ~_1159_;
	assign _1161_ = _1896_ & ~_1074_;
	assign _1162_ = \mchip.vga.h_idx [4] & ~_1161_;
	assign _1163_ = _1157_ & ~_1162_;
	assign _1164_ = _1116_ & ~_1163_;
	assign _1165_ = _1164_ | \mchip.vga.h_idx [9];
	assign _1166_ = _1165_ | _1160_;
	assign _1167_ = _1166_ | _1156_;
	assign _1168_ = _1167_ | _0998_;
	assign _1169_ = ~(_1168_ | _1029_);
	assign _1170_ = _1169_ ^ _1148_;
	assign _1171_ = _1755_ | ~_0936_;
	assign _1172_ = _0936_ | _1755_;
	assign _1173_ = _0968_ & ~_1753_;
	assign _1174_ = _1173_ & ~_1172_;
	assign _1175_ = _1171_ & ~_1174_;
	assign _1176_ = _1009_ & ~_1175_;
	assign _1177_ = ~(_1057_ | _1753_);
	assign _1178_ = _1009_ & _1001_;
	assign _1179_ = ~(_1178_ & _1177_);
	assign _1180_ = _0967_ & ~_1179_;
	assign _1181_ = _1755_ | ~_1009_;
	assign _1182_ = \mchip.vga.h_idx [5] & ~_1177_;
	assign _1183_ = _1178_ & ~_1182_;
	assign _1184_ = _1181_ & ~_1183_;
	assign _1185_ = _1184_ | _1180_;
	assign _1186_ = _1185_ | _1176_;
	assign _1187_ = _1186_ | _0998_;
	assign _1188_ = _1187_ | _1029_;
	assign _1189_ = _1746_ | ~_0986_;
	assign _1190_ = \mchip.vga.h_idx [6] | ~\mchip.vga.h_idx [5];
	assign _1191_ = _0986_ & ~_1190_;
	assign _1192_ = _1896_ & ~_1109_;
	assign _1193_ = \mchip.vga.h_idx [4] & ~_1192_;
	assign _1194_ = _1191_ & ~_1193_;
	assign _1195_ = _1189_ & ~_1194_;
	assign _1196_ = _1195_ | \mchip.vga.h_idx [9];
	assign _1197_ = \mchip.vga.h_idx [1] | ~\mchip.vga.h_idx [0];
	assign _1198_ = _1197_ | _1753_;
	assign _1199_ = _1198_ | _1172_;
	assign _1200_ = _1009_ & ~_1199_;
	assign _1201_ = _1200_ | _1196_;
	assign _1202_ = _1892_ | _1753_;
	assign _1203_ = _0941_ | _1755_;
	assign _1204_ = _1203_ | _1202_;
	assign _1205_ = _1009_ & ~_1204_;
	assign _1206_ = _1205_ | _1201_;
	assign _1207_ = _1206_ | _0998_;
	assign _1208_ = ~(_1207_ | _1029_);
	assign _1209_ = _1208_ ^ _1188_;
	assign _1210_ = _1209_ ^ _1170_;
	assign _1211_ = ~(_1210_ ^ _1128_);
	assign _1212_ = _1036_ | _1080_;
	assign _1213_ = ~(_1212_ | _1054_);
	assign _1214_ = _1213_ ^ _1055_;
	assign _1215_ = _1036_ | _1099_;
	assign _1216_ = _1215_ | _1054_;
	assign _1217_ = _1036_ | _1124_;
	assign _1218_ = ~(_1217_ | _1054_);
	assign _1219_ = _1218_ ^ _1216_;
	assign _1220_ = _1219_ ^ _1214_;
	assign _1221_ = _1036_ | _1146_;
	assign _1222_ = ~(_1221_ | _1054_);
	assign _1223_ = _1036_ | _1167_;
	assign _1224_ = ~(_1223_ | _1054_);
	assign _1225_ = _1224_ ^ _1222_;
	assign _1226_ = _1036_ | _1186_;
	assign _1227_ = _1226_ | _1054_;
	assign _1228_ = _1036_ | _1206_;
	assign _1229_ = ~(_1228_ | _1054_);
	assign _1230_ = _1229_ ^ _1227_;
	assign _1231_ = _1230_ ^ _1225_;
	assign _1232_ = ~(_1231_ ^ _1220_);
	assign _1233_ = ~(_1232_ & _1211_);
	assign _1234_ = _1232_ | _1211_;
	assign _1235_ = ~(_1234_ & _1233_);
	assign _1236_ = _0929_ & ~_0961_;
	assign _1237_ = _0929_ & ~_1236_;
	assign _1238_ = _0951_ & ~_1237_;
	assign _1239_ = ~(_1238_ | _1020_);
	assign _1240_ = ~_0914_;
	assign _1241_ = _1905_ & _1902_;
	assign _1242_ = _1900_ & ~_0719_;
	assign _1243_ = ~(_1242_ & _1241_);
	assign _1244_ = ~(_1243_ | _1240_);
	assign _1245_ = _1902_ & ~_0717_;
	assign _1246_ = \mchip.vga.v_idx [5] & ~_1245_;
	assign _1247_ = _1242_ & ~_1246_;
	assign _1248_ = _0952_ & ~_1247_;
	assign _1249_ = _1248_ | _1244_;
	assign _1250_ = _1249_ | ~_1239_;
	assign _1251_ = _1238_ | _1080_;
	assign _1252_ = ~(_1251_ | _1249_);
	assign _1253_ = _1252_ ^ _1250_;
	assign _1254_ = _1238_ | _1099_;
	assign _1255_ = _1254_ | _1249_;
	assign _1256_ = _1238_ | _1124_;
	assign _1257_ = ~(_1256_ | _1249_);
	assign _1258_ = _1257_ ^ _1255_;
	assign _1259_ = _1258_ ^ _1253_;
	assign _1260_ = _1238_ | _1146_;
	assign _1261_ = ~(_1260_ | _1249_);
	assign _1262_ = _1238_ | _1167_;
	assign _1263_ = ~(_1262_ | _1249_);
	assign _1264_ = _1263_ ^ _1261_;
	assign _1265_ = _1238_ | _1186_;
	assign _1266_ = _1265_ | _1249_;
	assign _1267_ = _1238_ | _1206_;
	assign _1268_ = ~(_1267_ | _1249_);
	assign _1269_ = _1268_ ^ _1266_;
	assign _1270_ = _1269_ ^ _1264_;
	assign _1271_ = ~(_1270_ ^ _1259_);
	assign _1272_ = _0720_ & _1903_;
	assign _1273_ = _0726_ & _1905_;
	assign _1274_ = \mchip.vga.v_idx [3] & ~_1273_;
	assign _1275_ = _1272_ & ~_1274_;
	assign _1276_ = _1903_ & ~_1275_;
	assign _1277_ = _0951_ & ~_1276_;
	assign _1278_ = ~(_1277_ | _1020_);
	assign _1279_ = ~(\mchip.vga.v_idx [2] | \mchip.vga.v_idx [1]);
	assign _1280_ = _1279_ & _1040_;
	assign _1281_ = ~(\mchip.vga.v_idx [5] & \mchip.vga.v_idx [6]);
	assign _1282_ = \mchip.vga.v_idx [7] & ~\mchip.vga.v_idx [8];
	assign _1283_ = _1282_ & ~_1281_;
	assign _1284_ = ~(_1283_ & _1280_);
	assign _1285_ = ~(_1284_ | _1038_);
	assign _1286_ = \mchip.vga.v_idx [8] | \mchip.vga.v_idx [7];
	assign _1287_ = _1282_ & _1281_;
	assign _1288_ = _1286_ & ~_1287_;
	assign _1289_ = _1040_ & ~_1279_;
	assign _1290_ = _1283_ & ~_1289_;
	assign _1291_ = _1288_ & ~_1290_;
	assign _1292_ = _1291_ | \mchip.vga.v_idx [9];
	assign _1293_ = _1292_ | _1285_;
	assign _1294_ = _1293_ | ~_1278_;
	assign _1295_ = _1277_ | _1080_;
	assign _1296_ = ~(_1295_ | _1293_);
	assign _1297_ = _1296_ ^ _1294_;
	assign _1298_ = _1277_ | _1099_;
	assign _1299_ = _1298_ | _1293_;
	assign _1300_ = _1277_ | _1124_;
	assign _1301_ = ~(_1300_ | _1293_);
	assign _1302_ = _1301_ ^ _1299_;
	assign _1303_ = _1302_ ^ _1297_;
	assign _1304_ = _1277_ | _1146_;
	assign _1305_ = ~(_1304_ | _1293_);
	assign _1306_ = _1277_ | _1167_;
	assign _1307_ = ~(_1306_ | _1293_);
	assign _1308_ = _1307_ ^ _1305_;
	assign _1309_ = _1277_ | _1186_;
	assign _1310_ = _1309_ | _1293_;
	assign _1311_ = _1277_ | _1206_;
	assign _1312_ = ~(_1311_ | _1293_);
	assign _1313_ = _1312_ ^ _1310_;
	assign _1314_ = _1313_ ^ _1308_;
	assign _1315_ = _1314_ ^ _1303_;
	assign _1316_ = _1315_ | _1271_;
	assign _1317_ = ~(_1315_ & _1271_);
	assign _1318_ = _1317_ & _1316_;
	assign _1319_ = _1318_ ^ _1235_;
	assign _1320_ = _0992_ & ~_1022_;
	assign _1321_ = \mchip.vga.v_idx [3] | ~\mchip.vga.v_idx [2];
	assign _1322_ = ~(_1321_ | _0914_);
	assign _1323_ = _0978_ & ~_1322_;
	assign _1324_ = _1320_ & ~_1323_;
	assign _1325_ = _1026_ & ~_1324_;
	assign _1326_ = _0951_ & ~_1325_;
	assign _1327_ = ~(_1326_ | _1020_);
	assign _1328_ = \mchip.vga.v_idx [4] | \mchip.vga.v_idx [3];
	assign _1329_ = ~(_1328_ | _1043_);
	assign _1330_ = _1282_ & ~_1038_;
	assign _1331_ = ~(_1330_ & _1329_);
	assign _1332_ = ~(_1331_ | _1049_);
	assign _1333_ = \mchip.vga.v_idx [6] & ~_1329_;
	assign _1334_ = _1282_ & ~_1333_;
	assign _1335_ = _1286_ & ~_1334_;
	assign _1336_ = _1335_ | \mchip.vga.v_idx [9];
	assign _1337_ = _1336_ | _1332_;
	assign _1338_ = _1337_ | ~_1327_;
	assign _1339_ = _1326_ | _1080_;
	assign _1340_ = ~(_1339_ | _1337_);
	assign _1341_ = _1340_ ^ _1338_;
	assign _1342_ = _1326_ | _1099_;
	assign _1343_ = _1342_ | _1337_;
	assign _1344_ = _1326_ | _1124_;
	assign _1345_ = ~(_1344_ | _1337_);
	assign _1346_ = _1345_ ^ _1343_;
	assign _1347_ = _1346_ ^ _1341_;
	assign _1348_ = _1326_ | _1146_;
	assign _1349_ = ~(_1348_ | _1337_);
	assign _1350_ = _1326_ | _1167_;
	assign _1351_ = ~(_1350_ | _1337_);
	assign _1352_ = _1351_ ^ _1349_;
	assign _1353_ = _1326_ | _1186_;
	assign _1354_ = _1353_ | _1337_;
	assign _1355_ = _1326_ | _1206_;
	assign _1356_ = ~(_1355_ | _1337_);
	assign _1357_ = _1356_ ^ _1354_;
	assign _1358_ = _1357_ ^ _1352_;
	assign _1359_ = ~(_1358_ ^ _1347_);
	assign _1360_ = _0920_ & ~_0989_;
	assign _1361_ = _0719_ & ~_1360_;
	assign _1362_ = _1902_ & ~_0989_;
	assign _1363_ = _0726_ & ~_1321_;
	assign _1364_ = _0978_ & ~_1363_;
	assign _1365_ = _1362_ & ~_1364_;
	assign _1366_ = _1361_ & ~_1365_;
	assign _1367_ = _0951_ & ~_1366_;
	assign _1368_ = ~(_1367_ | _1020_);
	assign _1369_ = \mchip.vga.v_idx [3] | ~\mchip.vga.v_idx [4];
	assign _1370_ = ~(_1369_ | _1039_);
	assign _1371_ = \mchip.vga.v_idx [5] | \mchip.vga.v_idx [6];
	assign _1372_ = _1282_ & ~_1371_;
	assign _1373_ = ~(_1372_ & _1370_);
	assign _1374_ = ~(_1373_ | _1038_);
	assign _1375_ = _1049_ & ~_1369_;
	assign _1376_ = \mchip.vga.v_idx [4] & ~_1375_;
	assign _1377_ = _1372_ & ~_1376_;
	assign _1378_ = _1286_ & ~_1377_;
	assign _1379_ = _1378_ | \mchip.vga.v_idx [9];
	assign _1380_ = _1379_ | _1374_;
	assign _1381_ = _1368_ & ~_1380_;
	assign _1382_ = _1367_ | _1080_;
	assign _1383_ = ~(_1382_ | _1380_);
	assign _1384_ = _1383_ ^ _1381_;
	assign _1385_ = _1367_ | _1099_;
	assign _1386_ = _1385_ | _1380_;
	assign _1387_ = _1367_ | _1124_;
	assign _1388_ = ~(_1387_ | _1380_);
	assign _1389_ = _1388_ ^ _1386_;
	assign _1390_ = _1389_ ^ _1384_;
	assign _1391_ = _1367_ | _1146_;
	assign _1392_ = ~(_1391_ | _1380_);
	assign _1393_ = _1367_ | _1167_;
	assign _1394_ = ~(_1393_ | _1380_);
	assign _1395_ = _1394_ ^ _1392_;
	assign _1396_ = _1367_ | _1186_;
	assign _1397_ = _1396_ | _1380_;
	assign _1398_ = _1367_ | _1206_;
	assign _1399_ = ~(_1398_ | _1380_);
	assign _1400_ = _1399_ ^ _1397_;
	assign _1401_ = _1400_ ^ _1395_;
	assign _1402_ = _1401_ ^ _1390_;
	assign _1403_ = _1359_ | ~_1402_;
	assign _1404_ = _1402_ | ~_1359_;
	assign _1405_ = ~(_1404_ & _1403_);
	assign _1406_ = _0719_ | ~_0924_;
	assign _1407_ = _0924_ | _0719_;
	assign _1408_ = ~(_0978_ | _0914_);
	assign _1409_ = _1408_ & ~_1407_;
	assign _1410_ = _1406_ & ~_1409_;
	assign _1411_ = _0951_ & ~_1410_;
	assign _1412_ = _1411_ | _1020_;
	assign _1413_ = _1902_ & ~_0978_;
	assign _1414_ = _0951_ & ~_0989_;
	assign _1415_ = ~(_1414_ & _1413_);
	assign _1416_ = ~(_1415_ | _1240_);
	assign _1417_ = _0719_ | ~_0951_;
	assign _1418_ = \mchip.vga.v_idx [5] & ~_1413_;
	assign _1419_ = _1414_ & ~_1418_;
	assign _1420_ = _1417_ & ~_1419_;
	assign _1421_ = _1420_ | _1416_;
	assign _1422_ = _1421_ | _1412_;
	assign _1423_ = _1411_ | _1080_;
	assign _1424_ = ~(_1423_ | _1421_);
	assign _1425_ = _1424_ ^ _1422_;
	assign _1426_ = _1411_ | _1099_;
	assign _1427_ = _1426_ | _1421_;
	assign _1428_ = _1411_ | _1124_;
	assign _1429_ = ~(_1428_ | _1421_);
	assign _1430_ = _1429_ ^ _1427_;
	assign _1431_ = _1430_ ^ _1425_;
	assign _1432_ = _1411_ | _1146_;
	assign _1433_ = _1432_ | _1421_;
	assign _1434_ = _1411_ | _1167_;
	assign _1435_ = ~(_1434_ | _1421_);
	assign _1436_ = _1435_ ^ _1433_;
	assign _1437_ = _1411_ | _1186_;
	assign _1438_ = _1437_ | _1421_;
	assign _1439_ = _1411_ | _1206_;
	assign _1440_ = ~(_1439_ | _1421_);
	assign _1441_ = _1440_ ^ _1438_;
	assign _1442_ = _1441_ ^ _1436_;
	assign _1443_ = _1442_ ^ _1431_;
	assign _1444_ = _0979_ | _0721_;
	assign _1445_ = _0951_ & ~_1444_;
	assign _1446_ = _1445_ | _1020_;
	assign _1447_ = _0978_ | _0716_;
	assign _1448_ = _1447_ | _1407_;
	assign _1449_ = _0951_ & ~_1448_;
	assign _1450_ = _1371_ | _1286_;
	assign _1451_ = \mchip.vga.v_idx [5] & ~\mchip.vga.v_idx [6];
	assign _1452_ = _1451_ & ~_1286_;
	assign _1453_ = _1279_ & ~_1369_;
	assign _1454_ = \mchip.vga.v_idx [4] & ~_1453_;
	assign _1455_ = _1452_ & ~_1454_;
	assign _1456_ = _1450_ & ~_1455_;
	assign _1457_ = _1456_ | \mchip.vga.v_idx [9];
	assign _1458_ = _1457_ | _1449_;
	assign _1459_ = _1458_ | _1446_;
	assign _1460_ = _1445_ | _1080_;
	assign _1461_ = ~(_1460_ | _1458_);
	assign _1462_ = _1461_ ^ _1459_;
	assign _1463_ = _1445_ | _1099_;
	assign _1464_ = _1463_ | _1458_;
	assign _1465_ = _1445_ | _1124_;
	assign _1466_ = ~(_1465_ | _1458_);
	assign _1467_ = _1466_ ^ _1464_;
	assign _1468_ = _1467_ ^ _1462_;
	assign _1469_ = _1445_ | _1146_;
	assign _1470_ = _1469_ | _1458_;
	assign _1471_ = _1445_ | _1167_;
	assign _1472_ = ~(_1471_ | _1458_);
	assign _1473_ = _1472_ ^ _1470_;
	assign _1474_ = _1445_ | _1186_;
	assign _1475_ = _1474_ | _1458_;
	assign _1476_ = _1445_ | _1206_;
	assign _1477_ = ~(_1476_ | _1458_);
	assign _1478_ = _1477_ ^ _1475_;
	assign _1479_ = _1478_ ^ _1473_;
	assign _1480_ = _1479_ ^ _1468_;
	assign _1481_ = _1443_ | ~_1480_;
	assign _1482_ = _1480_ | ~_1443_;
	assign _1483_ = _1482_ & _1481_;
	assign _1484_ = _1483_ ^ _1405_;
	assign _1485_ = _1484_ ^ _1319_;
	assign _1486_ = _1232_ | ~_1211_;
	assign _1487_ = _1271_ | ~_1315_;
	assign _1488_ = ~(_1487_ | _1486_);
	assign _1489_ = _1402_ | _1359_;
	assign _1490_ = _1489_ | _1481_;
	assign _1491_ = _1488_ & ~_1490_;
	assign _1492_ = _1486_ | _1316_;
	assign _1493_ = _1480_ | _1443_;
	assign _1494_ = _1493_ | _1489_;
	assign _1495_ = _1494_ | _1492_;
	assign _1496_ = _1487_ | _1234_;
	assign _1497_ = _1496_ | _1494_;
	assign _1498_ = ~(_1493_ | _1489_);
	assign _1499_ = _1487_ | _1233_;
	assign _1500_ = _1498_ & ~_1499_;
	assign _1501_ = _1500_ | _1497_;
	assign _1502_ = _1486_ | _1317_;
	assign _1503_ = _1498_ & ~_1502_;
	assign _1504_ = _1501_ & ~_1503_;
	assign _1505_ = _1504_ | ~_1495_;
	assign _1506_ = _1493_ | _1404_;
	assign _1507_ = _1488_ & ~_1506_;
	assign _1508_ = _1505_ & ~_1507_;
	assign _1509_ = _1493_ | _1403_;
	assign _1510_ = _1488_ & ~_1509_;
	assign _1511_ = _1510_ | _1508_;
	assign _1512_ = _1489_ | _1482_;
	assign _1513_ = _1488_ & ~_1512_;
	assign _1514_ = _1511_ & ~_1513_;
	assign _1515_ = _1514_ | _1491_;
	assign _1516_ = _1485_ & ~_1515_;
	assign _1517_ = (_1516_ ? _1030_ : _1055_);
	assign _1518_ = _1500_ | ~_1497_;
	assign _1519_ = _1503_ | ~_1518_;
	assign _1520_ = _1495_ & ~_1519_;
	assign _1521_ = _1520_ | _1507_;
	assign _1522_ = ~(_1521_ | _1510_);
	assign _1523_ = _1522_ | _1513_;
	assign _1524_ = _1523_ | _1491_;
	assign _1525_ = _1485_ & ~_1524_;
	assign _1526_ = (_1516_ ? _1250_ : _1294_);
	assign _1527_ = (_1525_ ? _1517_ : _1526_);
	assign _1528_ = _1518_ | _1503_;
	assign _1529_ = _1495_ & ~_1528_;
	assign _1530_ = _1529_ | _1507_;
	assign _1531_ = _1530_ | _1510_;
	assign _1532_ = _1531_ | _1513_;
	assign _1533_ = _1532_ | _1491_;
	assign _1534_ = _1485_ & ~_1533_;
	assign _1535_ = ~_1381_;
	assign _1536_ = (_1516_ ? _1338_ : _1535_);
	assign _1537_ = (_1516_ ? _1422_ : _1459_);
	assign _1538_ = (_1525_ ? _1536_ : _1537_);
	assign _1539_ = (_1534_ ? _1527_ : _1538_);
	assign _1540_ = (_1516_ ? _1082_ : _1213_);
	assign _1541_ = (_1516_ ? _1252_ : _1296_);
	assign _1542_ = (_1525_ ? _1540_ : _1541_);
	assign _1543_ = (_1516_ ? _1340_ : _1383_);
	assign _1544_ = (_1516_ ? _1424_ : _1461_);
	assign _1545_ = (_1525_ ? _1543_ : _1544_);
	assign _1546_ = (_1534_ ? _1542_ : _1545_);
	assign _1547_ = ~(_1546_ & _1539_);
	assign _1548_ = _1546_ | _1539_;
	assign _1549_ = _1548_ & _1547_;
	assign _1550_ = (_1516_ ? _1101_ : _1216_);
	assign _1551_ = (_1516_ ? _1255_ : _1299_);
	assign _1552_ = (_1525_ ? _1550_ : _1551_);
	assign _1553_ = (_1516_ ? _1343_ : _1386_);
	assign _1554_ = (_1516_ ? _1427_ : _1464_);
	assign _1555_ = (_1525_ ? _1553_ : _1554_);
	assign _1556_ = (_1534_ ? _1552_ : _1555_);
	assign _1557_ = (_1516_ ? _1126_ : _1218_);
	assign _1558_ = (_1516_ ? _1257_ : _1301_);
	assign _1559_ = (_1525_ ? _1557_ : _1558_);
	assign _1560_ = (_1516_ ? _1345_ : _1388_);
	assign _1561_ = (_1516_ ? _1429_ : _1466_);
	assign _1562_ = (_1525_ ? _1560_ : _1561_);
	assign _1563_ = (_1534_ ? _1559_ : _1562_);
	assign _1564_ = ~(_1563_ & _1556_);
	assign _1565_ = _1563_ | _1556_;
	assign _1566_ = _1565_ & _1564_;
	assign _1567_ = _1566_ ^ _1549_;
	assign _1568_ = ~_1148_;
	assign _1569_ = ~_1222_;
	assign _1570_ = (_1516_ ? _1568_ : _1569_);
	assign _1571_ = ~_1261_;
	assign _1572_ = ~_1305_;
	assign _1573_ = (_1516_ ? _1571_ : _1572_);
	assign _1574_ = (_1525_ ? _1570_ : _1573_);
	assign _1575_ = ~_1349_;
	assign _1576_ = ~_1392_;
	assign _1577_ = (_1516_ ? _1575_ : _1576_);
	assign _1578_ = (_1516_ ? _1433_ : _1470_);
	assign _1579_ = (_1525_ ? _1577_ : _1578_);
	assign _1580_ = (_1534_ ? _1574_ : _1579_);
	assign _1581_ = (_1516_ ? _1169_ : _1224_);
	assign _1582_ = (_1516_ ? _1263_ : _1307_);
	assign _1583_ = (_1525_ ? _1581_ : _1582_);
	assign _1584_ = (_1516_ ? _1351_ : _1394_);
	assign _1585_ = (_1516_ ? _1435_ : _1472_);
	assign _1586_ = (_1525_ ? _1584_ : _1585_);
	assign _1587_ = (_1534_ ? _1583_ : _1586_);
	assign _1588_ = ~(_1587_ & _1580_);
	assign _1589_ = _1587_ | _1580_;
	assign _1590_ = ~(_1589_ & _1588_);
	assign _1591_ = ~_1188_;
	assign _1592_ = ~_1227_;
	assign _1593_ = (_1516_ ? _1591_ : _1592_);
	assign _1594_ = ~_1266_;
	assign _1595_ = ~_1310_;
	assign _1596_ = (_1516_ ? _1594_ : _1595_);
	assign _1597_ = (_1525_ ? _1593_ : _1596_);
	assign _1598_ = ~_1354_;
	assign _1599_ = ~_1397_;
	assign _1600_ = (_1516_ ? _1598_ : _1599_);
	assign _1601_ = ~_1438_;
	assign _1602_ = ~_1475_;
	assign _1603_ = (_1516_ ? _1601_ : _1602_);
	assign _1604_ = (_1525_ ? _1600_ : _1603_);
	assign _1605_ = (_1534_ ? _1597_ : _1604_);
	assign _1606_ = (_1516_ ? _1208_ : _1229_);
	assign _1607_ = (_1516_ ? _1268_ : _1312_);
	assign _1608_ = (_1525_ ? _1606_ : _1607_);
	assign _1609_ = (_1516_ ? _1356_ : _1399_);
	assign _1610_ = (_1516_ ? _1440_ : _1477_);
	assign _1611_ = (_1525_ ? _1609_ : _1610_);
	assign _1612_ = (_1534_ ? _1608_ : _1611_);
	assign _1613_ = _1605_ | ~_1612_;
	assign _1614_ = _1612_ | ~_1605_;
	assign _1615_ = _1614_ & _1613_;
	assign _1616_ = _1615_ ^ _1590_;
	assign _1617_ = ~(_1616_ ^ _1567_);
	assign _1618_ = ~_1617_;
	assign _1619_ = _1546_ | ~_1539_;
	assign _1620_ = _1563_ | ~_1556_;
	assign _1621_ = ~(_1620_ | _1619_);
	assign _1622_ = _1587_ | ~_1580_;
	assign _1623_ = _1622_ | _1613_;
	assign _1624_ = _1621_ & ~_1623_;
	assign _1625_ = _1619_ | _1564_;
	assign _1626_ = _1612_ | _1605_;
	assign _1627_ = _1626_ | _1622_;
	assign _1628_ = _1627_ | _1625_;
	assign _1629_ = _1620_ | _1548_;
	assign _1630_ = _1629_ | _1627_;
	assign _1631_ = ~(_1626_ | _1622_);
	assign _1632_ = _1620_ | _1547_;
	assign _1633_ = _1631_ & ~_1632_;
	assign _1634_ = _1633_ | _1630_;
	assign _1635_ = _1619_ | _1565_;
	assign _1636_ = _1631_ & ~_1635_;
	assign _1637_ = _1634_ & ~_1636_;
	assign _1638_ = _1637_ | ~_1628_;
	assign _1639_ = _1626_ | _1589_;
	assign _1640_ = _1621_ & ~_1639_;
	assign _1641_ = _1638_ & ~_1640_;
	assign _1642_ = _1626_ | _1588_;
	assign _1643_ = _1621_ & ~_1642_;
	assign _1644_ = _1643_ | _1641_;
	assign _1645_ = _1622_ | _1614_;
	assign _1646_ = _1621_ & ~_1645_;
	assign _1647_ = _1644_ & ~_1646_;
	assign _1648_ = _1647_ | _1624_;
	assign _1649_ = _1648_ | _1618_;
	assign _1650_ = (_1649_ ? \mchip.row_sel[7].col_sel[6].tile_state.state  : \mchip.row_sel[7].col_sel[7].tile_state.state );
	assign _1651_ = _1633_ | ~_1630_;
	assign _1652_ = _1636_ | ~_1651_;
	assign _1653_ = _1628_ & ~_1652_;
	assign _1654_ = _1653_ | _1640_;
	assign _1655_ = ~(_1654_ | _1643_);
	assign _1656_ = _1655_ | _1646_;
	assign _1657_ = _1656_ | _1624_;
	assign _1658_ = _1617_ & ~_1657_;
	assign _1659_ = (_1649_ ? \mchip.row_sel[7].col_sel[4].tile_state.state  : \mchip.row_sel[7].col_sel[5].tile_state.state );
	assign _1660_ = (_1658_ ? _1650_ : _1659_);
	assign _1661_ = _1651_ | _1636_;
	assign _1662_ = _1628_ & ~_1661_;
	assign _1663_ = _1662_ | _1640_;
	assign _1664_ = _1663_ | _1643_;
	assign _1665_ = _1664_ | _1646_;
	assign _1666_ = _1665_ | _1624_;
	assign _1667_ = _1617_ & ~_1666_;
	assign _1668_ = (_1649_ ? \mchip.row_sel[7].col_sel[2].tile_state.state  : \mchip.row_sel[7].col_sel[3].tile_state.state );
	assign _1669_ = (_1649_ ? \mchip.row_sel[7].col_sel[0].tile_state.state  : \mchip.row_sel[7].col_sel[1].tile_state.state );
	assign _1670_ = (_1658_ ? _1668_ : _1669_);
	assign _1671_ = (_1667_ ? _1660_ : _1670_);
	assign _1672_ = (_1649_ ? \mchip.row_sel[6].col_sel[6].tile_state.state  : \mchip.row_sel[6].col_sel[7].tile_state.state );
	assign _1673_ = (_1649_ ? \mchip.row_sel[6].col_sel[4].tile_state.state  : \mchip.row_sel[6].col_sel[5].tile_state.state );
	assign _1674_ = (_1658_ ? _1672_ : _1673_);
	assign _1675_ = (_1649_ ? \mchip.row_sel[6].col_sel[2].tile_state.state  : \mchip.row_sel[6].col_sel[3].tile_state.state );
	assign _1676_ = (_1649_ ? \mchip.row_sel[6].col_sel[0].tile_state.state  : \mchip.row_sel[6].col_sel[1].tile_state.state );
	assign _1677_ = (_1658_ ? _1675_ : _1676_);
	assign _1678_ = (_1667_ ? _1674_ : _1677_);
	assign _1679_ = (_1516_ ? _1671_ : _1678_);
	assign _1680_ = (_1649_ ? \mchip.row_sel[5].col_sel[6].tile_state.state  : \mchip.row_sel[5].col_sel[7].tile_state.state );
	assign _1681_ = (_1649_ ? \mchip.row_sel[5].col_sel[4].tile_state.state  : \mchip.row_sel[5].col_sel[5].tile_state.state );
	assign _1682_ = (_1658_ ? _1680_ : _1681_);
	assign _1683_ = (_1649_ ? \mchip.row_sel[5].col_sel[2].tile_state.state  : \mchip.row_sel[5].col_sel[3].tile_state.state );
	assign _1684_ = (_1649_ ? \mchip.row_sel[5].col_sel[0].tile_state.state  : \mchip.row_sel[5].col_sel[1].tile_state.state );
	assign _1685_ = (_1658_ ? _1683_ : _1684_);
	assign _1686_ = (_1667_ ? _1682_ : _1685_);
	assign _1687_ = (_1649_ ? \mchip.row_sel[4].col_sel[6].tile_state.state  : \mchip.row_sel[4].col_sel[7].tile_state.state );
	assign _1688_ = (_1649_ ? \mchip.row_sel[4].col_sel[4].tile_state.state  : \mchip.row_sel[4].col_sel[5].tile_state.state );
	assign _1689_ = (_1658_ ? _1687_ : _1688_);
	assign _1690_ = (_1649_ ? \mchip.row_sel[4].col_sel[2].tile_state.state  : \mchip.row_sel[4].col_sel[3].tile_state.state );
	assign _1691_ = (_1649_ ? \mchip.row_sel[4].col_sel[0].tile_state.state  : \mchip.row_sel[4].col_sel[1].tile_state.state );
	assign _1692_ = (_1658_ ? _1690_ : _1691_);
	assign _1693_ = (_1667_ ? _1689_ : _1692_);
	assign _1694_ = (_1516_ ? _1686_ : _1693_);
	assign _1695_ = (_1525_ ? _1679_ : _1694_);
	assign _1696_ = (_1649_ ? \mchip.row_sel[3].col_sel[6].tile_state.state  : \mchip.row_sel[3].col_sel[7].tile_state.state );
	assign _1697_ = (_1649_ ? \mchip.row_sel[3].col_sel[4].tile_state.state  : \mchip.row_sel[3].col_sel[5].tile_state.state );
	assign _1698_ = (_1658_ ? _1696_ : _1697_);
	assign _1699_ = (_1649_ ? \mchip.row_sel[3].col_sel[2].tile_state.state  : \mchip.row_sel[3].col_sel[3].tile_state.state );
	assign _1700_ = (_1649_ ? \mchip.row_sel[3].col_sel[0].tile_state.state  : \mchip.row_sel[3].col_sel[1].tile_state.state );
	assign _1701_ = (_1658_ ? _1699_ : _1700_);
	assign _1702_ = (_1667_ ? _1698_ : _1701_);
	assign _1703_ = (_1649_ ? \mchip.row_sel[2].col_sel[6].tile_state.state  : \mchip.row_sel[2].col_sel[7].tile_state.state );
	assign _1704_ = (_1649_ ? \mchip.row_sel[2].col_sel[4].tile_state.state  : \mchip.row_sel[2].col_sel[5].tile_state.state );
	assign _1705_ = (_1658_ ? _1703_ : _1704_);
	assign _1706_ = (_1649_ ? \mchip.row_sel[2].col_sel[2].tile_state.state  : \mchip.row_sel[2].col_sel[3].tile_state.state );
	assign _1707_ = (_1649_ ? \mchip.row_sel[2].col_sel[0].tile_state.state  : \mchip.row_sel[2].col_sel[1].tile_state.state );
	assign _1708_ = (_1658_ ? _1706_ : _1707_);
	assign _1709_ = (_1667_ ? _1705_ : _1708_);
	assign _1710_ = (_1516_ ? _1702_ : _1709_);
	assign _1711_ = (_1649_ ? \mchip.row_sel[1].col_sel[6].tile_state.state  : \mchip.row_sel[1].col_sel[7].tile_state.state );
	assign _1712_ = (_1649_ ? \mchip.row_sel[1].col_sel[4].tile_state.state  : \mchip.row_sel[1].col_sel[5].tile_state.state );
	assign _1713_ = (_1658_ ? _1711_ : _1712_);
	assign _1714_ = (_1649_ ? \mchip.row_sel[1].col_sel[2].tile_state.state  : \mchip.row_sel[1].col_sel[3].tile_state.state );
	assign _1715_ = (_1649_ ? \mchip.row_sel[1].col_sel[0].tile_state.state  : \mchip.row_sel[1].col_sel[1].tile_state.state );
	assign _1716_ = (_1658_ ? _1714_ : _1715_);
	assign _1717_ = (_1667_ ? _1713_ : _1716_);
	assign _1718_ = (_1649_ ? \mchip.row_sel[0].col_sel[6].tile_state.state  : \mchip.row_sel[0].col_sel[7].tile_state.state );
	assign _1719_ = (_1649_ ? \mchip.row_sel[0].col_sel[4].tile_state.state  : \mchip.row_sel[0].col_sel[5].tile_state.state );
	assign _1720_ = (_1658_ ? _1718_ : _1719_);
	assign _1721_ = (_1649_ ? \mchip.row_sel[0].col_sel[2].tile_state.state  : \mchip.row_sel[0].col_sel[3].tile_state.state );
	assign _1722_ = (_1649_ ? \mchip.row_sel[0].col_sel[0].tile_state.state  : \mchip.row_sel[0].col_sel[1].tile_state.state );
	assign _1723_ = (_1658_ ? _1721_ : _1722_);
	assign _1724_ = (_1667_ ? _1720_ : _1723_);
	assign _1725_ = (_1516_ ? _1717_ : _1724_);
	assign _1726_ = (_1525_ ? _1710_ : _1725_);
	assign _1727_ = (_1534_ ? _1695_ : _1726_);
	assign _1728_ = ~(_1727_ & _1617_);
	assign \mchip.gn16  = _0988_ & ~_1728_;
	assign _1729_ = _1727_ | _1618_;
	assign \mchip.gp23  = _0988_ & ~_1729_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [0] <= 1'h0;
		else
			\mchip.vga.frame_count [0] <= _0071_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [1] <= 1'h0;
		else
			\mchip.vga.frame_count [1] <= _0082_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [2] <= 1'h0;
		else
			\mchip.vga.frame_count [2] <= _0093_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [3] <= 1'h0;
		else
			\mchip.vga.frame_count [3] <= _0096_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [4] <= 1'h0;
		else
			\mchip.vga.frame_count [4] <= _0097_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [5] <= 1'h0;
		else
			\mchip.vga.frame_count [5] <= _0098_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [6] <= 1'h0;
		else
			\mchip.vga.frame_count [6] <= _0099_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [7] <= 1'h0;
		else
			\mchip.vga.frame_count [7] <= _0100_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [8] <= 1'h0;
		else
			\mchip.vga.frame_count [8] <= _0101_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [9] <= 1'h0;
		else
			\mchip.vga.frame_count [9] <= _0102_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [10] <= 1'h0;
		else
			\mchip.vga.frame_count [10] <= _0072_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [11] <= 1'h0;
		else
			\mchip.vga.frame_count [11] <= _0073_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [12] <= 1'h0;
		else
			\mchip.vga.frame_count [12] <= _0074_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [13] <= 1'h0;
		else
			\mchip.vga.frame_count [13] <= _0075_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [14] <= 1'h0;
		else
			\mchip.vga.frame_count [14] <= _0076_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [15] <= 1'h0;
		else
			\mchip.vga.frame_count [15] <= _0077_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [16] <= 1'h0;
		else
			\mchip.vga.frame_count [16] <= _0078_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [17] <= 1'h0;
		else
			\mchip.vga.frame_count [17] <= _0079_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [18] <= 1'h0;
		else
			\mchip.vga.frame_count [18] <= _0080_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [19] <= 1'h0;
		else
			\mchip.vga.frame_count [19] <= _0081_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [20] <= 1'h0;
		else
			\mchip.vga.frame_count [20] <= _0083_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [21] <= 1'h0;
		else
			\mchip.vga.frame_count [21] <= _0084_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [22] <= 1'h0;
		else
			\mchip.vga.frame_count [22] <= _0085_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [23] <= 1'h0;
		else
			\mchip.vga.frame_count [23] <= _0086_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [24] <= 1'h0;
		else
			\mchip.vga.frame_count [24] <= _0087_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [25] <= 1'h0;
		else
			\mchip.vga.frame_count [25] <= _0088_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [26] <= 1'h0;
		else
			\mchip.vga.frame_count [26] <= _0089_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [27] <= 1'h0;
		else
			\mchip.vga.frame_count [27] <= _0090_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [28] <= 1'h0;
		else
			\mchip.vga.frame_count [28] <= _0091_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [29] <= 1'h0;
		else
			\mchip.vga.frame_count [29] <= _0092_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [30] <= 1'h0;
		else
			\mchip.vga.frame_count [30] <= _0094_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.frame_count [31] <= 1'h0;
		else
			\mchip.vga.frame_count [31] <= _0095_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[4].tile_state.state_locked  <= 1'h0;
		else if (_0166_)
			\mchip.row_sel[3].col_sel[4].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[4].tile_state.state  <= 1'h0;
		else if (_0035_)
			\mchip.row_sel[3].col_sel[4].tile_state.state  <= _0167_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[7].tile_state.state_locked  <= 1'h0;
		else if (_0156_)
			\mchip.row_sel[2].col_sel[7].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[7].tile_state.state  <= 1'h0;
		else if (_0040_)
			\mchip.row_sel[2].col_sel[7].tile_state.state  <= _0157_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[6].tile_state.state_locked  <= 1'h0;
		else if (_0218_)
			\mchip.row_sel[6].col_sel[6].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[6].tile_state.state  <= 1'h0;
		else if (_0009_)
			\mchip.row_sel[6].col_sel[6].tile_state.state  <= _0219_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[7].tile_state.state_locked  <= 1'h0;
		else if (_0140_)
			\mchip.row_sel[1].col_sel[7].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[7].tile_state.state  <= 1'h0;
		else if (_0048_)
			\mchip.row_sel[1].col_sel[7].tile_state.state  <= _0141_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[7].tile_state.state_locked  <= 1'h0;
		else if (_0172_)
			\mchip.row_sel[3].col_sel[7].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[7].tile_state.state  <= 1'h0;
		else if (_0032_)
			\mchip.row_sel[3].col_sel[7].tile_state.state  <= _0173_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[0].tile_state.state_locked  <= 1'h0;
		else if (_0206_)
			\mchip.row_sel[6].col_sel[0].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[0].tile_state.state  <= 1'h0;
		else if (_0015_)
			\mchip.row_sel[6].col_sel[0].tile_state.state  <= _0207_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[4].tile_state.state_locked  <= 1'h0;
		else if (_0198_)
			\mchip.row_sel[5].col_sel[4].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[4].tile_state.state  <= 1'h0;
		else if (_0019_)
			\mchip.row_sel[5].col_sel[4].tile_state.state  <= _0199_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[1].tile_state.state_locked  <= 1'h0;
		else if (_0176_)
			\mchip.row_sel[4].col_sel[1].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[1].tile_state.state  <= 1'h0;
		else if (_0030_)
			\mchip.row_sel[4].col_sel[1].tile_state.state  <= _0177_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[6].tile_state.state_locked  <= 1'h0;
		else if (_0138_)
			\mchip.row_sel[1].col_sel[6].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[6].tile_state.state  <= 1'h0;
		else if (_0049_)
			\mchip.row_sel[1].col_sel[6].tile_state.state  <= _0139_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[7].tile_state.state_locked  <= 1'h0;
		else if (_0220_)
			\mchip.row_sel[6].col_sel[7].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[7].tile_state.state  <= 1'h0;
		else if (_0008_)
			\mchip.row_sel[6].col_sel[7].tile_state.state  <= _0221_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[6].tile_state.state_locked  <= 1'h0;
		else if (_0154_)
			\mchip.row_sel[2].col_sel[6].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[6].tile_state.state  <= 1'h0;
		else if (_0041_)
			\mchip.row_sel[2].col_sel[6].tile_state.state  <= _0155_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[3].tile_state.state_locked  <= 1'h0;
		else if (_0180_)
			\mchip.row_sel[4].col_sel[3].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[3].tile_state.state  <= 1'h0;
		else if (_0028_)
			\mchip.row_sel[4].col_sel[3].tile_state.state  <= _0181_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[3].tile_state.state_locked  <= 1'h0;
		else if (_0164_)
			\mchip.row_sel[3].col_sel[3].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[3].tile_state.state  <= 1'h0;
		else if (_0036_)
			\mchip.row_sel[3].col_sel[3].tile_state.state  <= _0165_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[5].tile_state.state_locked  <= 1'h0;
		else if (_0136_)
			\mchip.row_sel[1].col_sel[5].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[5].tile_state.state  <= 1'h0;
		else if (_0050_)
			\mchip.row_sel[1].col_sel[5].tile_state.state  <= _0137_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[1].tile_state.state_locked  <= 1'h0;
		else if (_0208_)
			\mchip.row_sel[6].col_sel[1].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[1].tile_state.state  <= 1'h0;
		else if (_0014_)
			\mchip.row_sel[6].col_sel[1].tile_state.state  <= _0209_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[0].tile_state.state_locked  <= 1'h0;
		else if (_0222_)
			\mchip.row_sel[7].col_sel[0].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[0].tile_state.state  <= 1'h0;
		else if (_0007_)
			\mchip.row_sel[7].col_sel[0].tile_state.state  <= _0223_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[0].tile_state.state_locked  <= 1'h0;
		else if (_0190_)
			\mchip.row_sel[5].col_sel[0].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[0].tile_state.state  <= 1'h0;
		else if (_0023_)
			\mchip.row_sel[5].col_sel[0].tile_state.state  <= _0191_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[5].tile_state.state_locked  <= 1'h0;
		else if (_0152_)
			\mchip.row_sel[2].col_sel[5].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[5].tile_state.state  <= 1'h0;
		else if (_0042_)
			\mchip.row_sel[2].col_sel[5].tile_state.state  <= _0153_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[4].tile_state.state_locked  <= 1'h0;
		else if (_0134_)
			\mchip.row_sel[1].col_sel[4].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[4].tile_state.state  <= 1'h0;
		else if (_0051_)
			\mchip.row_sel[1].col_sel[4].tile_state.state  <= _0135_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[2].tile_state.state_locked  <= 1'h0;
		else if (_0194_)
			\mchip.row_sel[5].col_sel[2].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[2].tile_state.state  <= 1'h0;
		else if (_0021_)
			\mchip.row_sel[5].col_sel[2].tile_state.state  <= _0195_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[5].tile_state.state_locked  <= 1'h0;
		else if (_0200_)
			\mchip.row_sel[5].col_sel[5].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[5].tile_state.state  <= 1'h0;
		else if (_0018_)
			\mchip.row_sel[5].col_sel[5].tile_state.state  <= _0201_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[1].tile_state.state_locked  <= 1'h0;
		else if (_0224_)
			\mchip.row_sel[7].col_sel[1].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[1].tile_state.state  <= 1'h0;
		else if (_0006_)
			\mchip.row_sel[7].col_sel[1].tile_state.state  <= _0225_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[6].tile_state.state_locked  <= 1'h0;
		else if (_0170_)
			\mchip.row_sel[3].col_sel[6].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[6].tile_state.state  <= 1'h0;
		else if (_0033_)
			\mchip.row_sel[3].col_sel[6].tile_state.state  <= _0171_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[3].tile_state.state_locked  <= 1'h0;
		else if (_0132_)
			\mchip.row_sel[1].col_sel[3].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[3].tile_state.state  <= 1'h0;
		else if (_0052_)
			\mchip.row_sel[1].col_sel[3].tile_state.state  <= _0133_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[2].tile_state.state_locked  <= 1'h0;
		else if (_0210_)
			\mchip.row_sel[6].col_sel[2].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[2].tile_state.state  <= 1'h0;
		else if (_0013_)
			\mchip.row_sel[6].col_sel[2].tile_state.state  <= _0211_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[4].tile_state.state_locked  <= 1'h0;
		else if (_0150_)
			\mchip.row_sel[2].col_sel[4].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[4].tile_state.state  <= 1'h0;
		else if (_0043_)
			\mchip.row_sel[2].col_sel[4].tile_state.state  <= _0151_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[2].tile_state.state_locked  <= 1'h0;
		else if (_0162_)
			\mchip.row_sel[3].col_sel[2].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[2].tile_state.state  <= 1'h0;
		else if (_0037_)
			\mchip.row_sel[3].col_sel[2].tile_state.state  <= _0163_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[2].tile_state.state_locked  <= 1'h0;
		else if (_0226_)
			\mchip.row_sel[7].col_sel[2].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[2].tile_state.state  <= 1'h0;
		else if (_0005_)
			\mchip.row_sel[7].col_sel[2].tile_state.state  <= _0227_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[2].tile_state.state_locked  <= 1'h0;
		else if (_0130_)
			\mchip.row_sel[1].col_sel[2].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[2].tile_state.state  <= 1'h0;
		else if (_0053_)
			\mchip.row_sel[1].col_sel[2].tile_state.state  <= _0131_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[2].tile_state.state_locked  <= 1'h0;
		else if (_0178_)
			\mchip.row_sel[4].col_sel[2].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[2].tile_state.state  <= 1'h0;
		else if (_0029_)
			\mchip.row_sel[4].col_sel[2].tile_state.state  <= _0179_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[7].tile_state.state_locked  <= 1'h0;
		else if (_0188_)
			\mchip.row_sel[4].col_sel[7].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[7].tile_state.state  <= 1'h0;
		else if (_0024_)
			\mchip.row_sel[4].col_sel[7].tile_state.state  <= _0189_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[0].tile_state.state_locked  <= 1'h0;
		else if (_0174_)
			\mchip.row_sel[4].col_sel[0].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[0].tile_state.state  <= 1'h0;
		else if (_0031_)
			\mchip.row_sel[4].col_sel[0].tile_state.state  <= _0175_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[3].tile_state.state_locked  <= 1'h0;
		else if (_0148_)
			\mchip.row_sel[2].col_sel[3].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[3].tile_state.state  <= 1'h0;
		else if (_0044_)
			\mchip.row_sel[2].col_sel[3].tile_state.state  <= _0149_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[1].tile_state.state_locked  <= 1'h0;
		else if (_0128_)
			\mchip.row_sel[1].col_sel[1].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[1].tile_state.state  <= 1'h0;
		else if (_0054_)
			\mchip.row_sel[1].col_sel[1].tile_state.state  <= _0129_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[3].tile_state.state_locked  <= 1'h0;
		else if (_0228_)
			\mchip.row_sel[7].col_sel[3].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[3].tile_state.state  <= 1'h0;
		else if (_0004_)
			\mchip.row_sel[7].col_sel[3].tile_state.state  <= _0229_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[3].tile_state.state_locked  <= 1'h0;
		else if (_0212_)
			\mchip.row_sel[6].col_sel[3].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[3].tile_state.state  <= 1'h0;
		else if (_0012_)
			\mchip.row_sel[6].col_sel[3].tile_state.state  <= _0213_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[6].tile_state.state_locked  <= 1'h0;
		else if (_0202_)
			\mchip.row_sel[5].col_sel[6].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[6].tile_state.state  <= 1'h0;
		else if (_0017_)
			\mchip.row_sel[5].col_sel[6].tile_state.state  <= _0203_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[1].tile_state.state_locked  <= 1'h0;
		else if (_0160_)
			\mchip.row_sel[3].col_sel[1].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[1].tile_state.state  <= 1'h0;
		else if (_0038_)
			\mchip.row_sel[3].col_sel[1].tile_state.state  <= _0161_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[0].tile_state.state_locked  <= 1'h0;
		else if (_0126_)
			\mchip.row_sel[1].col_sel[0].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[1].col_sel[0].tile_state.state  <= 1'h0;
		else if (_0055_)
			\mchip.row_sel[1].col_sel[0].tile_state.state  <= _0127_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[4].tile_state.state_locked  <= 1'h0;
		else if (_0182_)
			\mchip.row_sel[4].col_sel[4].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[4].tile_state.state  <= 1'h0;
		else if (_0027_)
			\mchip.row_sel[4].col_sel[4].tile_state.state  <= _0183_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[4].tile_state.state_locked  <= 1'h0;
		else if (_0230_)
			\mchip.row_sel[7].col_sel[4].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[4].tile_state.state  <= 1'h0;
		else if (_0003_)
			\mchip.row_sel[7].col_sel[4].tile_state.state  <= _0231_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[2].tile_state.state_locked  <= 1'h0;
		else if (_0146_)
			\mchip.row_sel[2].col_sel[2].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[2].tile_state.state  <= 1'h0;
		else if (_0045_)
			\mchip.row_sel[2].col_sel[2].tile_state.state  <= _0147_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[5].tile_state.state_locked  <= 1'h0;
		else if (_0168_)
			\mchip.row_sel[3].col_sel[5].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[5].tile_state.state  <= 1'h0;
		else if (_0034_)
			\mchip.row_sel[3].col_sel[5].tile_state.state  <= _0169_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[7].tile_state.state_locked  <= 1'h0;
		else if (_0124_)
			\mchip.row_sel[0].col_sel[7].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[7].tile_state.state  <= 1'h0;
		else if (_0056_)
			\mchip.row_sel[0].col_sel[7].tile_state.state  <= _0125_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[4].tile_state.state_locked  <= 1'h0;
		else if (_0214_)
			\mchip.row_sel[6].col_sel[4].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[4].tile_state.state  <= 1'h0;
		else if (_0011_)
			\mchip.row_sel[6].col_sel[4].tile_state.state  <= _0215_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[3].tile_state.state_locked  <= 1'h0;
		else if (_0196_)
			\mchip.row_sel[5].col_sel[3].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[3].tile_state.state  <= 1'h0;
		else if (_0020_)
			\mchip.row_sel[5].col_sel[3].tile_state.state  <= _0197_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[5].tile_state.state_locked  <= 1'h0;
		else if (_0232_)
			\mchip.row_sel[7].col_sel[5].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[5].tile_state.state  <= 1'h0;
		else if (_0002_)
			\mchip.row_sel[7].col_sel[5].tile_state.state  <= _0233_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[5].tile_state.state_locked  <= 1'h0;
		else if (_0184_)
			\mchip.row_sel[4].col_sel[5].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[5].tile_state.state  <= 1'h0;
		else if (_0026_)
			\mchip.row_sel[4].col_sel[5].tile_state.state  <= _0185_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[6].tile_state.state_locked  <= 1'h0;
		else if (_0122_)
			\mchip.row_sel[0].col_sel[6].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[6].tile_state.state  <= 1'h0;
		else if (_0057_)
			\mchip.row_sel[0].col_sel[6].tile_state.state  <= _0123_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[1].tile_state.state_locked  <= 1'h0;
		else if (_0144_)
			\mchip.row_sel[2].col_sel[1].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[1].tile_state.state  <= 1'h0;
		else if (_0046_)
			\mchip.row_sel[2].col_sel[1].tile_state.state  <= _0145_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[0].tile_state.state_locked  <= 1'h0;
		else if (_0158_)
			\mchip.row_sel[3].col_sel[0].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[3].col_sel[0].tile_state.state  <= 1'h0;
		else if (_0039_)
			\mchip.row_sel[3].col_sel[0].tile_state.state  <= _0159_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[7].tile_state.state_locked  <= 1'h0;
		else if (_0204_)
			\mchip.row_sel[5].col_sel[7].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[7].tile_state.state  <= 1'h0;
		else if (_0016_)
			\mchip.row_sel[5].col_sel[7].tile_state.state  <= _0205_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[6].tile_state.state_locked  <= 1'h0;
		else if (_0234_)
			\mchip.row_sel[7].col_sel[6].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[6].tile_state.state  <= 1'h0;
		else if (_0001_)
			\mchip.row_sel[7].col_sel[6].tile_state.state  <= _0235_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[5].tile_state.state_locked  <= 1'h0;
		else if (_0120_)
			\mchip.row_sel[0].col_sel[5].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[5].tile_state.state  <= 1'h0;
		else if (_0058_)
			\mchip.row_sel[0].col_sel[5].tile_state.state  <= _0121_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[5].tile_state.state_locked  <= 1'h0;
		else if (_0216_)
			\mchip.row_sel[6].col_sel[5].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[6].col_sel[5].tile_state.state  <= 1'h0;
		else if (_0010_)
			\mchip.row_sel[6].col_sel[5].tile_state.state  <= _0217_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[1].tile_state.state_locked  <= 1'h0;
		else if (_0192_)
			\mchip.row_sel[5].col_sel[1].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[5].col_sel[1].tile_state.state  <= 1'h0;
		else if (_0022_)
			\mchip.row_sel[5].col_sel[1].tile_state.state  <= _0193_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[0].tile_state.state_locked  <= 1'h0;
		else if (_0142_)
			\mchip.row_sel[2].col_sel[0].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[2].col_sel[0].tile_state.state  <= 1'h0;
		else if (_0047_)
			\mchip.row_sel[2].col_sel[0].tile_state.state  <= _0143_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[6].tile_state.state_locked  <= 1'h0;
		else if (_0186_)
			\mchip.row_sel[4].col_sel[6].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[4].col_sel[6].tile_state.state  <= 1'h0;
		else if (_0025_)
			\mchip.row_sel[4].col_sel[6].tile_state.state  <= _0187_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[4].tile_state.state_locked  <= 1'h0;
		else if (_0118_)
			\mchip.row_sel[0].col_sel[4].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[4].tile_state.state  <= 1'h0;
		else if (_0059_)
			\mchip.row_sel[0].col_sel[4].tile_state.state  <= _0119_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[7].tile_state.state_locked  <= 1'h0;
		else if (_0236_)
			\mchip.row_sel[7].col_sel[7].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[7].col_sel[7].tile_state.state  <= 1'h0;
		else if (_0000_)
			\mchip.row_sel[7].col_sel[7].tile_state.state  <= _0237_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[3].tile_state.state_locked  <= 1'h0;
		else if (_0116_)
			\mchip.row_sel[0].col_sel[3].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[3].tile_state.state  <= 1'h0;
		else if (_0060_)
			\mchip.row_sel[0].col_sel[3].tile_state.state  <= _0117_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[2].tile_state.state_locked  <= 1'h0;
		else if (_0114_)
			\mchip.row_sel[0].col_sel[2].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[2].tile_state.state  <= 1'h0;
		else if (_0061_)
			\mchip.row_sel[0].col_sel[2].tile_state.state  <= _0115_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[1].tile_state.state_locked  <= 1'h0;
		else if (_0112_)
			\mchip.row_sel[0].col_sel[1].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[1].tile_state.state  <= 1'h0;
		else if (_0062_)
			\mchip.row_sel[0].col_sel[1].tile_state.state  <= _0113_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[0].tile_state.state_locked  <= 1'h0;
		else if (_0110_)
			\mchip.row_sel[0].col_sel[0].tile_state.state_locked  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.row_sel[0].col_sel[0].tile_state.state  <= 1'h0;
		else if (_0063_)
			\mchip.row_sel[0].col_sel[0].tile_state.state  <= _0111_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.vsync  <= 1'h1;
		else if (!_0252_)
			\mchip.vga.vsync  <= _0251_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.hsync  <= 1'h1;
		else
			\mchip.vga.hsync  <= _0240_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [0] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [0] <= _0241_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [1] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [1] <= _0242_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [2] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [2] <= _0243_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [3] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [3] <= _0244_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [4] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [4] <= _0245_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [5] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [5] <= _0246_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [6] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [6] <= _0247_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [7] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [7] <= _0248_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [8] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [8] <= _0249_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.vga.v_idx [9] <= 1'h0;
		else if (!_0252_)
			\mchip.vga.v_idx [9] <= _0250_;
	always @(posedge io_in[12])
		if (_0069_)
			\mchip.vga.refresh  <= 1'h0;
		else
			\mchip.vga.refresh  <= _0238_;
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [0] <= 1'h0;
		else
			\mchip.vga.h_idx [0] <= _2115_[0];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [1] <= 1'h0;
		else
			\mchip.vga.h_idx [1] <= _2116_[1];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [2] <= 1'h0;
		else
			\mchip.vga.h_idx [2] <= _2116_[2];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [3] <= 1'h0;
		else
			\mchip.vga.h_idx [3] <= _2116_[3];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [4] <= 1'h0;
		else
			\mchip.vga.h_idx [4] <= _2116_[4];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [5] <= 1'h0;
		else
			\mchip.vga.h_idx [5] <= _2116_[5];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [6] <= 1'h0;
		else
			\mchip.vga.h_idx [6] <= _2116_[6];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [7] <= 1'h0;
		else
			\mchip.vga.h_idx [7] <= _2116_[7];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [8] <= 1'h0;
		else
			\mchip.vga.h_idx [8] <= _2116_[8];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.vga.h_idx [9] <= 1'h0;
		else
			\mchip.vga.h_idx [9] <= _2116_[9];
	always @(posedge io_in[12])
		if (_0067_)
			\mchip.vga.frame_end  <= 1'h0;
		else
			\mchip.vga.frame_end  <= _0239_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.fsm_state  <= 1'h0;
		else if (_0066_)
			\mchip.fsm_state  <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.focus_row [0] <= 1'h0;
		else if (_0065_)
			\mchip.focus_row [0] <= _0107_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.focus_row [1] <= 1'h0;
		else if (_0065_)
			\mchip.focus_row [1] <= _0108_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.focus_row [2] <= 1'h0;
		else if (_0065_)
			\mchip.focus_row [2] <= _0109_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.focus_col [0] <= 1'h0;
		else if (_0103_)
			\mchip.focus_col [0] <= _0104_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.focus_col [1] <= 1'h0;
		else if (_0103_)
			\mchip.focus_col [1] <= _0105_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.focus_col [2] <= 1'h0;
		else if (_0103_)
			\mchip.focus_col [2] <= _0106_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.lock_state  <= 1'h0;
		else if (_0064_)
			\mchip.lock_state  <= _0070_;
	always @(posedge io_in[12]) \mchip.btn3_tmp  <= io_in[0];
	always @(posedge io_in[12]) \mchip.btn3_sync  <= \mchip.btn3_tmp ;
	always @(posedge io_in[12]) \mchip.btn4_tmp  <= io_in[1];
	always @(posedge io_in[12]) \mchip.btn4_sync  <= \mchip.btn4_tmp ;
	assign _2115_[9:1] = 9'h000;
	assign _2116_[0] = _2115_[0];
	assign io_out = {5'h00, \mchip.gn16 , 2'h0, \mchip.gp23 , 3'h0, \mchip.vga.hsync , \mchip.vga.vsync };
	assign \mchip.COLS  = 32'd640;
	assign \mchip.ROWS  = 32'd480;
	assign \mchip.TILE_COLS  = 32'd8;
	assign \mchip.TILE_HEIGHT  = 32'd50;
	assign \mchip.TILE_ROWS  = 32'd8;
	assign \mchip.TILE_WIDTH  = 32'd50;
	assign \mchip.blue  = 3'h0;
	assign \mchip.bottom  = 640'h63d8f63d8f63d8f63d8f5755d5755d5755d5755d4ad2b4ad2b4ad2b4ad2b3e4f93e4f93e4f93e4f931cc731cc731cc731cc72549525495254952549518c6318c6318c6318c630c4310c4310c4310c431;
	assign \mchip.btn  = {io_in[3:0], 3'h0};
	assign \mchip.clock  = io_in[12];
	assign \mchip.frame_end  = \mchip.vga.frame_end ;
	assign \mchip.gn14  = 1'h0;
	assign \mchip.gn15  = 1'h0;
	assign \mchip.gn17  = 1'h0;
	assign \mchip.gn21  = 1'h0;
	assign \mchip.gn22  = 1'h0;
	assign \mchip.gn23  = 1'h0;
	assign \mchip.gn24  = 1'h0;
	assign \mchip.gp16  = \mchip.vga.vsync ;
	assign \mchip.gp17  = \mchip.vga.hsync ;
	assign \mchip.gp21  = 1'h0;
	assign \mchip.gp22  = 1'h0;
	assign \mchip.gp24  = 1'h0;
	assign \mchip.green  = 3'h0;
	assign \mchip.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.hsync  = \mchip.vga.hsync ;
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {3'h0, \mchip.gn16 , 2'h0, \mchip.gp23 , 3'h0, \mchip.vga.hsync , \mchip.vga.vsync };
	assign \mchip.left  = 640'h5792c3e8c8258640c8005792c3e8c8258640c8005792c3e8c8258640c8005792c3e8c8258640c8005792c3e8c8258640c8005792c3e8c8258640c8005792c3e8c8258640c8005792c3e8c8258640c800;
	assign \mchip.red  = 3'h0;
	assign \mchip.refresh  = \mchip.vga.refresh ;
	assign \mchip.reset  = io_in[13];
	assign \mchip.right  = 640'h63d5d4acf931c9518c3163d5d4acf931c9518c3163d5d4acf931c9518c3163d5d4acf931c9518c3163d5d4acf931c9518c3163d5d4acf931c9518c3163d5d4acf931c9518c3163d5d4acf931c9518c31;
	assign \mchip.row_sel[0].col_sel[0].tile.bottom  = 10'h031;
	assign \mchip.row_sel[0].col_sel[0].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[0].col_sel[0].tile.left  = 10'h000;
	assign \mchip.row_sel[0].col_sel[0].tile.right  = 10'h031;
	assign \mchip.row_sel[0].col_sel[0].tile.top  = 10'h000;
	assign \mchip.row_sel[0].col_sel[0].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[0].col_sel[0].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[0].col_sel[0].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[0].col_sel[0].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[0].col_sel[0].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[0].col_sel[0].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[0].col_sel[0].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[0].col_sel[0].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[0].col_sel[0].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[0].col_sel[1].tile.bottom  = 10'h031;
	assign \mchip.row_sel[0].col_sel[1].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[0].col_sel[1].tile.left  = 10'h032;
	assign \mchip.row_sel[0].col_sel[1].tile.right  = 10'h063;
	assign \mchip.row_sel[0].col_sel[1].tile.top  = 10'h000;
	assign \mchip.row_sel[0].col_sel[1].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[0].col_sel[1].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[0].col_sel[1].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[0].col_sel[1].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[0].col_sel[1].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[0].col_sel[1].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[0].col_sel[1].tile_state.neighbors_vert  = {\mchip.row_sel[1].col_sel[1].tile_state.state , 1'h0};
	assign \mchip.row_sel[0].col_sel[1].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[0].col_sel[1].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[0].col_sel[1].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[0].col_sel[2].tile.bottom  = 10'h031;
	assign \mchip.row_sel[0].col_sel[2].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[0].col_sel[2].tile.left  = 10'h064;
	assign \mchip.row_sel[0].col_sel[2].tile.right  = 10'h095;
	assign \mchip.row_sel[0].col_sel[2].tile.top  = 10'h000;
	assign \mchip.row_sel[0].col_sel[2].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[0].col_sel[2].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[0].col_sel[2].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[0].col_sel[2].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[0].col_sel[2].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[0].col_sel[2].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[0].col_sel[2].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[0].col_sel[2].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[0].col_sel[2].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[0].col_sel[3].tile.bottom  = 10'h031;
	assign \mchip.row_sel[0].col_sel[3].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[0].col_sel[3].tile.left  = 10'h096;
	assign \mchip.row_sel[0].col_sel[3].tile.right  = 10'h0c7;
	assign \mchip.row_sel[0].col_sel[3].tile.top  = 10'h000;
	assign \mchip.row_sel[0].col_sel[3].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[0].col_sel[3].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[0].col_sel[3].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[0].col_sel[3].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[0].col_sel[3].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[0].col_sel[3].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[0].col_sel[3].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[0].col_sel[3].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[0].col_sel[3].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[0].col_sel[4].tile.bottom  = 10'h031;
	assign \mchip.row_sel[0].col_sel[4].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[0].col_sel[4].tile.left  = 10'h0c8;
	assign \mchip.row_sel[0].col_sel[4].tile.right  = 10'h0f9;
	assign \mchip.row_sel[0].col_sel[4].tile.top  = 10'h000;
	assign \mchip.row_sel[0].col_sel[4].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[0].col_sel[4].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[0].col_sel[4].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[0].col_sel[4].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[0].col_sel[4].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[0].col_sel[4].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[0].col_sel[4].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[0].col_sel[4].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[0].col_sel[4].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[0].col_sel[5].tile.bottom  = 10'h031;
	assign \mchip.row_sel[0].col_sel[5].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[0].col_sel[5].tile.left  = 10'h0fa;
	assign \mchip.row_sel[0].col_sel[5].tile.right  = 10'h12b;
	assign \mchip.row_sel[0].col_sel[5].tile.top  = 10'h000;
	assign \mchip.row_sel[0].col_sel[5].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[0].col_sel[5].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[0].col_sel[5].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[0].col_sel[5].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[0].col_sel[5].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[0].col_sel[5].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[0].col_sel[5].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[0].col_sel[5].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[0].col_sel[5].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[0].col_sel[6].tile.bottom  = 10'h031;
	assign \mchip.row_sel[0].col_sel[6].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[0].col_sel[6].tile.left  = 10'h12c;
	assign \mchip.row_sel[0].col_sel[6].tile.right  = 10'h15d;
	assign \mchip.row_sel[0].col_sel[6].tile.top  = 10'h000;
	assign \mchip.row_sel[0].col_sel[6].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[0].col_sel[6].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[0].col_sel[6].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[0].col_sel[6].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[0].col_sel[6].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[0].col_sel[6].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[0].col_sel[6].tile_state.neighbors_vert  = {\mchip.row_sel[1].col_sel[6].tile_state.state , 1'h0};
	assign \mchip.row_sel[0].col_sel[6].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[0].col_sel[6].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[0].col_sel[6].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[0].col_sel[7].tile.bottom  = 10'h031;
	assign \mchip.row_sel[0].col_sel[7].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[0].col_sel[7].tile.left  = 10'h15e;
	assign \mchip.row_sel[0].col_sel[7].tile.right  = 10'h18f;
	assign \mchip.row_sel[0].col_sel[7].tile.top  = 10'h000;
	assign \mchip.row_sel[0].col_sel[7].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[0].col_sel[7].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[0].col_sel[7].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[0].col_sel[7].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[0].col_sel[7].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[0].col_sel[7].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[0].col_sel[7].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[0].col_sel[7].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[0].col_sel[7].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[1].col_sel[0].tile.bottom  = 10'h063;
	assign \mchip.row_sel[1].col_sel[0].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[1].col_sel[0].tile.left  = 10'h000;
	assign \mchip.row_sel[1].col_sel[0].tile.right  = 10'h031;
	assign \mchip.row_sel[1].col_sel[0].tile.top  = 10'h032;
	assign \mchip.row_sel[1].col_sel[0].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[1].col_sel[0].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[1].col_sel[0].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[1].col_sel[0].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[1].col_sel[0].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[1].col_sel[0].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[1].col_sel[0].tile_state.neighbors_hori  = {\mchip.row_sel[1].col_sel[1].tile_state.state , 1'h0};
	assign \mchip.row_sel[1].col_sel[0].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[1].col_sel[0].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[1].col_sel[0].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[1].col_sel[1].tile.bottom  = 10'h063;
	assign \mchip.row_sel[1].col_sel[1].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[1].col_sel[1].tile.left  = 10'h032;
	assign \mchip.row_sel[1].col_sel[1].tile.right  = 10'h063;
	assign \mchip.row_sel[1].col_sel[1].tile.top  = 10'h032;
	assign \mchip.row_sel[1].col_sel[1].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[1].col_sel[1].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[1].col_sel[1].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[1].col_sel[1].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[1].col_sel[1].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[1].col_sel[1].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[1].col_sel[1].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[1].col_sel[1].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[1].col_sel[1].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[1].col_sel[2].tile.bottom  = 10'h063;
	assign \mchip.row_sel[1].col_sel[2].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[1].col_sel[2].tile.left  = 10'h064;
	assign \mchip.row_sel[1].col_sel[2].tile.right  = 10'h095;
	assign \mchip.row_sel[1].col_sel[2].tile.top  = 10'h032;
	assign \mchip.row_sel[1].col_sel[2].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[1].col_sel[2].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[1].col_sel[2].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[1].col_sel[2].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[1].col_sel[2].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[1].col_sel[2].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[1].col_sel[2].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[1].col_sel[2].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[1].col_sel[2].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[1].col_sel[3].tile.bottom  = 10'h063;
	assign \mchip.row_sel[1].col_sel[3].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[1].col_sel[3].tile.left  = 10'h096;
	assign \mchip.row_sel[1].col_sel[3].tile.right  = 10'h0c7;
	assign \mchip.row_sel[1].col_sel[3].tile.top  = 10'h032;
	assign \mchip.row_sel[1].col_sel[3].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[1].col_sel[3].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[1].col_sel[3].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[1].col_sel[3].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[1].col_sel[3].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[1].col_sel[3].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[1].col_sel[3].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[1].col_sel[3].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[1].col_sel[3].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[1].col_sel[4].tile.bottom  = 10'h063;
	assign \mchip.row_sel[1].col_sel[4].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[1].col_sel[4].tile.left  = 10'h0c8;
	assign \mchip.row_sel[1].col_sel[4].tile.right  = 10'h0f9;
	assign \mchip.row_sel[1].col_sel[4].tile.top  = 10'h032;
	assign \mchip.row_sel[1].col_sel[4].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[1].col_sel[4].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[1].col_sel[4].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[1].col_sel[4].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[1].col_sel[4].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[1].col_sel[4].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[1].col_sel[4].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[1].col_sel[4].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[1].col_sel[4].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[1].col_sel[5].tile.bottom  = 10'h063;
	assign \mchip.row_sel[1].col_sel[5].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[1].col_sel[5].tile.left  = 10'h0fa;
	assign \mchip.row_sel[1].col_sel[5].tile.right  = 10'h12b;
	assign \mchip.row_sel[1].col_sel[5].tile.top  = 10'h032;
	assign \mchip.row_sel[1].col_sel[5].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[1].col_sel[5].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[1].col_sel[5].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[1].col_sel[5].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[1].col_sel[5].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[1].col_sel[5].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[1].col_sel[5].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[1].col_sel[5].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[1].col_sel[5].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[1].col_sel[6].tile.bottom  = 10'h063;
	assign \mchip.row_sel[1].col_sel[6].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[1].col_sel[6].tile.left  = 10'h12c;
	assign \mchip.row_sel[1].col_sel[6].tile.right  = 10'h15d;
	assign \mchip.row_sel[1].col_sel[6].tile.top  = 10'h032;
	assign \mchip.row_sel[1].col_sel[6].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[1].col_sel[6].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[1].col_sel[6].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[1].col_sel[6].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[1].col_sel[6].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[1].col_sel[6].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[1].col_sel[6].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[1].col_sel[6].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[1].col_sel[6].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[1].col_sel[7].tile.bottom  = 10'h063;
	assign \mchip.row_sel[1].col_sel[7].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[1].col_sel[7].tile.left  = 10'h15e;
	assign \mchip.row_sel[1].col_sel[7].tile.right  = 10'h18f;
	assign \mchip.row_sel[1].col_sel[7].tile.top  = 10'h032;
	assign \mchip.row_sel[1].col_sel[7].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[1].col_sel[7].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[1].col_sel[7].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[1].col_sel[7].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[1].col_sel[7].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[1].col_sel[7].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[1].col_sel[7].tile_state.neighbors_hori  = {\mchip.row_sel[1].col_sel[6].tile_state.state , 1'h0};
	assign \mchip.row_sel[1].col_sel[7].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[1].col_sel[7].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[1].col_sel[7].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[2].col_sel[0].tile.bottom  = 10'h095;
	assign \mchip.row_sel[2].col_sel[0].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[2].col_sel[0].tile.left  = 10'h000;
	assign \mchip.row_sel[2].col_sel[0].tile.right  = 10'h031;
	assign \mchip.row_sel[2].col_sel[0].tile.top  = 10'h064;
	assign \mchip.row_sel[2].col_sel[0].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[2].col_sel[0].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[2].col_sel[0].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[2].col_sel[0].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[2].col_sel[0].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[2].col_sel[0].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[2].col_sel[0].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[2].col_sel[0].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[2].col_sel[0].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[2].col_sel[1].tile.bottom  = 10'h095;
	assign \mchip.row_sel[2].col_sel[1].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[2].col_sel[1].tile.left  = 10'h032;
	assign \mchip.row_sel[2].col_sel[1].tile.right  = 10'h063;
	assign \mchip.row_sel[2].col_sel[1].tile.top  = 10'h064;
	assign \mchip.row_sel[2].col_sel[1].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[2].col_sel[1].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[2].col_sel[1].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[2].col_sel[1].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[2].col_sel[1].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[2].col_sel[1].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[2].col_sel[1].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[2].col_sel[1].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[2].col_sel[1].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[2].col_sel[2].tile.bottom  = 10'h095;
	assign \mchip.row_sel[2].col_sel[2].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[2].col_sel[2].tile.left  = 10'h064;
	assign \mchip.row_sel[2].col_sel[2].tile.right  = 10'h095;
	assign \mchip.row_sel[2].col_sel[2].tile.top  = 10'h064;
	assign \mchip.row_sel[2].col_sel[2].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[2].col_sel[2].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[2].col_sel[2].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[2].col_sel[2].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[2].col_sel[2].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[2].col_sel[2].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[2].col_sel[2].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[2].col_sel[2].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[2].col_sel[2].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[2].col_sel[3].tile.bottom  = 10'h095;
	assign \mchip.row_sel[2].col_sel[3].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[2].col_sel[3].tile.left  = 10'h096;
	assign \mchip.row_sel[2].col_sel[3].tile.right  = 10'h0c7;
	assign \mchip.row_sel[2].col_sel[3].tile.top  = 10'h064;
	assign \mchip.row_sel[2].col_sel[3].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[2].col_sel[3].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[2].col_sel[3].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[2].col_sel[3].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[2].col_sel[3].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[2].col_sel[3].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[2].col_sel[3].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[2].col_sel[3].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[2].col_sel[3].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[2].col_sel[4].tile.bottom  = 10'h095;
	assign \mchip.row_sel[2].col_sel[4].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[2].col_sel[4].tile.left  = 10'h0c8;
	assign \mchip.row_sel[2].col_sel[4].tile.right  = 10'h0f9;
	assign \mchip.row_sel[2].col_sel[4].tile.top  = 10'h064;
	assign \mchip.row_sel[2].col_sel[4].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[2].col_sel[4].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[2].col_sel[4].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[2].col_sel[4].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[2].col_sel[4].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[2].col_sel[4].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[2].col_sel[4].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[2].col_sel[4].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[2].col_sel[4].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[2].col_sel[5].tile.bottom  = 10'h095;
	assign \mchip.row_sel[2].col_sel[5].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[2].col_sel[5].tile.left  = 10'h0fa;
	assign \mchip.row_sel[2].col_sel[5].tile.right  = 10'h12b;
	assign \mchip.row_sel[2].col_sel[5].tile.top  = 10'h064;
	assign \mchip.row_sel[2].col_sel[5].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[2].col_sel[5].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[2].col_sel[5].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[2].col_sel[5].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[2].col_sel[5].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[2].col_sel[5].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[2].col_sel[5].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[2].col_sel[5].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[2].col_sel[5].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[2].col_sel[6].tile.bottom  = 10'h095;
	assign \mchip.row_sel[2].col_sel[6].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[2].col_sel[6].tile.left  = 10'h12c;
	assign \mchip.row_sel[2].col_sel[6].tile.right  = 10'h15d;
	assign \mchip.row_sel[2].col_sel[6].tile.top  = 10'h064;
	assign \mchip.row_sel[2].col_sel[6].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[2].col_sel[6].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[2].col_sel[6].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[2].col_sel[6].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[2].col_sel[6].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[2].col_sel[6].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[2].col_sel[6].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[2].col_sel[6].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[2].col_sel[6].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[2].col_sel[7].tile.bottom  = 10'h095;
	assign \mchip.row_sel[2].col_sel[7].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[2].col_sel[7].tile.left  = 10'h15e;
	assign \mchip.row_sel[2].col_sel[7].tile.right  = 10'h18f;
	assign \mchip.row_sel[2].col_sel[7].tile.top  = 10'h064;
	assign \mchip.row_sel[2].col_sel[7].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[2].col_sel[7].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[2].col_sel[7].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[2].col_sel[7].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[2].col_sel[7].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[2].col_sel[7].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[2].col_sel[7].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[2].col_sel[7].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[2].col_sel[7].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[3].col_sel[0].tile.bottom  = 10'h0c7;
	assign \mchip.row_sel[3].col_sel[0].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[3].col_sel[0].tile.left  = 10'h000;
	assign \mchip.row_sel[3].col_sel[0].tile.right  = 10'h031;
	assign \mchip.row_sel[3].col_sel[0].tile.top  = 10'h096;
	assign \mchip.row_sel[3].col_sel[0].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[3].col_sel[0].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[3].col_sel[0].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[3].col_sel[0].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[3].col_sel[0].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[3].col_sel[0].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[3].col_sel[0].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[3].col_sel[0].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[3].col_sel[0].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[3].col_sel[1].tile.bottom  = 10'h0c7;
	assign \mchip.row_sel[3].col_sel[1].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[3].col_sel[1].tile.left  = 10'h032;
	assign \mchip.row_sel[3].col_sel[1].tile.right  = 10'h063;
	assign \mchip.row_sel[3].col_sel[1].tile.top  = 10'h096;
	assign \mchip.row_sel[3].col_sel[1].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[3].col_sel[1].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[3].col_sel[1].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[3].col_sel[1].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[3].col_sel[1].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[3].col_sel[1].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[3].col_sel[1].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[3].col_sel[1].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[3].col_sel[1].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[3].col_sel[2].tile.bottom  = 10'h0c7;
	assign \mchip.row_sel[3].col_sel[2].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[3].col_sel[2].tile.left  = 10'h064;
	assign \mchip.row_sel[3].col_sel[2].tile.right  = 10'h095;
	assign \mchip.row_sel[3].col_sel[2].tile.top  = 10'h096;
	assign \mchip.row_sel[3].col_sel[2].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[3].col_sel[2].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[3].col_sel[2].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[3].col_sel[2].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[3].col_sel[2].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[3].col_sel[2].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[3].col_sel[2].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[3].col_sel[2].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[3].col_sel[2].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[3].col_sel[3].tile.bottom  = 10'h0c7;
	assign \mchip.row_sel[3].col_sel[3].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[3].col_sel[3].tile.left  = 10'h096;
	assign \mchip.row_sel[3].col_sel[3].tile.right  = 10'h0c7;
	assign \mchip.row_sel[3].col_sel[3].tile.top  = 10'h096;
	assign \mchip.row_sel[3].col_sel[3].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[3].col_sel[3].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[3].col_sel[3].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[3].col_sel[3].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[3].col_sel[3].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[3].col_sel[3].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[3].col_sel[3].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[3].col_sel[3].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[3].col_sel[3].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[3].col_sel[4].tile.bottom  = 10'h0c7;
	assign \mchip.row_sel[3].col_sel[4].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[3].col_sel[4].tile.left  = 10'h0c8;
	assign \mchip.row_sel[3].col_sel[4].tile.right  = 10'h0f9;
	assign \mchip.row_sel[3].col_sel[4].tile.top  = 10'h096;
	assign \mchip.row_sel[3].col_sel[4].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[3].col_sel[4].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[3].col_sel[4].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[3].col_sel[4].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[3].col_sel[4].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[3].col_sel[4].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[3].col_sel[4].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[3].col_sel[4].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[3].col_sel[4].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[3].col_sel[5].tile.bottom  = 10'h0c7;
	assign \mchip.row_sel[3].col_sel[5].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[3].col_sel[5].tile.left  = 10'h0fa;
	assign \mchip.row_sel[3].col_sel[5].tile.right  = 10'h12b;
	assign \mchip.row_sel[3].col_sel[5].tile.top  = 10'h096;
	assign \mchip.row_sel[3].col_sel[5].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[3].col_sel[5].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[3].col_sel[5].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[3].col_sel[5].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[3].col_sel[5].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[3].col_sel[5].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[3].col_sel[5].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[3].col_sel[5].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[3].col_sel[5].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[3].col_sel[6].tile.bottom  = 10'h0c7;
	assign \mchip.row_sel[3].col_sel[6].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[3].col_sel[6].tile.left  = 10'h12c;
	assign \mchip.row_sel[3].col_sel[6].tile.right  = 10'h15d;
	assign \mchip.row_sel[3].col_sel[6].tile.top  = 10'h096;
	assign \mchip.row_sel[3].col_sel[6].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[3].col_sel[6].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[3].col_sel[6].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[3].col_sel[6].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[3].col_sel[6].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[3].col_sel[6].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[3].col_sel[6].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[3].col_sel[6].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[3].col_sel[6].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[3].col_sel[7].tile.bottom  = 10'h0c7;
	assign \mchip.row_sel[3].col_sel[7].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[3].col_sel[7].tile.left  = 10'h15e;
	assign \mchip.row_sel[3].col_sel[7].tile.right  = 10'h18f;
	assign \mchip.row_sel[3].col_sel[7].tile.top  = 10'h096;
	assign \mchip.row_sel[3].col_sel[7].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[3].col_sel[7].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[3].col_sel[7].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[3].col_sel[7].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[3].col_sel[7].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[3].col_sel[7].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[3].col_sel[7].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[3].col_sel[7].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[3].col_sel[7].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[4].col_sel[0].tile.bottom  = 10'h0f9;
	assign \mchip.row_sel[4].col_sel[0].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[4].col_sel[0].tile.left  = 10'h000;
	assign \mchip.row_sel[4].col_sel[0].tile.right  = 10'h031;
	assign \mchip.row_sel[4].col_sel[0].tile.top  = 10'h0c8;
	assign \mchip.row_sel[4].col_sel[0].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[4].col_sel[0].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[4].col_sel[0].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[4].col_sel[0].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[4].col_sel[0].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[4].col_sel[0].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[4].col_sel[0].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[4].col_sel[0].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[4].col_sel[0].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[4].col_sel[1].tile.bottom  = 10'h0f9;
	assign \mchip.row_sel[4].col_sel[1].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[4].col_sel[1].tile.left  = 10'h032;
	assign \mchip.row_sel[4].col_sel[1].tile.right  = 10'h063;
	assign \mchip.row_sel[4].col_sel[1].tile.top  = 10'h0c8;
	assign \mchip.row_sel[4].col_sel[1].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[4].col_sel[1].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[4].col_sel[1].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[4].col_sel[1].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[4].col_sel[1].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[4].col_sel[1].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[4].col_sel[1].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[4].col_sel[1].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[4].col_sel[1].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[4].col_sel[2].tile.bottom  = 10'h0f9;
	assign \mchip.row_sel[4].col_sel[2].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[4].col_sel[2].tile.left  = 10'h064;
	assign \mchip.row_sel[4].col_sel[2].tile.right  = 10'h095;
	assign \mchip.row_sel[4].col_sel[2].tile.top  = 10'h0c8;
	assign \mchip.row_sel[4].col_sel[2].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[4].col_sel[2].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[4].col_sel[2].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[4].col_sel[2].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[4].col_sel[2].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[4].col_sel[2].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[4].col_sel[2].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[4].col_sel[2].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[4].col_sel[2].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[4].col_sel[3].tile.bottom  = 10'h0f9;
	assign \mchip.row_sel[4].col_sel[3].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[4].col_sel[3].tile.left  = 10'h096;
	assign \mchip.row_sel[4].col_sel[3].tile.right  = 10'h0c7;
	assign \mchip.row_sel[4].col_sel[3].tile.top  = 10'h0c8;
	assign \mchip.row_sel[4].col_sel[3].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[4].col_sel[3].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[4].col_sel[3].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[4].col_sel[3].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[4].col_sel[3].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[4].col_sel[3].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[4].col_sel[3].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[4].col_sel[3].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[4].col_sel[3].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[4].col_sel[4].tile.bottom  = 10'h0f9;
	assign \mchip.row_sel[4].col_sel[4].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[4].col_sel[4].tile.left  = 10'h0c8;
	assign \mchip.row_sel[4].col_sel[4].tile.right  = 10'h0f9;
	assign \mchip.row_sel[4].col_sel[4].tile.top  = 10'h0c8;
	assign \mchip.row_sel[4].col_sel[4].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[4].col_sel[4].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[4].col_sel[4].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[4].col_sel[4].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[4].col_sel[4].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[4].col_sel[4].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[4].col_sel[4].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[4].col_sel[4].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[4].col_sel[4].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[4].col_sel[5].tile.bottom  = 10'h0f9;
	assign \mchip.row_sel[4].col_sel[5].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[4].col_sel[5].tile.left  = 10'h0fa;
	assign \mchip.row_sel[4].col_sel[5].tile.right  = 10'h12b;
	assign \mchip.row_sel[4].col_sel[5].tile.top  = 10'h0c8;
	assign \mchip.row_sel[4].col_sel[5].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[4].col_sel[5].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[4].col_sel[5].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[4].col_sel[5].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[4].col_sel[5].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[4].col_sel[5].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[4].col_sel[5].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[4].col_sel[5].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[4].col_sel[5].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[4].col_sel[6].tile.bottom  = 10'h0f9;
	assign \mchip.row_sel[4].col_sel[6].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[4].col_sel[6].tile.left  = 10'h12c;
	assign \mchip.row_sel[4].col_sel[6].tile.right  = 10'h15d;
	assign \mchip.row_sel[4].col_sel[6].tile.top  = 10'h0c8;
	assign \mchip.row_sel[4].col_sel[6].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[4].col_sel[6].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[4].col_sel[6].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[4].col_sel[6].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[4].col_sel[6].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[4].col_sel[6].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[4].col_sel[6].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[4].col_sel[6].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[4].col_sel[6].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[4].col_sel[7].tile.bottom  = 10'h0f9;
	assign \mchip.row_sel[4].col_sel[7].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[4].col_sel[7].tile.left  = 10'h15e;
	assign \mchip.row_sel[4].col_sel[7].tile.right  = 10'h18f;
	assign \mchip.row_sel[4].col_sel[7].tile.top  = 10'h0c8;
	assign \mchip.row_sel[4].col_sel[7].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[4].col_sel[7].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[4].col_sel[7].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[4].col_sel[7].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[4].col_sel[7].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[4].col_sel[7].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[4].col_sel[7].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[4].col_sel[7].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[4].col_sel[7].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[5].col_sel[0].tile.bottom  = 10'h12b;
	assign \mchip.row_sel[5].col_sel[0].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[5].col_sel[0].tile.left  = 10'h000;
	assign \mchip.row_sel[5].col_sel[0].tile.right  = 10'h031;
	assign \mchip.row_sel[5].col_sel[0].tile.top  = 10'h0fa;
	assign \mchip.row_sel[5].col_sel[0].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[5].col_sel[0].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[5].col_sel[0].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[5].col_sel[0].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[5].col_sel[0].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[5].col_sel[0].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[5].col_sel[0].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[5].col_sel[0].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[5].col_sel[0].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[5].col_sel[1].tile.bottom  = 10'h12b;
	assign \mchip.row_sel[5].col_sel[1].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[5].col_sel[1].tile.left  = 10'h032;
	assign \mchip.row_sel[5].col_sel[1].tile.right  = 10'h063;
	assign \mchip.row_sel[5].col_sel[1].tile.top  = 10'h0fa;
	assign \mchip.row_sel[5].col_sel[1].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[5].col_sel[1].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[5].col_sel[1].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[5].col_sel[1].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[5].col_sel[1].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[5].col_sel[1].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[5].col_sel[1].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[5].col_sel[1].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[5].col_sel[1].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[5].col_sel[2].tile.bottom  = 10'h12b;
	assign \mchip.row_sel[5].col_sel[2].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[5].col_sel[2].tile.left  = 10'h064;
	assign \mchip.row_sel[5].col_sel[2].tile.right  = 10'h095;
	assign \mchip.row_sel[5].col_sel[2].tile.top  = 10'h0fa;
	assign \mchip.row_sel[5].col_sel[2].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[5].col_sel[2].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[5].col_sel[2].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[5].col_sel[2].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[5].col_sel[2].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[5].col_sel[2].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[5].col_sel[2].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[5].col_sel[2].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[5].col_sel[2].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[5].col_sel[3].tile.bottom  = 10'h12b;
	assign \mchip.row_sel[5].col_sel[3].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[5].col_sel[3].tile.left  = 10'h096;
	assign \mchip.row_sel[5].col_sel[3].tile.right  = 10'h0c7;
	assign \mchip.row_sel[5].col_sel[3].tile.top  = 10'h0fa;
	assign \mchip.row_sel[5].col_sel[3].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[5].col_sel[3].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[5].col_sel[3].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[5].col_sel[3].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[5].col_sel[3].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[5].col_sel[3].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[5].col_sel[3].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[5].col_sel[3].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[5].col_sel[3].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[5].col_sel[4].tile.bottom  = 10'h12b;
	assign \mchip.row_sel[5].col_sel[4].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[5].col_sel[4].tile.left  = 10'h0c8;
	assign \mchip.row_sel[5].col_sel[4].tile.right  = 10'h0f9;
	assign \mchip.row_sel[5].col_sel[4].tile.top  = 10'h0fa;
	assign \mchip.row_sel[5].col_sel[4].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[5].col_sel[4].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[5].col_sel[4].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[5].col_sel[4].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[5].col_sel[4].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[5].col_sel[4].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[5].col_sel[4].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[5].col_sel[4].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[5].col_sel[4].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[5].col_sel[5].tile.bottom  = 10'h12b;
	assign \mchip.row_sel[5].col_sel[5].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[5].col_sel[5].tile.left  = 10'h0fa;
	assign \mchip.row_sel[5].col_sel[5].tile.right  = 10'h12b;
	assign \mchip.row_sel[5].col_sel[5].tile.top  = 10'h0fa;
	assign \mchip.row_sel[5].col_sel[5].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[5].col_sel[5].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[5].col_sel[5].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[5].col_sel[5].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[5].col_sel[5].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[5].col_sel[5].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[5].col_sel[5].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[5].col_sel[5].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[5].col_sel[5].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[5].col_sel[6].tile.bottom  = 10'h12b;
	assign \mchip.row_sel[5].col_sel[6].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[5].col_sel[6].tile.left  = 10'h12c;
	assign \mchip.row_sel[5].col_sel[6].tile.right  = 10'h15d;
	assign \mchip.row_sel[5].col_sel[6].tile.top  = 10'h0fa;
	assign \mchip.row_sel[5].col_sel[6].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[5].col_sel[6].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[5].col_sel[6].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[5].col_sel[6].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[5].col_sel[6].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[5].col_sel[6].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[5].col_sel[6].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[5].col_sel[6].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[5].col_sel[6].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[5].col_sel[7].tile.bottom  = 10'h12b;
	assign \mchip.row_sel[5].col_sel[7].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[5].col_sel[7].tile.left  = 10'h15e;
	assign \mchip.row_sel[5].col_sel[7].tile.right  = 10'h18f;
	assign \mchip.row_sel[5].col_sel[7].tile.top  = 10'h0fa;
	assign \mchip.row_sel[5].col_sel[7].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[5].col_sel[7].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[5].col_sel[7].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[5].col_sel[7].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[5].col_sel[7].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[5].col_sel[7].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[5].col_sel[7].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[5].col_sel[7].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[5].col_sel[7].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[6].col_sel[0].tile.bottom  = 10'h15d;
	assign \mchip.row_sel[6].col_sel[0].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[6].col_sel[0].tile.left  = 10'h000;
	assign \mchip.row_sel[6].col_sel[0].tile.right  = 10'h031;
	assign \mchip.row_sel[6].col_sel[0].tile.top  = 10'h12c;
	assign \mchip.row_sel[6].col_sel[0].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[6].col_sel[0].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[6].col_sel[0].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[6].col_sel[0].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[6].col_sel[0].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[6].col_sel[0].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[6].col_sel[0].tile_state.neighbors_hori  = {\mchip.row_sel[6].col_sel[1].tile_state.state , 1'h0};
	assign \mchip.row_sel[6].col_sel[0].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[6].col_sel[0].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[6].col_sel[0].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[6].col_sel[1].tile.bottom  = 10'h15d;
	assign \mchip.row_sel[6].col_sel[1].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[6].col_sel[1].tile.left  = 10'h032;
	assign \mchip.row_sel[6].col_sel[1].tile.right  = 10'h063;
	assign \mchip.row_sel[6].col_sel[1].tile.top  = 10'h12c;
	assign \mchip.row_sel[6].col_sel[1].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[6].col_sel[1].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[6].col_sel[1].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[6].col_sel[1].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[6].col_sel[1].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[6].col_sel[1].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[6].col_sel[1].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[6].col_sel[1].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[6].col_sel[1].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[6].col_sel[2].tile.bottom  = 10'h15d;
	assign \mchip.row_sel[6].col_sel[2].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[6].col_sel[2].tile.left  = 10'h064;
	assign \mchip.row_sel[6].col_sel[2].tile.right  = 10'h095;
	assign \mchip.row_sel[6].col_sel[2].tile.top  = 10'h12c;
	assign \mchip.row_sel[6].col_sel[2].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[6].col_sel[2].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[6].col_sel[2].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[6].col_sel[2].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[6].col_sel[2].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[6].col_sel[2].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[6].col_sel[2].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[6].col_sel[2].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[6].col_sel[2].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[6].col_sel[3].tile.bottom  = 10'h15d;
	assign \mchip.row_sel[6].col_sel[3].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[6].col_sel[3].tile.left  = 10'h096;
	assign \mchip.row_sel[6].col_sel[3].tile.right  = 10'h0c7;
	assign \mchip.row_sel[6].col_sel[3].tile.top  = 10'h12c;
	assign \mchip.row_sel[6].col_sel[3].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[6].col_sel[3].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[6].col_sel[3].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[6].col_sel[3].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[6].col_sel[3].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[6].col_sel[3].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[6].col_sel[3].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[6].col_sel[3].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[6].col_sel[3].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[6].col_sel[4].tile.bottom  = 10'h15d;
	assign \mchip.row_sel[6].col_sel[4].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[6].col_sel[4].tile.left  = 10'h0c8;
	assign \mchip.row_sel[6].col_sel[4].tile.right  = 10'h0f9;
	assign \mchip.row_sel[6].col_sel[4].tile.top  = 10'h12c;
	assign \mchip.row_sel[6].col_sel[4].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[6].col_sel[4].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[6].col_sel[4].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[6].col_sel[4].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[6].col_sel[4].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[6].col_sel[4].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[6].col_sel[4].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[6].col_sel[4].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[6].col_sel[4].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[6].col_sel[5].tile.bottom  = 10'h15d;
	assign \mchip.row_sel[6].col_sel[5].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[6].col_sel[5].tile.left  = 10'h0fa;
	assign \mchip.row_sel[6].col_sel[5].tile.right  = 10'h12b;
	assign \mchip.row_sel[6].col_sel[5].tile.top  = 10'h12c;
	assign \mchip.row_sel[6].col_sel[5].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[6].col_sel[5].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[6].col_sel[5].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[6].col_sel[5].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[6].col_sel[5].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[6].col_sel[5].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[6].col_sel[5].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[6].col_sel[5].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[6].col_sel[5].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[6].col_sel[6].tile.bottom  = 10'h15d;
	assign \mchip.row_sel[6].col_sel[6].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[6].col_sel[6].tile.left  = 10'h12c;
	assign \mchip.row_sel[6].col_sel[6].tile.right  = 10'h15d;
	assign \mchip.row_sel[6].col_sel[6].tile.top  = 10'h12c;
	assign \mchip.row_sel[6].col_sel[6].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[6].col_sel[6].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[6].col_sel[6].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[6].col_sel[6].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[6].col_sel[6].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[6].col_sel[6].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[6].col_sel[6].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[6].col_sel[6].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[6].col_sel[6].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[6].col_sel[7].tile.bottom  = 10'h15d;
	assign \mchip.row_sel[6].col_sel[7].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[6].col_sel[7].tile.left  = 10'h15e;
	assign \mchip.row_sel[6].col_sel[7].tile.right  = 10'h18f;
	assign \mchip.row_sel[6].col_sel[7].tile.top  = 10'h12c;
	assign \mchip.row_sel[6].col_sel[7].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[6].col_sel[7].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[6].col_sel[7].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[6].col_sel[7].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[6].col_sel[7].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[6].col_sel[7].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[6].col_sel[7].tile_state.neighbors_hori  = {\mchip.row_sel[6].col_sel[6].tile_state.state , 1'h0};
	assign \mchip.row_sel[6].col_sel[7].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[6].col_sel[7].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[6].col_sel[7].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[7].col_sel[0].tile.bottom  = 10'h18f;
	assign \mchip.row_sel[7].col_sel[0].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[7].col_sel[0].tile.left  = 10'h000;
	assign \mchip.row_sel[7].col_sel[0].tile.right  = 10'h031;
	assign \mchip.row_sel[7].col_sel[0].tile.top  = 10'h15e;
	assign \mchip.row_sel[7].col_sel[0].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[7].col_sel[0].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[7].col_sel[0].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[7].col_sel[0].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[7].col_sel[0].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[7].col_sel[0].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[7].col_sel[0].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[7].col_sel[0].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[7].col_sel[0].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[7].col_sel[1].tile.bottom  = 10'h18f;
	assign \mchip.row_sel[7].col_sel[1].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[7].col_sel[1].tile.left  = 10'h032;
	assign \mchip.row_sel[7].col_sel[1].tile.right  = 10'h063;
	assign \mchip.row_sel[7].col_sel[1].tile.top  = 10'h15e;
	assign \mchip.row_sel[7].col_sel[1].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[7].col_sel[1].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[7].col_sel[1].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[7].col_sel[1].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[7].col_sel[1].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[7].col_sel[1].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[7].col_sel[1].tile_state.neighbors_vert  = {\mchip.row_sel[6].col_sel[1].tile_state.state , 1'h0};
	assign \mchip.row_sel[7].col_sel[1].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[7].col_sel[1].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[7].col_sel[1].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[7].col_sel[2].tile.bottom  = 10'h18f;
	assign \mchip.row_sel[7].col_sel[2].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[7].col_sel[2].tile.left  = 10'h064;
	assign \mchip.row_sel[7].col_sel[2].tile.right  = 10'h095;
	assign \mchip.row_sel[7].col_sel[2].tile.top  = 10'h15e;
	assign \mchip.row_sel[7].col_sel[2].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[7].col_sel[2].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[7].col_sel[2].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[7].col_sel[2].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[7].col_sel[2].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[7].col_sel[2].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[7].col_sel[2].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[7].col_sel[2].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[7].col_sel[2].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[7].col_sel[3].tile.bottom  = 10'h18f;
	assign \mchip.row_sel[7].col_sel[3].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[7].col_sel[3].tile.left  = 10'h096;
	assign \mchip.row_sel[7].col_sel[3].tile.right  = 10'h0c7;
	assign \mchip.row_sel[7].col_sel[3].tile.top  = 10'h15e;
	assign \mchip.row_sel[7].col_sel[3].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[7].col_sel[3].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[7].col_sel[3].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[7].col_sel[3].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[7].col_sel[3].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[7].col_sel[3].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[7].col_sel[3].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[7].col_sel[3].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[7].col_sel[3].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[7].col_sel[4].tile.bottom  = 10'h18f;
	assign \mchip.row_sel[7].col_sel[4].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[7].col_sel[4].tile.left  = 10'h0c8;
	assign \mchip.row_sel[7].col_sel[4].tile.right  = 10'h0f9;
	assign \mchip.row_sel[7].col_sel[4].tile.top  = 10'h15e;
	assign \mchip.row_sel[7].col_sel[4].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[7].col_sel[4].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[7].col_sel[4].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[7].col_sel[4].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[7].col_sel[4].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[7].col_sel[4].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[7].col_sel[4].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[7].col_sel[4].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[7].col_sel[4].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[7].col_sel[5].tile.bottom  = 10'h18f;
	assign \mchip.row_sel[7].col_sel[5].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[7].col_sel[5].tile.left  = 10'h0fa;
	assign \mchip.row_sel[7].col_sel[5].tile.right  = 10'h12b;
	assign \mchip.row_sel[7].col_sel[5].tile.top  = 10'h15e;
	assign \mchip.row_sel[7].col_sel[5].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[7].col_sel[5].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[7].col_sel[5].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[7].col_sel[5].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[7].col_sel[5].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[7].col_sel[5].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[7].col_sel[5].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[7].col_sel[5].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[7].col_sel[5].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[7].col_sel[6].tile.bottom  = 10'h18f;
	assign \mchip.row_sel[7].col_sel[6].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[7].col_sel[6].tile.left  = 10'h12c;
	assign \mchip.row_sel[7].col_sel[6].tile.right  = 10'h15d;
	assign \mchip.row_sel[7].col_sel[6].tile.top  = 10'h15e;
	assign \mchip.row_sel[7].col_sel[6].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[7].col_sel[6].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[7].col_sel[6].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[7].col_sel[6].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[7].col_sel[6].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[7].col_sel[6].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[7].col_sel[6].tile_state.neighbors_vert  = {\mchip.row_sel[6].col_sel[6].tile_state.state , 1'h0};
	assign \mchip.row_sel[7].col_sel[6].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[7].col_sel[6].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[7].col_sel[6].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.row_sel[7].col_sel[7].tile.bottom  = 10'h18f;
	assign \mchip.row_sel[7].col_sel[7].tile.h_idx  = \mchip.vga.h_idx ;
	assign \mchip.row_sel[7].col_sel[7].tile.left  = 10'h15e;
	assign \mchip.row_sel[7].col_sel[7].tile.right  = 10'h18f;
	assign \mchip.row_sel[7].col_sel[7].tile.top  = 10'h15e;
	assign \mchip.row_sel[7].col_sel[7].tile.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.row_sel[7].col_sel[7].tile_state.clk  = io_in[12];
	assign \mchip.row_sel[7].col_sel[7].tile_state.focus_col  = \mchip.focus_col ;
	assign \mchip.row_sel[7].col_sel[7].tile_state.focus_row  = \mchip.focus_row ;
	assign \mchip.row_sel[7].col_sel[7].tile_state.fsm_state  = \mchip.fsm_state ;
	assign \mchip.row_sel[7].col_sel[7].tile_state.lock_state  = \mchip.lock_state ;
	assign \mchip.row_sel[7].col_sel[7].tile_state.refresh  = \mchip.vga.refresh ;
	assign \mchip.row_sel[7].col_sel[7].tile_state.rst  = io_in[13];
	assign \mchip.row_sel[7].col_sel[7].tile_state.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.tile_states  = {\mchip.row_sel[7].col_sel[7].tile_state.state , \mchip.row_sel[7].col_sel[6].tile_state.state , \mchip.row_sel[7].col_sel[5].tile_state.state , \mchip.row_sel[7].col_sel[4].tile_state.state , \mchip.row_sel[7].col_sel[3].tile_state.state , \mchip.row_sel[7].col_sel[2].tile_state.state , \mchip.row_sel[7].col_sel[1].tile_state.state , \mchip.row_sel[7].col_sel[0].tile_state.state , \mchip.row_sel[6].col_sel[7].tile_state.state , \mchip.row_sel[6].col_sel[6].tile_state.state , \mchip.row_sel[6].col_sel[5].tile_state.state , \mchip.row_sel[6].col_sel[4].tile_state.state , \mchip.row_sel[6].col_sel[3].tile_state.state , \mchip.row_sel[6].col_sel[2].tile_state.state , \mchip.row_sel[6].col_sel[1].tile_state.state , \mchip.row_sel[6].col_sel[0].tile_state.state , \mchip.row_sel[5].col_sel[7].tile_state.state , \mchip.row_sel[5].col_sel[6].tile_state.state , \mchip.row_sel[5].col_sel[5].tile_state.state , \mchip.row_sel[5].col_sel[4].tile_state.state , \mchip.row_sel[5].col_sel[3].tile_state.state , \mchip.row_sel[5].col_sel[2].tile_state.state , \mchip.row_sel[5].col_sel[1].tile_state.state , \mchip.row_sel[5].col_sel[0].tile_state.state , \mchip.row_sel[4].col_sel[7].tile_state.state , \mchip.row_sel[4].col_sel[6].tile_state.state , \mchip.row_sel[4].col_sel[5].tile_state.state , \mchip.row_sel[4].col_sel[4].tile_state.state , \mchip.row_sel[4].col_sel[3].tile_state.state , \mchip.row_sel[4].col_sel[2].tile_state.state , \mchip.row_sel[4].col_sel[1].tile_state.state , \mchip.row_sel[4].col_sel[0].tile_state.state , \mchip.row_sel[3].col_sel[7].tile_state.state , \mchip.row_sel[3].col_sel[6].tile_state.state , \mchip.row_sel[3].col_sel[5].tile_state.state , \mchip.row_sel[3].col_sel[4].tile_state.state , \mchip.row_sel[3].col_sel[3].tile_state.state , \mchip.row_sel[3].col_sel[2].tile_state.state , \mchip.row_sel[3].col_sel[1].tile_state.state , \mchip.row_sel[3].col_sel[0].tile_state.state , \mchip.row_sel[2].col_sel[7].tile_state.state , \mchip.row_sel[2].col_sel[6].tile_state.state , \mchip.row_sel[2].col_sel[5].tile_state.state , \mchip.row_sel[2].col_sel[4].tile_state.state , \mchip.row_sel[2].col_sel[3].tile_state.state , \mchip.row_sel[2].col_sel[2].tile_state.state , \mchip.row_sel[2].col_sel[1].tile_state.state , \mchip.row_sel[2].col_sel[0].tile_state.state , \mchip.row_sel[1].col_sel[7].tile_state.state , \mchip.row_sel[1].col_sel[6].tile_state.state , \mchip.row_sel[1].col_sel[5].tile_state.state , \mchip.row_sel[1].col_sel[4].tile_state.state , \mchip.row_sel[1].col_sel[3].tile_state.state , \mchip.row_sel[1].col_sel[2].tile_state.state , \mchip.row_sel[1].col_sel[1].tile_state.state , \mchip.row_sel[1].col_sel[0].tile_state.state , \mchip.row_sel[0].col_sel[7].tile_state.state , \mchip.row_sel[0].col_sel[6].tile_state.state , \mchip.row_sel[0].col_sel[5].tile_state.state , \mchip.row_sel[0].col_sel[4].tile_state.state , \mchip.row_sel[0].col_sel[3].tile_state.state , \mchip.row_sel[0].col_sel[2].tile_state.state , \mchip.row_sel[0].col_sel[1].tile_state.state , \mchip.row_sel[0].col_sel[0].tile_state.state };
	assign \mchip.top  = 640'h5795e5795e5795e5795e4b12c4b12c4b12c4b12c3e8fa3e8fa3e8fa3e8fa320c8320c8320c8320c825896258962589625896190641906419064190640c8320c8320c8320c83200000000000000000000;
	assign \mchip.v_idx  = \mchip.vga.v_idx ;
	assign \mchip.vga.clk  = io_in[12];
	assign \mchip.vga.rst  = io_in[13];
	assign \mchip.vsync  = \mchip.vga.vsync ;
endmodule
module d13_thomaska_cordic (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	reg _0064_;
	reg _0065_;
	reg _0066_;
	reg _0067_;
	reg _0068_;
	reg _0069_;
	reg _0070_;
	reg _0071_;
	reg _0072_;
	reg _0073_;
	reg _0074_;
	reg _0075_;
	reg _0076_;
	reg _0077_;
	reg _0078_;
	reg _0079_;
	reg _0080_;
	reg _0081_;
	reg _0082_;
	reg _0083_;
	reg _0084_;
	reg _0085_;
	reg _0086_;
	reg _0087_;
	reg _0088_;
	reg _0089_;
	reg _0090_;
	reg _0091_;
	reg _0092_;
	reg _0093_;
	reg _0094_;
	reg _0095_;
	reg _0096_;
	reg _0097_;
	reg _0098_;
	reg _0099_;
	reg _0100_;
	reg _0101_;
	reg _0102_;
	reg _0103_;
	reg _0104_;
	reg _0105_;
	reg _0106_;
	reg _0107_;
	reg _0108_;
	reg _0109_;
	reg _0110_;
	reg _0111_;
	reg _0112_;
	reg _0113_;
	reg _0114_;
	reg _0115_;
	reg _0116_;
	reg _0117_;
	reg _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire _2025_;
	wire _2026_;
	wire _2027_;
	wire _2028_;
	wire _2029_;
	wire _2030_;
	wire _2031_;
	wire _2032_;
	wire _2033_;
	wire _2034_;
	wire _2035_;
	wire _2036_;
	wire _2037_;
	wire _2038_;
	wire _2039_;
	wire _2040_;
	wire _2041_;
	wire _2042_;
	wire _2043_;
	wire _2044_;
	wire _2045_;
	wire _2046_;
	wire _2047_;
	wire _2048_;
	wire _2049_;
	wire _2050_;
	wire _2051_;
	wire _2052_;
	wire _2053_;
	wire _2054_;
	wire _2055_;
	wire _2056_;
	wire _2057_;
	wire _2058_;
	wire _2059_;
	wire _2060_;
	wire _2061_;
	wire _2062_;
	wire _2063_;
	wire _2064_;
	wire _2065_;
	wire _2066_;
	wire _2067_;
	wire _2068_;
	wire _2069_;
	wire _2070_;
	wire _2071_;
	wire _2072_;
	wire _2073_;
	wire _2074_;
	wire _2075_;
	wire _2076_;
	wire _2077_;
	wire _2078_;
	wire _2079_;
	wire _2080_;
	wire _2081_;
	wire _2082_;
	wire _2083_;
	wire _2084_;
	wire _2085_;
	wire _2086_;
	wire _2087_;
	wire _2088_;
	wire _2089_;
	wire _2090_;
	wire _2091_;
	wire _2092_;
	wire _2093_;
	wire _2094_;
	wire _2095_;
	wire _2096_;
	wire _2097_;
	wire _2098_;
	wire _2099_;
	wire _2100_;
	wire _2101_;
	wire _2102_;
	wire _2103_;
	wire _2104_;
	wire _2105_;
	wire _2106_;
	wire _2107_;
	wire _2108_;
	wire _2109_;
	wire _2110_;
	wire _2111_;
	wire _2112_;
	wire _2113_;
	wire _2114_;
	wire _2115_;
	wire _2116_;
	wire _2117_;
	wire _2118_;
	wire _2119_;
	wire _2120_;
	wire _2121_;
	wire _2122_;
	wire _2123_;
	wire _2124_;
	wire _2125_;
	wire _2126_;
	wire _2127_;
	wire _2128_;
	wire _2129_;
	wire _2130_;
	wire _2131_;
	wire _2132_;
	wire _2133_;
	wire [2:0] _2134_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire \mchip.cordic_module.clk ;
	wire \mchip.cordic_module.done ;
	wire \mchip.cordic_module.fstage_0.clk ;
	wire \mchip.cordic_module.fstage_0.mode ;
	wire [16:0] \mchip.cordic_module.fstage_0.out_x ;
	wire \mchip.cordic_module.fstage_0.reset ;
	wire \mchip.cordic_module.fstage_0.stage_0.clk ;
	wire \mchip.cordic_module.fstage_0.stage_0.mode ;
	wire \mchip.cordic_module.fstage_0.stage_0.reset ;
	wire [4:0] \mchip.cordic_module.fstage_0.stage_0.step_ctr ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_0.subx.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_0.suby.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_0.subz.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_0.subz.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_0.subz.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_0.x_coeff ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_0.y_coeff ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_0.z_coeff ;
	wire \mchip.cordic_module.fstage_0.stage_1.clk ;
	wire \mchip.cordic_module.fstage_0.stage_1.mode ;
	wire \mchip.cordic_module.fstage_0.stage_1.reset ;
	wire [4:0] \mchip.cordic_module.fstage_0.stage_1.step_ctr ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_1.subx.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_1.subx.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_1.suby.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_1.suby.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_1.subz.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_1.subz.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_1.subz.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_1.z_coeff ;
	wire \mchip.cordic_module.fstage_0.stage_2.clk ;
	wire \mchip.cordic_module.fstage_0.stage_2.mode ;
	wire \mchip.cordic_module.fstage_0.stage_2.reset ;
	wire [4:0] \mchip.cordic_module.fstage_0.stage_2.step_ctr ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_2.subx.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_2.subx.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_2.suby.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_2.suby.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_2.subz.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_2.subz.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_2.subz.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_2.z_coeff ;
	wire \mchip.cordic_module.fstage_0.stage_3.clk ;
	wire \mchip.cordic_module.fstage_0.stage_3.mode ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.out_x ;
	wire \mchip.cordic_module.fstage_0.stage_3.reset ;
	wire [4:0] \mchip.cordic_module.fstage_0.stage_3.step_ctr ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.subx.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.subx.inside_add.out ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.subx.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.subx.out ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.suby.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.suby.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.subz.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.subz.inside_add.in_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.subz.modified_b ;
	wire [16:0] \mchip.cordic_module.fstage_0.stage_3.z_coeff ;
	wire [4:0] \mchip.cordic_module.fstage_0.step_ctr ;
	wire [16:0] \mchip.cordic_module.fstage_0.z_coeff_0 ;
	wire [16:0] \mchip.cordic_module.fstage_0.z_coeff_1 ;
	wire [16:0] \mchip.cordic_module.fstage_0.z_coeff_2 ;
	wire [16:0] \mchip.cordic_module.fstage_0.z_coeff_3 ;
	wire [9:0] \mchip.cordic_module.in_val ;
	wire [16:0] \mchip.cordic_module.in_val_32768 ;
	wire [16:0] \mchip.cordic_module.in_x_32768 ;
	wire [16:0] \mchip.cordic_module.in_y_32768 ;
	wire [16:0] \mchip.cordic_module.init_x ;
	wire [16:0] \mchip.cordic_module.init_y ;
	wire [16:0] \mchip.cordic_module.init_z ;
	wire \mchip.cordic_module.mode_toggle ;
	wire [16:0] \mchip.cordic_module.next_x ;
	wire [16:0] \mchip.cordic_module.out1 ;
	wire [16:0] \mchip.cordic_module.out2 ;
	wire \mchip.cordic_module.out_toggle ;
	wire \mchip.cordic_module.rst ;
	wire [4:0] \mchip.cordic_module.step_ctr_4 ;
	wire [10:0] \mchip.cordic_module.val ;
	wire [16:0] \mchip.cordic_module.z_coeff[0] ;
	wire [16:0] \mchip.cordic_module.z_coeff[10] ;
	wire [16:0] \mchip.cordic_module.z_coeff[11] ;
	wire [16:0] \mchip.cordic_module.z_coeff[12] ;
	wire [16:0] \mchip.cordic_module.z_coeff[13] ;
	wire [16:0] \mchip.cordic_module.z_coeff[14] ;
	wire [16:0] \mchip.cordic_module.z_coeff[15] ;
	wire [16:0] \mchip.cordic_module.z_coeff[1] ;
	wire [16:0] \mchip.cordic_module.z_coeff[2] ;
	wire [16:0] \mchip.cordic_module.z_coeff[3] ;
	wire [16:0] \mchip.cordic_module.z_coeff[4] ;
	wire [16:0] \mchip.cordic_module.z_coeff[5] ;
	wire [16:0] \mchip.cordic_module.z_coeff[6] ;
	wire [16:0] \mchip.cordic_module.z_coeff[7] ;
	wire [16:0] \mchip.cordic_module.z_coeff[8] ;
	wire [16:0] \mchip.cordic_module.z_coeff[9] ;
	wire [16:0] \mchip.cordic_module.z_coeff_group[0] ;
	wire [16:0] \mchip.cordic_module.z_coeff_group[1] ;
	wire [16:0] \mchip.cordic_module.z_coeff_group[2] ;
	wire [16:0] \mchip.cordic_module.z_coeff_group[3] ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign \mchip.cordic_module.fstage_0.stage_0.step_ctr [2] = io_in[13] | ~_0099_;
	assign _0936_ = _0100_ & ~io_in[13];
	assign _0946_ = \mchip.cordic_module.fstage_0.stage_0.step_ctr [2] & ~_0936_;
	assign _0957_ = _0101_ & ~io_in[13];
	assign _0001_ = ~(_0957_ & _0946_);
	assign _0000_ = ~(_0001_ | io_in[13]);
	assign io_out[0] = (io_in[11] ? \mchip.cordic_module.out1 [6] : \mchip.cordic_module.out2 [6]);
	assign io_out[1] = (io_in[11] ? \mchip.cordic_module.out1 [7] : \mchip.cordic_module.out2 [7]);
	assign io_out[2] = (io_in[11] ? \mchip.cordic_module.out1 [8] : \mchip.cordic_module.out2 [8]);
	assign io_out[3] = (io_in[11] ? \mchip.cordic_module.out1 [9] : \mchip.cordic_module.out2 [9]);
	assign io_out[4] = (io_in[11] ? \mchip.cordic_module.out1 [10] : \mchip.cordic_module.out2 [10]);
	assign io_out[5] = (io_in[11] ? \mchip.cordic_module.out1 [11] : \mchip.cordic_module.out2 [11]);
	assign io_out[6] = (io_in[11] ? \mchip.cordic_module.out1 [12] : \mchip.cordic_module.out2 [12]);
	assign io_out[7] = (io_in[11] ? \mchip.cordic_module.out1 [13] : \mchip.cordic_module.out2 [13]);
	assign io_out[8] = (io_in[11] ? \mchip.cordic_module.out1 [14] : \mchip.cordic_module.out2 [14]);
	assign io_out[9] = (io_in[11] ? \mchip.cordic_module.out1 [15] : \mchip.cordic_module.out2 [15]);
	assign io_out[10] = (io_in[11] ? \mchip.cordic_module.out1 [16] : \mchip.cordic_module.out2 [16]);
	assign _1091_ = ~io_in[10];
	assign _1102_ = _0957_ ^ _0946_;
	assign _1113_ = io_in[13] | ~_0096_;
	assign _1123_ = io_in[13] | ~_0097_;
	assign _1131_ = _0080_ & ~io_in[13];
	assign _1137_ = (io_in[10] ? _1123_ : _1131_);
	assign _1143_ = io_in[13] | ~_0118_;
	assign _1150_ = _0936_ ^ \mchip.cordic_module.fstage_0.stage_0.step_ctr [2];
	assign _1158_ = io_in[13] | ~_0117_;
	assign _1163_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1143_ : _1158_);
	assign _1169_ = (_1150_ ? _1143_ : _1163_);
	assign _1177_ = (_1102_ ? _1143_ : _1169_);
	assign _1187_ = ~(_1177_ ^ _1137_);
	assign _1197_ = _1187_ ^ _1113_;
	assign _1208_ = io_in[13] | ~_0095_;
	assign _1218_ = io_in[13] | ~_0116_;
	assign _1228_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1143_ : _1218_);
	assign _1238_ = (_1150_ ? _1143_ : _1228_);
	assign _1248_ = (_1102_ ? _1143_ : _1238_);
	assign _1257_ = ~(_1248_ ^ _1137_);
	assign _1266_ = _1208_ | ~_1257_;
	assign _1277_ = ~(_1257_ ^ _1208_);
	assign _1286_ = io_in[13] | ~_0094_;
	assign _1295_ = io_in[13] | ~_0115_;
	assign _1304_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1143_ : _1295_);
	assign _1313_ = (_1150_ ? _1143_ : _1304_);
	assign _1324_ = (_1102_ ? _1143_ : _1313_);
	assign _1332_ = ~(_1324_ ^ _1137_);
	assign _1341_ = _1286_ | ~_1332_;
	assign _1349_ = io_in[13] | ~_0093_;
	assign _1360_ = io_in[13] | ~_0114_;
	assign _1363_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1143_ : _1360_);
	assign _1364_ = (_1150_ ? _1143_ : _1363_);
	assign _1365_ = (_1102_ ? _1143_ : _1364_);
	assign _1366_ = ~(_1365_ ^ _1137_);
	assign _1367_ = _1366_ & ~_1349_;
	assign _1368_ = ~(_1332_ ^ _1286_);
	assign _1369_ = _1368_ & _1367_;
	assign _1370_ = _1341_ & ~_1369_;
	assign _1371_ = _1366_ ^ _1349_;
	assign _1372_ = _1368_ & ~_1371_;
	assign _1373_ = io_in[13] | ~_0092_;
	assign _1374_ = ~_1373_;
	assign _1375_ = io_in[13] | ~_0113_;
	assign _1376_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1158_ : _1375_);
	assign _1377_ = (_1150_ ? _1143_ : _1376_);
	assign _1378_ = (_1102_ ? _1143_ : _1377_);
	assign _1379_ = ~(_1378_ ^ _1137_);
	assign _1380_ = ~(_1379_ & _1374_);
	assign _1381_ = _1379_ ^ _1374_;
	assign _1382_ = io_in[13] | ~_0091_;
	assign _1383_ = io_in[13] | ~_0112_;
	assign _1384_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1218_ : _1383_);
	assign _1385_ = (_1150_ ? _1143_ : _1384_);
	assign _1386_ = (_1102_ ? _1143_ : _1385_);
	assign _1387_ = ~(_1386_ ^ _1137_);
	assign _1388_ = _1382_ | ~_1387_;
	assign _1389_ = _1381_ & ~_1388_;
	assign _1390_ = _1380_ & ~_1389_;
	assign _1391_ = _1387_ ^ _1382_;
	assign _1392_ = _1381_ & ~_1391_;
	assign _1393_ = io_in[13] | ~_0090_;
	assign _1394_ = io_in[13] | ~_0111_;
	assign _1395_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1295_ : _1394_);
	assign _1396_ = (_1150_ ? _1143_ : _1395_);
	assign _1397_ = (_1102_ ? _1143_ : _1396_);
	assign _1398_ = ~(_1397_ ^ _1137_);
	assign _1399_ = _1398_ & ~_1393_;
	assign _1400_ = _1398_ ^ _1393_;
	assign _1401_ = io_in[13] | ~_0089_;
	assign _1402_ = ~_1143_;
	assign _1403_ = _0114_ & ~io_in[13];
	assign _1404_ = _0110_ & ~io_in[13];
	assign _1405_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1403_ : _1404_);
	assign _1406_ = (_1150_ ? _1402_ : _1405_);
	assign _1407_ = (_1102_ ? _1402_ : _1406_);
	assign _1408_ = _1407_ ^ _1137_;
	assign _1409_ = _1401_ | ~_1408_;
	assign _1410_ = _1409_ | _1400_;
	assign _1411_ = _1410_ & ~_1399_;
	assign _1412_ = _1392_ & ~_1411_;
	assign _1413_ = _1390_ & ~_1412_;
	assign _1414_ = _1408_ ^ _1401_;
	assign _1415_ = _1414_ | _1400_;
	assign _1416_ = _1392_ & ~_1415_;
	assign _1417_ = io_in[13] | ~_0088_;
	assign _1418_ = ~_1417_;
	assign _1419_ = io_in[13] | ~_0109_;
	assign _1420_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1375_ : _1419_);
	assign _1421_ = (_1150_ ? _1163_ : _1420_);
	assign _1422_ = (_1102_ ? _1143_ : _1421_);
	assign _1423_ = ~(_1422_ ^ _1137_);
	assign _1424_ = ~(_1423_ & _1418_);
	assign _1425_ = _1423_ ^ _1418_;
	assign _1426_ = io_in[13] | ~_0087_;
	assign _1427_ = io_in[13] | ~_0108_;
	assign _1428_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1383_ : _1427_);
	assign _1429_ = (_1150_ ? _1228_ : _1428_);
	assign _1430_ = (_1102_ ? _1143_ : _1429_);
	assign _1431_ = ~(_1430_ ^ _1137_);
	assign _1432_ = _1426_ | ~_1431_;
	assign _1433_ = _1425_ & ~_1432_;
	assign _1434_ = _1424_ & ~_1433_;
	assign _1435_ = _1431_ ^ _1426_;
	assign _1436_ = _1425_ & ~_1435_;
	assign _1437_ = io_in[13] | ~_0086_;
	assign _1438_ = ~_1437_;
	assign _1439_ = io_in[13] | ~_0107_;
	assign _1440_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1394_ : _1439_);
	assign _1441_ = (_1150_ ? _1304_ : _1440_);
	assign _1442_ = (_1102_ ? _1143_ : _1441_);
	assign _1443_ = ~(_1442_ ^ _1137_);
	assign _1444_ = ~(_1443_ & _1438_);
	assign _1445_ = _1443_ ^ _1438_;
	assign _1446_ = io_in[13] | ~_0085_;
	assign _1447_ = io_in[13] | ~_0110_;
	assign _1448_ = io_in[13] | ~_0106_;
	assign _1449_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1447_ : _1448_);
	assign _1450_ = (_1150_ ? _1363_ : _1449_);
	assign _1451_ = (_1102_ ? _1143_ : _1450_);
	assign _1452_ = ~(_1451_ ^ _1137_);
	assign _1453_ = _1446_ | ~_1452_;
	assign _1454_ = _1445_ & ~_1453_;
	assign _1455_ = _1444_ & ~_1454_;
	assign _1456_ = _1436_ & ~_1455_;
	assign _1457_ = _1434_ & ~_1456_;
	assign _1458_ = _1452_ ^ _1446_;
	assign _1459_ = _1458_ | ~_1445_;
	assign _1460_ = _1436_ & ~_1459_;
	assign _1461_ = io_in[13] | ~_0084_;
	assign _1462_ = ~_1461_;
	assign _1463_ = io_in[13] | ~_0105_;
	assign _1464_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1419_ : _1463_);
	assign _1465_ = (_1150_ ? _1376_ : _1464_);
	assign _1466_ = (_1102_ ? _1143_ : _1465_);
	assign _1467_ = ~(_1466_ ^ _1137_);
	assign _1468_ = ~(_1467_ & _1462_);
	assign _1469_ = _1467_ ^ _1462_;
	assign _1470_ = io_in[13] | ~_0083_;
	assign _1471_ = io_in[13] | ~_0104_;
	assign _1472_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1427_ : _1471_);
	assign _1473_ = (_1150_ ? _1384_ : _1472_);
	assign _1474_ = (_1102_ ? _1143_ : _1473_);
	assign _1475_ = ~(_1474_ ^ _1137_);
	assign _1476_ = _1470_ | ~_1475_;
	assign _1477_ = _1469_ & ~_1476_;
	assign _1478_ = _1468_ & ~_1477_;
	assign _1479_ = _1475_ ^ _1470_;
	assign _1480_ = _1469_ & ~_1479_;
	assign _1481_ = io_in[13] | ~_0082_;
	assign _1482_ = ~_1481_;
	assign _1483_ = io_in[13] | ~_0103_;
	assign _1484_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1439_ : _1483_);
	assign _1485_ = (_1150_ ? _1395_ : _1484_);
	assign _1486_ = (_1102_ ? _1143_ : _1485_);
	assign _1487_ = ~(_1486_ ^ _1137_);
	assign _1488_ = ~(_1487_ & _1482_);
	assign _1489_ = _1487_ ^ _1482_;
	assign _1490_ = io_in[13] | ~_0081_;
	assign _1491_ = ~_1137_;
	assign _1492_ = _0106_ & ~io_in[13];
	assign _1493_ = _0102_ & ~io_in[13];
	assign _1494_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1492_ : _1493_);
	assign _1495_ = (_1150_ ? _1405_ : _1494_);
	assign _1496_ = (_1102_ ? _1402_ : _1495_);
	assign _1497_ = (_1496_ ? _1490_ : _1491_);
	assign _1498_ = _1489_ & ~_1497_;
	assign _1499_ = _1488_ & ~_1498_;
	assign _1500_ = _1480_ & ~_1499_;
	assign _1501_ = _1478_ & ~_1500_;
	assign _1502_ = _1460_ & ~_1501_;
	assign _1503_ = _1457_ & ~_1502_;
	assign _1504_ = _1416_ & ~_1503_;
	assign _1505_ = _1413_ & ~_1504_;
	assign _1506_ = _1372_ & ~_1505_;
	assign _1507_ = _1370_ & ~_1506_;
	assign _1508_ = _1277_ & ~_1507_;
	assign _1509_ = _1266_ & ~_1508_;
	assign _1510_ = _1509_ ^ _1197_;
	assign _1511_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1123_ : _1113_);
	assign _1512_ = (_1150_ ? _1123_ : _1511_);
	assign _1513_ = (_1102_ ? _1123_ : _1512_);
	assign _1514_ = ~_1123_;
	assign _1515_ = ~_1131_;
	assign _1516_ = (io_in[10] ? _1514_ : _1515_);
	assign _1517_ = ~_1516_;
	assign _1518_ = _1517_ ^ _1513_;
	assign _1519_ = _1518_ & ~_1158_;
	assign _1520_ = _1158_ ^ _1518_;
	assign _1521_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1123_ : _1208_);
	assign _1522_ = (_1150_ ? _1123_ : _1521_);
	assign _1523_ = (_1102_ ? _1123_ : _1522_);
	assign _1524_ = _1523_ ^ _1516_;
	assign _1525_ = _1218_ | _1524_;
	assign _1526_ = ~(_1525_ | _1520_);
	assign _1527_ = ~(_1526_ | _1519_);
	assign _1528_ = _1218_ ^ _1524_;
	assign _1529_ = _1528_ & ~_1520_;
	assign _1530_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1123_ : _1286_);
	assign _1531_ = (_1150_ ? _1123_ : _1530_);
	assign _1532_ = (_1102_ ? _1123_ : _1531_);
	assign _1533_ = _1532_ ^ _1516_;
	assign _1534_ = _1295_ | _1533_;
	assign _1535_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1123_ : _1349_);
	assign _1536_ = (_1150_ ? _1123_ : _1535_);
	assign _1537_ = (_1102_ ? _1123_ : _1536_);
	assign _1538_ = _1537_ ^ _1517_;
	assign _1539_ = _1538_ & ~_1360_;
	assign _1540_ = _1295_ ^ _1533_;
	assign _1541_ = _1540_ & _1539_;
	assign _1542_ = _1534_ & ~_1541_;
	assign _1543_ = _1529_ & ~_1542_;
	assign _1544_ = _1527_ & ~_1543_;
	assign _1545_ = _1360_ ^ _1538_;
	assign _1546_ = _1540_ & ~_1545_;
	assign _1547_ = _1546_ & _1529_;
	assign _1548_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1113_ : _1373_);
	assign _1549_ = (_1150_ ? _1123_ : _1548_);
	assign _1550_ = (_1102_ ? _1123_ : _1549_);
	assign _1551_ = _1550_ ^ _1517_;
	assign _1552_ = ~_1375_;
	assign _1553_ = ~(_1552_ & _1551_);
	assign _1554_ = _1552_ ^ _1551_;
	assign _1555_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1208_ : _1382_);
	assign _1556_ = (_1150_ ? _1123_ : _1555_);
	assign _1557_ = (_1102_ ? _1123_ : _1556_);
	assign _1558_ = _1557_ ^ _1516_;
	assign _1559_ = _1383_ | _1558_;
	assign _1560_ = _1554_ & ~_1559_;
	assign _1561_ = _1553_ & ~_1560_;
	assign _1562_ = ~(_1383_ ^ _1558_);
	assign _1563_ = _1554_ & ~_1562_;
	assign _1564_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1286_ : _1393_);
	assign _1565_ = (_1150_ ? _1123_ : _1564_);
	assign _1566_ = (_1102_ ? _1123_ : _1565_);
	assign _1567_ = _1566_ ^ _1516_;
	assign _1568_ = _1394_ | _1567_;
	assign _1569_ = ~(_1394_ ^ _1567_);
	assign _1570_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1349_ : _1401_);
	assign _1571_ = (_1150_ ? _1123_ : _1570_);
	assign _1572_ = (_1102_ ? _1123_ : _1571_);
	assign _1573_ = _1572_ ^ _1516_;
	assign _1574_ = _1447_ | _1573_;
	assign _1575_ = ~(_1574_ | _1569_);
	assign _1576_ = _1568_ & ~_1575_;
	assign _1577_ = _1563_ & ~_1576_;
	assign _1578_ = _1561_ & ~_1577_;
	assign _1579_ = _1547_ & ~_1578_;
	assign _1580_ = _1544_ & ~_1579_;
	assign _1581_ = _1404_ ^ _1573_;
	assign _1582_ = _1581_ | _1569_;
	assign _1583_ = _1563_ & ~_1582_;
	assign _1584_ = _1583_ & _1547_;
	assign _1585_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1373_ : _1417_);
	assign _1586_ = (_1150_ ? _1511_ : _1585_);
	assign _1587_ = (_1102_ ? _1123_ : _1586_);
	assign _1588_ = _1587_ ^ _1516_;
	assign _1589_ = _1419_ | _1588_;
	assign _1590_ = _1419_ ^ _1588_;
	assign _1591_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1382_ : _1426_);
	assign _1592_ = (_1150_ ? _1521_ : _1591_);
	assign _1593_ = (_1102_ ? _1123_ : _1592_);
	assign _1594_ = _1593_ ^ _1516_;
	assign _1595_ = _1427_ | _1594_;
	assign _1596_ = _1590_ & ~_1595_;
	assign _1597_ = _1589_ & ~_1596_;
	assign _1598_ = ~(_1427_ ^ _1594_);
	assign _1599_ = _1590_ & ~_1598_;
	assign _1600_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1393_ : _1437_);
	assign _1601_ = (_1150_ ? _1530_ : _1600_);
	assign _1602_ = (_1102_ ? _1123_ : _1601_);
	assign _1603_ = _1602_ ^ _1516_;
	assign _1604_ = _1439_ | _1603_;
	assign _1605_ = _1439_ ^ _1603_;
	assign _1606_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1401_ : _1446_);
	assign _1607_ = (_1150_ ? _1535_ : _1606_);
	assign _1608_ = (_1102_ ? _1123_ : _1607_);
	assign _1609_ = _1608_ ^ _1516_;
	assign _1610_ = _1448_ | _1609_;
	assign _1611_ = _1605_ & ~_1610_;
	assign _1612_ = _1604_ & ~_1611_;
	assign _1613_ = _1599_ & ~_1612_;
	assign _1614_ = _1597_ & ~_1613_;
	assign _1615_ = _1492_ ^ _1609_;
	assign _1616_ = _1615_ | ~_1605_;
	assign _1617_ = _1599_ & ~_1616_;
	assign _1618_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1417_ : _1461_);
	assign _1619_ = (_1150_ ? _1548_ : _1618_);
	assign _1620_ = (_1102_ ? _1123_ : _1619_);
	assign _1621_ = _1620_ ^ _1516_;
	assign _1622_ = _1463_ | _1621_;
	assign _1623_ = _1463_ ^ _1621_;
	assign _1624_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1426_ : _1470_);
	assign _1625_ = (_1150_ ? _1555_ : _1624_);
	assign _1626_ = (_1102_ ? _1123_ : _1625_);
	assign _1627_ = _1626_ ^ _1516_;
	assign _1628_ = _1471_ | _1627_;
	assign _1629_ = _1623_ & ~_1628_;
	assign _1630_ = _1622_ & ~_1629_;
	assign _1631_ = ~_1471_;
	assign _1632_ = _1631_ ^ _1627_;
	assign _1633_ = _1623_ & ~_1632_;
	assign _1634_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1437_ : _1481_);
	assign _1635_ = (_1150_ ? _1564_ : _1634_);
	assign _1636_ = (_1102_ ? _1123_ : _1635_);
	assign _1637_ = _1636_ ^ _1516_;
	assign _1638_ = _1483_ | _1637_;
	assign _1639_ = _1483_ ^ _1637_;
	assign _1640_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1446_ : _1490_);
	assign _1641_ = (_1150_ ? _1570_ : _1640_);
	assign _1642_ = (_1102_ ? _1123_ : _1641_);
	assign _1643_ = ~_1493_;
	assign _1644_ = (_1642_ ? _1517_ : _1643_);
	assign _1645_ = _1639_ & ~_1644_;
	assign _1646_ = _1638_ & ~_1645_;
	assign _1647_ = _1633_ & ~_1646_;
	assign _1648_ = _1630_ & ~_1647_;
	assign _1649_ = _1617_ & ~_1648_;
	assign _1650_ = _1614_ & ~_1649_;
	assign _1651_ = _1584_ & ~_1650_;
	assign _1652_ = _1580_ & ~_1651_;
	assign _1653_ = ~(_1137_ ^ _1123_);
	assign _1654_ = _1402_ ^ _1653_;
	assign _1655_ = _1654_ ^ _1652_;
	assign _1656_ = _0079_ & ~io_in[13];
	assign _1657_ = _1656_ & ~_1137_;
	assign _1658_ = _1656_ ^ _1137_;
	assign _1659_ = _0936_ | \mchip.cordic_module.fstage_0.stage_0.step_ctr [2];
	assign _1660_ = _1659_ | _0957_;
	assign _1661_ = _1660_ ^ _1137_;
	assign _1662_ = _0078_ & ~io_in[13];
	assign _1663_ = ~(_1662_ & _1661_);
	assign _1664_ = ~(_1663_ | _1658_);
	assign _1665_ = ~(_1664_ | _1657_);
	assign _1666_ = _1662_ ^ _1661_;
	assign _1667_ = _1666_ & ~_1658_;
	assign _1668_ = _0077_ & ~io_in[13];
	assign _1669_ = ~(_1668_ & _1661_);
	assign _1670_ = _0076_ & ~io_in[13];
	assign _1671_ = _1670_ & _1516_;
	assign _1672_ = ~_1671_;
	assign _1673_ = _1668_ ^ _1661_;
	assign _1674_ = _1673_ & ~_1672_;
	assign _1675_ = _1669_ & ~_1674_;
	assign _1676_ = _1667_ & ~_1675_;
	assign _1677_ = _1665_ & ~_1676_;
	assign _1678_ = _1670_ ^ _1137_;
	assign _1679_ = _1673_ & ~_1678_;
	assign _1680_ = _1679_ & _1667_;
	assign _1681_ = _0075_ & ~io_in[13];
	assign _1682_ = ~(_1681_ & _1516_);
	assign _1683_ = ~(_1681_ ^ _1137_);
	assign _1684_ = ~(_0936_ & \mchip.cordic_module.fstage_0.stage_0.step_ctr [2]);
	assign _1685_ = ~(_1684_ | _0957_);
	assign _1686_ = _0936_ & ~\mchip.cordic_module.fstage_0.stage_0.step_ctr [2];
	assign _1687_ = (_0957_ ? _0946_ : _1686_);
	assign _1688_ = _1685_ | ~_1660_;
	assign _1689_ = _1688_ ^ _1517_;
	assign _1690_ = _0074_ & ~io_in[13];
	assign _1691_ = _1689_ | ~_1690_;
	assign _1692_ = _1683_ & ~_1691_;
	assign _1693_ = _1682_ & ~_1692_;
	assign _1694_ = _1690_ ^ _1689_;
	assign _1695_ = _1683_ & ~_1694_;
	assign _1696_ = _1660_ & ~_1685_;
	assign _1697_ = _1687_ | ~_1696_;
	assign _1698_ = _1697_ & _1685_;
	assign _1699_ = _1698_ ^ _1516_;
	assign _1700_ = _0073_ & ~io_in[13];
	assign _1701_ = ~(_1700_ & _1699_);
	assign _1702_ = _1700_ ^ _1699_;
	assign _1703_ = _0072_ & ~io_in[13];
	assign _1704_ = ~(_1703_ & _1699_);
	assign _1705_ = _1702_ & ~_1704_;
	assign _1706_ = _1701_ & ~_1705_;
	assign _1707_ = _1695_ & ~_1706_;
	assign _1708_ = _1693_ & ~_1707_;
	assign _1709_ = _1680_ & ~_1708_;
	assign _1710_ = _1677_ & ~_1709_;
	assign _1711_ = ~(_1703_ ^ _1699_);
	assign _1712_ = _1711_ | ~_1702_;
	assign _1713_ = _1695_ & ~_1712_;
	assign _1714_ = _1713_ & _1680_;
	assign _1715_ = _1686_ & ~_0957_;
	assign _1716_ = _1696_ & ~_1715_;
	assign _1717_ = _1697_ & ~_1716_;
	assign _1718_ = _1717_ ^ _1516_;
	assign _1719_ = _0071_ & ~io_in[13];
	assign _1720_ = ~(_1719_ & _1718_);
	assign _1721_ = ~(_1719_ ^ _1718_);
	assign _1722_ = _0070_ & ~io_in[13];
	assign _1723_ = ~(_1722_ & _1699_);
	assign _1724_ = ~(_1723_ | _1721_);
	assign _1725_ = _1720_ & ~_1724_;
	assign _1726_ = _1722_ ^ _1699_;
	assign _1727_ = _1726_ & ~_1721_;
	assign _1728_ = _0069_ & ~io_in[13];
	assign _1729_ = ~(_1728_ & _1699_);
	assign _1730_ = _1728_ ^ _1699_;
	assign _1731_ = _0068_ & ~io_in[13];
	assign _1732_ = ~(_1731_ & _1699_);
	assign _1733_ = _1730_ & ~_1732_;
	assign _1734_ = _1729_ & ~_1733_;
	assign _1735_ = _1727_ & ~_1734_;
	assign _1736_ = _1725_ & ~_1735_;
	assign _1737_ = ~(_1731_ ^ _1699_);
	assign _1738_ = _1730_ & ~_1737_;
	assign _1739_ = _1738_ & _1727_;
	assign _1740_ = _1696_ & _0001_;
	assign _1741_ = _1697_ & ~_1740_;
	assign _1742_ = _1741_ ^ _1516_;
	assign _1743_ = _0067_ & ~io_in[13];
	assign _1744_ = ~(_1743_ & _1742_);
	assign _1745_ = _1743_ ^ _1742_;
	assign _1746_ = _0066_ & ~io_in[13];
	assign _1747_ = ~(_1746_ & _1699_);
	assign _1748_ = _1745_ & ~_1747_;
	assign _1749_ = _1744_ & ~_1748_;
	assign _1750_ = ~(_1746_ ^ _1699_);
	assign _1751_ = _1745_ & ~_1750_;
	assign _1752_ = _0065_ & ~io_in[13];
	assign _1753_ = _1137_ | ~_1752_;
	assign _1754_ = _1752_ ^ _1137_;
	assign _1755_ = _0064_ & ~io_in[13];
	assign _1756_ = ~_1755_;
	assign _1757_ = (_1698_ ? _1756_ : _1517_);
	assign _1758_ = ~(_1757_ | _1754_);
	assign _1759_ = _1753_ & ~_1758_;
	assign _1760_ = _1751_ & ~_1759_;
	assign _1761_ = _1749_ & ~_1760_;
	assign _1762_ = _1739_ & ~_1761_;
	assign _1763_ = _1736_ & ~_1762_;
	assign _1764_ = _1714_ & ~_1763_;
	assign _1765_ = _1710_ & ~_1764_;
	assign _1766_ = _1137_ ^ _1515_;
	assign _1767_ = _1766_ ^ _1765_;
	assign _1768_ = _1187_ & ~_1113_;
	assign _1769_ = ~(_1266_ | _1197_);
	assign _1770_ = ~(_1769_ | _1768_);
	assign _1771_ = _1277_ & ~_1197_;
	assign _1772_ = _1771_ & ~_1370_;
	assign _1773_ = _1770_ & ~_1772_;
	assign _1774_ = _1372_ & _1771_;
	assign _1775_ = _1774_ & ~_1413_;
	assign _1776_ = _1773_ & ~_1775_;
	assign _1777_ = _1416_ & _1774_;
	assign _1778_ = _1777_ & ~_1503_;
	assign _1779_ = _1778_ | ~_1776_;
	assign _1780_ = ~(_1143_ ^ _1137_);
	assign _1781_ = _1780_ ^ _1514_;
	assign _1782_ = _1781_ ^ _1779_;
	assign _1783_ = (io_in[10] ? _1782_ : _1767_);
	assign _1784_ = ~(_1783_ ^ _1655_);
	assign _1785_ = ~_1784_;
	assign _1786_ = _1510_ & ~_1785_;
	assign _1787_ = _1583_ & ~_1650_;
	assign _1788_ = _1578_ & ~_1787_;
	assign _1789_ = _1546_ & ~_1788_;
	assign _1790_ = _1542_ & ~_1789_;
	assign _1791_ = _1528_ & ~_1790_;
	assign _1792_ = _1525_ & ~_1791_;
	assign _1793_ = _1792_ ^ _1520_;
	assign _1794_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1655_ : _1793_);
	assign _1795_ = (_1150_ ? _1655_ : _1794_);
	assign _1796_ = (_1102_ ? _1655_ : _1795_);
	assign _1797_ = ~(_1783_ ^ _1796_);
	assign _1798_ = ~(_1507_ ^ _1277_);
	assign _1799_ = _1798_ & _1797_;
	assign _1800_ = _1785_ ^ _1510_;
	assign _1801_ = _1799_ & ~_1800_;
	assign _1802_ = ~(_1801_ | _1786_);
	assign _1803_ = ~(_1790_ ^ _1528_);
	assign _1804_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1655_ : _1803_);
	assign _1805_ = (_1150_ ? _1655_ : _1804_);
	assign _1806_ = (_1102_ ? _1655_ : _1805_);
	assign _1807_ = ~(_1806_ ^ _1783_);
	assign _1808_ = _1505_ | _1371_;
	assign _1809_ = _1808_ & ~_1367_;
	assign _1810_ = ~(_1809_ ^ _1368_);
	assign _1811_ = ~_1810_;
	assign _1812_ = _1807_ & ~_1811_;
	assign _1813_ = _1788_ | _1545_;
	assign _1814_ = _1813_ & ~_1539_;
	assign _1815_ = ~(_1814_ ^ _1540_);
	assign _1816_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1655_ : _1815_);
	assign _1817_ = (_1150_ ? _1655_ : _1816_);
	assign _1818_ = (_1102_ ? _1655_ : _1817_);
	assign _1819_ = ~(_1818_ ^ _1783_);
	assign _1820_ = _1505_ ^ _1371_;
	assign _1821_ = _1820_ & _1819_;
	assign _1822_ = _1811_ ^ _1807_;
	assign _1823_ = _1821_ & ~_1822_;
	assign _1824_ = ~(_1823_ | _1812_);
	assign _1825_ = _1798_ ^ _1797_;
	assign _1826_ = _1800_ | ~_1825_;
	assign _1827_ = ~(_1826_ | _1824_);
	assign _1828_ = _1802_ & ~_1827_;
	assign _1829_ = _1788_ ^ _1545_;
	assign _1830_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1655_ : _1829_);
	assign _1831_ = (_1150_ ? _1655_ : _1830_);
	assign _1832_ = (_1102_ ? _1655_ : _1831_);
	assign _1833_ = ~(_1832_ ^ _1783_);
	assign _1834_ = ~(_1503_ | _1415_);
	assign _1835_ = _1411_ & ~_1834_;
	assign _1836_ = ~(_1835_ | _1391_);
	assign _1837_ = _1836_ | ~_1388_;
	assign _1838_ = _1837_ ^ _1381_;
	assign _1839_ = _1838_ & _1833_;
	assign _1840_ = _1838_ ^ _1833_;
	assign _1841_ = ~(_1650_ | _1582_);
	assign _1842_ = _1576_ & ~_1841_;
	assign _1843_ = ~(_1842_ | _1562_);
	assign _1844_ = _1843_ | ~_1559_;
	assign _1845_ = _1844_ ^ _1554_;
	assign _1846_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1793_ : _1845_);
	assign _1847_ = (_1150_ ? _1655_ : _1846_);
	assign _1848_ = (_1102_ ? _1655_ : _1847_);
	assign _1849_ = _1848_ ^ _1783_;
	assign _1850_ = _1835_ ^ _1391_;
	assign _1851_ = _1849_ | ~_1850_;
	assign _1852_ = _1840_ & ~_1851_;
	assign _1853_ = ~(_1852_ | _1839_);
	assign _1854_ = _1850_ ^ _1849_;
	assign _1855_ = _1840_ & ~_1854_;
	assign _1856_ = _1842_ ^ _1562_;
	assign _1857_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1803_ : _1856_);
	assign _1858_ = (_1150_ ? _1655_ : _1857_);
	assign _1859_ = (_1102_ ? _1655_ : _1858_);
	assign _1860_ = _1859_ ^ _1783_;
	assign _1861_ = ~(_1503_ | _1414_);
	assign _1862_ = _1409_ & ~_1861_;
	assign _1863_ = _1862_ ^ _1400_;
	assign _1864_ = _1860_ | ~_1863_;
	assign _1865_ = ~(_1863_ ^ _1860_);
	assign _1866_ = ~(_1650_ | _1581_);
	assign _1867_ = _1574_ & ~_1866_;
	assign _1868_ = _1867_ ^ _1569_;
	assign _1869_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1815_ : _1868_);
	assign _1870_ = (_1150_ ? _1655_ : _1869_);
	assign _1871_ = (_1102_ ? _1655_ : _1870_);
	assign _1872_ = _1871_ ^ _1783_;
	assign _1873_ = _1503_ ^ _1414_;
	assign _1874_ = _1872_ | ~_1873_;
	assign _1875_ = _1865_ & ~_1874_;
	assign _1876_ = _1864_ & ~_1875_;
	assign _1877_ = _1855_ & ~_1876_;
	assign _1878_ = _1853_ & ~_1877_;
	assign _1879_ = ~(_1820_ ^ _1819_);
	assign _1880_ = ~(_1879_ | _1822_);
	assign _1881_ = _1826_ | ~_1880_;
	assign _1882_ = ~(_1881_ | _1878_);
	assign _1883_ = _1828_ & ~_1882_;
	assign _1884_ = _1650_ ^ _1581_;
	assign _1885_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1829_ : _1884_);
	assign _1886_ = (_1150_ ? _1655_ : _1885_);
	assign _1887_ = (_1102_ ? _1655_ : _1886_);
	assign _1888_ = ~(_1887_ ^ _1783_);
	assign _1889_ = ~(_1501_ | _1459_);
	assign _1890_ = _1455_ & ~_1889_;
	assign _1891_ = ~(_1890_ | _1435_);
	assign _1892_ = _1891_ | ~_1432_;
	assign _1893_ = _1892_ ^ _1425_;
	assign _1894_ = ~(_1893_ & _1888_);
	assign _1895_ = ~(_1893_ ^ _1888_);
	assign _1896_ = ~_1895_;
	assign _1897_ = ~(_1648_ | _1616_);
	assign _1898_ = _1612_ & ~_1897_;
	assign _1899_ = ~(_1898_ | _1598_);
	assign _1900_ = _1899_ | ~_1595_;
	assign _1901_ = _1900_ ^ _1590_;
	assign _1902_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1845_ : _1901_);
	assign _1903_ = (_1150_ ? _1794_ : _1902_);
	assign _1904_ = (_1102_ ? _1655_ : _1903_);
	assign _1905_ = _1904_ ^ _1783_;
	assign _1906_ = _1890_ ^ _1435_;
	assign _1907_ = _1905_ | ~_1906_;
	assign _1908_ = _1896_ & ~_1907_;
	assign _1909_ = _1894_ & ~_1908_;
	assign _1910_ = _1906_ ^ _1905_;
	assign _1911_ = _1896_ & ~_1910_;
	assign _1912_ = _1898_ ^ _1598_;
	assign _1913_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1856_ : _1912_);
	assign _1914_ = (_1150_ ? _1804_ : _1913_);
	assign _1915_ = (_1102_ ? _1655_ : _1914_);
	assign _1916_ = _1915_ ^ _1783_;
	assign _1917_ = ~(_1501_ | _1458_);
	assign _1918_ = _1917_ | ~_1453_;
	assign _1919_ = _1918_ ^ _1445_;
	assign _1920_ = _1916_ | ~_1919_;
	assign _1921_ = ~(_1919_ ^ _1916_);
	assign _1922_ = ~(_1648_ | _1615_);
	assign _1923_ = _1922_ | ~_1610_;
	assign _1924_ = _1923_ ^ _1605_;
	assign _1925_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1868_ : _1924_);
	assign _1926_ = (_1150_ ? _1816_ : _1925_);
	assign _1927_ = (_1102_ ? _1655_ : _1926_);
	assign _1928_ = _1927_ ^ _1783_;
	assign _1929_ = _1501_ ^ _1458_;
	assign _1930_ = _1928_ | ~_1929_;
	assign _1931_ = _1921_ & ~_1930_;
	assign _1932_ = _1920_ & ~_1931_;
	assign _1933_ = _1911_ & ~_1932_;
	assign _1934_ = _1909_ & ~_1933_;
	assign _1935_ = _1929_ ^ _1928_;
	assign _1936_ = _1935_ | ~_1921_;
	assign _1937_ = _1911_ & ~_1936_;
	assign _1938_ = _1648_ ^ _1615_;
	assign _1939_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1884_ : _1938_);
	assign _1940_ = (_1150_ ? _1830_ : _1939_);
	assign _1941_ = (_1102_ ? _1655_ : _1940_);
	assign _1942_ = _1941_ ^ _1783_;
	assign _1943_ = ~(_1499_ | _1479_);
	assign _1944_ = _1943_ | ~_1476_;
	assign _1945_ = _1944_ ^ _1469_;
	assign _1946_ = _1942_ | ~_1945_;
	assign _1947_ = ~(_1945_ ^ _1942_);
	assign _1948_ = ~(_1646_ | _1632_);
	assign _1949_ = _1628_ & ~_1948_;
	assign _1950_ = ~(_1949_ ^ _1623_);
	assign _1951_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1901_ : _1950_);
	assign _1952_ = (_1150_ ? _1846_ : _1951_);
	assign _1953_ = (_1102_ ? _1655_ : _1952_);
	assign _1954_ = _1953_ ^ _1783_;
	assign _1955_ = _1499_ ^ _1479_;
	assign _1956_ = _1954_ | ~_1955_;
	assign _1957_ = _1947_ & ~_1956_;
	assign _1958_ = _1946_ & ~_1957_;
	assign _1959_ = _1955_ ^ _1954_;
	assign _1960_ = _1947_ & ~_1959_;
	assign _1961_ = _1646_ ^ _1632_;
	assign _1962_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1912_ : _1961_);
	assign _1963_ = (_1150_ ? _1857_ : _1962_);
	assign _1964_ = (_1102_ ? _1655_ : _1963_);
	assign _1965_ = _1964_ ^ _1783_;
	assign _1966_ = ~(_1497_ ^ _1489_);
	assign _1967_ = ~_1966_;
	assign _1968_ = _1967_ | _1965_;
	assign _1969_ = _1967_ ^ _1965_;
	assign _1970_ = _1496_ ^ _1491_;
	assign _1971_ = _1970_ ^ _1490_;
	assign _1972_ = _1971_ ^ _1517_;
	assign _1973_ = ~_1972_;
	assign _1974_ = ~_1655_;
	assign _1975_ = ~_1150_;
	assign _1976_ = ~(_1644_ ^ _1639_);
	assign _1977_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1924_ : _1976_);
	assign _1978_ = _1975_ & ~_1977_;
	assign _1979_ = _1150_ & ~_1869_;
	assign _1980_ = _1979_ | _1978_;
	assign _1981_ = (_1102_ ? _1974_ : _1980_);
	assign _1982_ = (_1981_ ? _1783_ : _1973_);
	assign _1983_ = _1969_ & ~_1982_;
	assign _1984_ = _1968_ & ~_1983_;
	assign _1985_ = _1960_ & ~_1984_;
	assign _1986_ = _1958_ & ~_1985_;
	assign _1987_ = _1937_ & ~_1986_;
	assign _1988_ = _1934_ & ~_1987_;
	assign _1989_ = _1873_ ^ _1872_;
	assign _1990_ = _1989_ | ~_1865_;
	assign _1991_ = _1855_ & ~_1990_;
	assign _1992_ = _1881_ | ~_1991_;
	assign _1993_ = ~(_1992_ | _1988_);
	assign _1994_ = _1883_ & ~_1993_;
	assign _1995_ = _1784_ ^ _1782_;
	assign _1996_ = ~(_1995_ ^ _1994_);
	assign _1997_ = ~_1996_;
	assign _1998_ = ~_1783_;
	assign _1999_ = _1713_ & ~_1763_;
	assign _2000_ = _1708_ & ~_1999_;
	assign _2001_ = _1679_ & ~_2000_;
	assign _2002_ = _1675_ & ~_2001_;
	assign _2003_ = _1666_ & ~_2002_;
	assign _2004_ = _1663_ & ~_2003_;
	assign _2005_ = _2004_ ^ _1658_;
	assign _2006_ = _2005_ & ~_1998_;
	assign _2007_ = _2005_ ^ _1998_;
	assign _2008_ = ~(_2002_ ^ _1666_);
	assign _2009_ = ~(_2008_ & _1783_);
	assign _2010_ = ~(_2009_ | _2007_);
	assign _2011_ = ~(_2010_ | _2006_);
	assign _2012_ = _2008_ ^ _1783_;
	assign _2013_ = _2012_ & ~_2007_;
	assign _2014_ = ~(_2000_ | _1678_);
	assign _2015_ = _1672_ & ~_2014_;
	assign _2016_ = ~(_2015_ ^ _1673_);
	assign _2017_ = ~_1660_;
	assign _2018_ = _1783_ ^ _2017_;
	assign _2019_ = ~(_2018_ & _2016_);
	assign _2020_ = _2000_ ^ _1678_;
	assign _2021_ = _2020_ & _2018_;
	assign _2022_ = _2018_ ^ _2016_;
	assign _2023_ = _2022_ & _2021_;
	assign _2024_ = _2019_ & ~_2023_;
	assign _2025_ = _2013_ & ~_2024_;
	assign _2026_ = _2011_ & ~_2025_;
	assign _2027_ = ~(_2020_ ^ _2018_);
	assign _2028_ = _2022_ & ~_2027_;
	assign _2029_ = _2028_ & _2013_;
	assign _2030_ = ~(_1763_ | _1712_);
	assign _2031_ = _1706_ & ~_2030_;
	assign _2032_ = ~(_2031_ | _1694_);
	assign _2033_ = _1691_ & ~_2032_;
	assign _2034_ = ~(_2033_ ^ _1683_);
	assign _2035_ = ~(_2034_ & _2018_);
	assign _2036_ = _2031_ ^ _1694_;
	assign _2037_ = ~_2036_;
	assign _2038_ = _1783_ ^ _1698_;
	assign _2039_ = _2038_ & ~_2037_;
	assign _2040_ = _2034_ ^ _2018_;
	assign _2041_ = _2040_ & _2039_;
	assign _2042_ = _2035_ & ~_2041_;
	assign _2043_ = _2038_ ^ _2037_;
	assign _2044_ = _2040_ & ~_2043_;
	assign _2045_ = ~(_1763_ | _1711_);
	assign _2046_ = _1704_ & ~_2045_;
	assign _2047_ = ~(_2046_ ^ _1702_);
	assign _2048_ = ~(_2047_ & _2018_);
	assign _2049_ = _1763_ ^ _1711_;
	assign _2050_ = _2049_ & _2018_;
	assign _2051_ = _2047_ ^ _2018_;
	assign _2052_ = _2051_ & _2050_;
	assign _2053_ = _2048_ & ~_2052_;
	assign _2054_ = _2044_ & ~_2053_;
	assign _2055_ = _2042_ & ~_2054_;
	assign _2056_ = _2029_ & ~_2055_;
	assign _2057_ = _2026_ & ~_2056_;
	assign _2058_ = ~(_2049_ ^ _2018_);
	assign _2059_ = _2058_ | ~_2051_;
	assign _2060_ = _2044_ & ~_2059_;
	assign _2061_ = _2060_ & _2029_;
	assign _2062_ = _1738_ & ~_1761_;
	assign _2063_ = _1734_ & ~_2062_;
	assign _2064_ = _1726_ & ~_2063_;
	assign _2065_ = _1723_ & ~_2064_;
	assign _2066_ = _2065_ ^ _1721_;
	assign _2067_ = ~(_2066_ & _1783_);
	assign _2068_ = ~(_2066_ ^ _1783_);
	assign _2069_ = _2063_ ^ _1726_;
	assign _2070_ = _1660_ & ~_1715_;
	assign _2071_ = _1697_ & ~_2070_;
	assign _2072_ = _2071_ ^ _1783_;
	assign _2073_ = _2069_ | ~_2072_;
	assign _2074_ = ~(_2073_ | _2068_);
	assign _2075_ = _2067_ & ~_2074_;
	assign _2076_ = ~(_2072_ ^ _2069_);
	assign _2077_ = _2076_ & ~_2068_;
	assign _2078_ = ~(_1761_ | _1737_);
	assign _2079_ = _1732_ & ~_2078_;
	assign _2080_ = ~(_2079_ ^ _1730_);
	assign _2081_ = ~(_2080_ & _1783_);
	assign _2082_ = _2080_ ^ _1783_;
	assign _2083_ = _1761_ ^ _1737_;
	assign _2084_ = ~(_2083_ & _2018_);
	assign _2085_ = _2082_ & ~_2084_;
	assign _2086_ = _2081_ & ~_2085_;
	assign _2087_ = _2077_ & ~_2086_;
	assign _2088_ = _2075_ & ~_2087_;
	assign _2089_ = ~(_2083_ ^ _2018_);
	assign _2090_ = _2082_ & ~_2089_;
	assign _2091_ = _2090_ & _2077_;
	assign _2092_ = ~_1750_;
	assign _2093_ = _2092_ & ~_1759_;
	assign _2094_ = _1747_ & ~_2093_;
	assign _2095_ = ~(_2094_ ^ _1745_);
	assign _2096_ = ~(_2095_ & _2018_);
	assign _2097_ = ~(_2095_ ^ _2018_);
	assign _2098_ = _1759_ ^ _2092_;
	assign _2099_ = _0957_ & _0946_;
	assign _2100_ = _2099_ ^ _1783_;
	assign _2101_ = _2098_ | ~_2100_;
	assign _2102_ = ~(_2101_ | _2097_);
	assign _2103_ = _2096_ & ~_2102_;
	assign _2104_ = ~(_2100_ ^ _2098_);
	assign _2105_ = _2104_ & ~_2097_;
	assign _2106_ = _1757_ ^ _1754_;
	assign _2107_ = ~(_2106_ & _1783_);
	assign _2108_ = ~(_2106_ ^ _1783_);
	assign _2109_ = _1755_ ^ _1699_;
	assign _2110_ = _2109_ ^ _1491_;
	assign _2111_ = (_1660_ ? _1783_ : _2110_);
	assign _2112_ = _2111_ & ~_2108_;
	assign _2113_ = _2107_ & ~_2112_;
	assign _2114_ = _2105_ & ~_2113_;
	assign _2115_ = _2103_ & ~_2114_;
	assign _2116_ = _2091_ & ~_2115_;
	assign _2117_ = _2088_ & ~_2116_;
	assign _2118_ = _2061_ & ~_2117_;
	assign _2119_ = _2057_ & ~_2118_;
	assign _2120_ = ~(_1783_ ^ _1767_);
	assign _2121_ = ~(_2120_ ^ _2119_);
	assign _2122_ = (io_in[10] ? _1997_ : _2121_);
	assign _2123_ = _2122_ ^ _1996_;
	assign _2124_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1782_ : _1510_);
	assign _2125_ = (_1150_ ? _1782_ : _2124_);
	assign _2126_ = (_1102_ ? _1782_ : _2125_);
	assign _2127_ = _2126_ ^ _1783_;
	assign _2128_ = _2127_ & _1803_;
	assign _2129_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1782_ : _1798_);
	assign _2130_ = (_1150_ ? _1782_ : _2129_);
	assign _2131_ = (_1102_ ? _1782_ : _2130_);
	assign _2132_ = ~(_2131_ ^ _1783_);
	assign _2133_ = _1815_ & ~_2132_;
	assign _0119_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1782_ : _1810_);
	assign _0120_ = (_1150_ ? _1782_ : _0119_);
	assign _0121_ = (_1102_ ? _1782_ : _0120_);
	assign _0122_ = _0121_ ^ _1783_;
	assign _0123_ = _0122_ & _1829_;
	assign _0124_ = _2132_ ^ _1815_;
	assign _0125_ = _0123_ & ~_0124_;
	assign _0126_ = _0125_ | _2133_;
	assign _0127_ = ~(_0122_ ^ _1829_);
	assign _0128_ = ~(_0127_ | _0124_);
	assign _0129_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1820_ : _1873_);
	assign _0130_ = (_1150_ ? _1782_ : _0129_);
	assign _0131_ = (_1102_ ? _1782_ : _0130_);
	assign _0132_ = _0131_ ^ _1783_;
	assign _0133_ = _0132_ & _1901_;
	assign _0134_ = ~(_0132_ ^ _1901_);
	assign _0135_ = ~_0134_;
	assign _0136_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1838_ : _1893_);
	assign _0137_ = (_1150_ ? _2124_ : _0136_);
	assign _0138_ = (_1102_ ? _1782_ : _0137_);
	assign _0139_ = _0138_ ^ _1783_;
	assign _0140_ = ~(_0139_ & _1912_);
	assign _0141_ = _0135_ & ~_0140_;
	assign _0142_ = _0141_ | _0133_;
	assign _0143_ = ~(_0139_ ^ _1912_);
	assign _0144_ = _0135_ & ~_0143_;
	assign _0145_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1850_ : _1906_);
	assign _0146_ = (_1150_ ? _2129_ : _0145_);
	assign _0147_ = (_1102_ ? _1782_ : _0146_);
	assign _0148_ = _0147_ ^ _1783_;
	assign _0149_ = ~(_0148_ & _1924_);
	assign _0150_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1863_ : _1919_);
	assign _0151_ = (_1150_ ? _0119_ : _0150_);
	assign _0152_ = (_1102_ ? _1782_ : _0151_);
	assign _0153_ = ~(_0152_ ^ _1783_);
	assign _0154_ = _1938_ & ~_0153_;
	assign _0155_ = ~(_0148_ ^ _1924_);
	assign _0156_ = _0154_ & ~_0155_;
	assign _0157_ = _0149_ & ~_0156_;
	assign _0158_ = _0144_ & ~_0157_;
	assign _0159_ = _0158_ | _0142_;
	assign _0160_ = _0153_ ^ _1938_;
	assign _0161_ = _0160_ | _0155_;
	assign _0162_ = _0144_ & ~_0161_;
	assign _0163_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1873_ : _1929_);
	assign _0164_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1782_ : _1820_);
	assign _0165_ = (_1150_ ? _0164_ : _0163_);
	assign _0166_ = (_1102_ ? _1782_ : _0165_);
	assign _0167_ = _0166_ ^ _1783_;
	assign _0168_ = ~(_0167_ & _1950_);
	assign _0169_ = _0167_ ^ _1950_;
	assign _0170_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1893_ : _1945_);
	assign _0171_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1510_ : _1838_);
	assign _0172_ = (_1150_ ? _0171_ : _0170_);
	assign _0173_ = (_1102_ ? _1782_ : _0172_);
	assign _0174_ = _0173_ ^ _1783_;
	assign _0175_ = ~(_0174_ & _1961_);
	assign _0176_ = _0169_ & ~_0175_;
	assign _0177_ = _0168_ & ~_0176_;
	assign _0178_ = ~(_0174_ ^ _1961_);
	assign _0179_ = _0169_ & ~_0178_;
	assign _0180_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1906_ : _1955_);
	assign _0181_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1798_ : _1850_);
	assign _0182_ = (_1150_ ? _0181_ : _0180_);
	assign _0183_ = (_1102_ ? _1782_ : _0182_);
	assign _0184_ = _0183_ ^ _1783_;
	assign _0185_ = ~(_0184_ & _1976_);
	assign _0186_ = _0184_ ^ _1976_;
	assign _0187_ = _1642_ ^ _1517_;
	assign _0188_ = _0187_ ^ _1493_;
	assign _0189_ = _0188_ ^ _1491_;
	assign _0190_ = ~_0189_;
	assign _0191_ = ~_1782_;
	assign _0192_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1919_ : _1966_);
	assign _0193_ = _1975_ & ~_0192_;
	assign _0194_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1810_ : _1863_);
	assign _0195_ = _1150_ & ~_0194_;
	assign _0196_ = _0195_ | _0193_;
	assign _0197_ = (_1102_ ? _0191_ : _0196_);
	assign _0198_ = (_0197_ ? _1998_ : _0190_);
	assign _0199_ = _0186_ & ~_0198_;
	assign _0200_ = _0185_ & ~_0199_;
	assign _0201_ = _0179_ & ~_0200_;
	assign _0202_ = _0177_ & ~_0201_;
	assign _0203_ = _0162_ & ~_0202_;
	assign _0204_ = _0203_ | _0159_;
	assign _0205_ = (_1150_ ? _1782_ : _0194_);
	assign _0206_ = (_1102_ ? _1782_ : _0205_);
	assign _0207_ = ~(_0206_ ^ _1783_);
	assign _0208_ = ~(_0207_ ^ _1884_);
	assign _0209_ = (_1150_ ? _1782_ : _0181_);
	assign _0210_ = (_1102_ ? _1782_ : _0209_);
	assign _0211_ = ~(_0210_ ^ _1783_);
	assign _0212_ = _0211_ ^ _1868_;
	assign _0213_ = _0212_ | ~_0208_;
	assign _0214_ = (_1150_ ? _1782_ : _0171_);
	assign _0215_ = (_1102_ ? _1782_ : _0214_);
	assign _0216_ = ~(_0215_ ^ _1783_);
	assign _0217_ = _0216_ ^ _1856_;
	assign _0218_ = (_1150_ ? _1782_ : _0164_);
	assign _0219_ = (_1102_ ? _1782_ : _0218_);
	assign _0220_ = _0219_ ^ _1783_;
	assign _0221_ = ~(_0220_ ^ _1845_);
	assign _0222_ = _0221_ | _0217_;
	assign _0223_ = _0222_ | _0213_;
	assign _0224_ = _0223_ | ~_0204_;
	assign _0225_ = _1868_ & ~_0211_;
	assign _0226_ = _1884_ & ~_0207_;
	assign _0227_ = _0226_ & ~_0212_;
	assign _0228_ = _0227_ | _0225_;
	assign _0229_ = _0228_ & ~_0222_;
	assign _0230_ = _0220_ & _1845_;
	assign _0231_ = _1856_ & ~_0216_;
	assign _0232_ = _0231_ & ~_0221_;
	assign _0233_ = _0232_ | _0230_;
	assign _0234_ = _0233_ | _0229_;
	assign _0235_ = _0224_ & ~_0234_;
	assign _0236_ = _0128_ & ~_0235_;
	assign _0237_ = _0236_ | _0126_;
	assign _0238_ = _2127_ ^ _1803_;
	assign _0239_ = ~_0238_;
	assign _0240_ = _0237_ & ~_0239_;
	assign _0241_ = _0240_ | _2128_;
	assign _0242_ = _1783_ ^ _1782_;
	assign _0243_ = _0242_ ^ _1793_;
	assign _0244_ = _0243_ ^ _0241_;
	assign _0245_ = _0244_ & ~_2123_;
	assign _0246_ = _0238_ ^ _0237_;
	assign _0247_ = _0246_ & ~_2123_;
	assign _0248_ = _0244_ ^ _2123_;
	assign _0249_ = _0247_ & ~_0248_;
	assign _0250_ = ~(_0249_ | _0245_);
	assign _0251_ = _0246_ ^ _2123_;
	assign _0252_ = ~(_0251_ | _0248_);
	assign _0253_ = ~_2122_;
	assign _0254_ = _1991_ & ~_1988_;
	assign _0255_ = _1878_ & ~_0254_;
	assign _0256_ = _1880_ & ~_0255_;
	assign _0257_ = _1824_ & ~_0256_;
	assign _0258_ = _1825_ & ~_0257_;
	assign _0259_ = ~(_0258_ | _1799_);
	assign _0260_ = _1800_ ^ _0259_;
	assign _0261_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1996_ : _0260_);
	assign _0262_ = (_1150_ ? _1996_ : _0261_);
	assign _0263_ = (_1102_ ? _1996_ : _0262_);
	assign _0264_ = ~(_0263_ ^ _0253_);
	assign _0265_ = _0235_ | _0127_;
	assign _0266_ = _0265_ & ~_0123_;
	assign _0267_ = _0266_ ^ _0124_;
	assign _0268_ = _0264_ | ~_0267_;
	assign _0269_ = ~(_0257_ ^ _1825_);
	assign _0270_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1996_ : _0269_);
	assign _0271_ = (_1150_ ? _1996_ : _0270_);
	assign _0272_ = (_1102_ ? _1996_ : _0271_);
	assign _0273_ = _0272_ ^ _0253_;
	assign _0274_ = _0235_ ^ _0127_;
	assign _0275_ = _0274_ & _0273_;
	assign _0276_ = _0267_ ^ _0264_;
	assign _0277_ = _0275_ & ~_0276_;
	assign _0278_ = _0268_ & ~_0277_;
	assign _0279_ = _0252_ & ~_0278_;
	assign _0280_ = _0250_ & ~_0279_;
	assign _0281_ = ~(_1988_ | _1990_);
	assign _0282_ = _1876_ & ~_0281_;
	assign _0283_ = ~(_0282_ | _1854_);
	assign _0284_ = _1851_ & ~_0283_;
	assign _0285_ = ~(_0284_ ^ _1840_);
	assign _0286_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0260_ : _0285_);
	assign _0287_ = (_1150_ ? _1996_ : _0286_);
	assign _0288_ = (_1102_ ? _1996_ : _0287_);
	assign _0289_ = _0253_ ^ _0288_;
	assign _0290_ = _0208_ & _0204_;
	assign _0291_ = ~(_0290_ | _0226_);
	assign _0292_ = _0212_ ^ _0291_;
	assign _0293_ = ~(_0292_ & _0289_);
	assign _0294_ = ~(_0292_ ^ _0289_);
	assign _0295_ = ~_0269_;
	assign _0296_ = _0282_ ^ _1854_;
	assign _0297_ = ~_0296_;
	assign _0298_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0295_ : _0297_);
	assign _0299_ = (_1150_ ? _1997_ : _0298_);
	assign _0300_ = (_1102_ ? _1997_ : _0299_);
	assign _0301_ = _0300_ ^ _0253_;
	assign _0302_ = _0208_ ^ _0204_;
	assign _0303_ = _0301_ | ~_0302_;
	assign _0304_ = ~(_0303_ | _0294_);
	assign _0305_ = _0304_ | ~_0293_;
	assign _0306_ = _0255_ ^ _1879_;
	assign _0307_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1996_ : _0306_);
	assign _0308_ = (_1150_ ? _1996_ : _0307_);
	assign _0309_ = (_1102_ ? _1996_ : _0308_);
	assign _0310_ = _0309_ ^ _0253_;
	assign _0311_ = _0204_ & ~_0213_;
	assign _0312_ = _0311_ | _0228_;
	assign _0313_ = ~(_0217_ ^ _0312_);
	assign _0314_ = _0313_ ^ _0310_;
	assign _0315_ = _0255_ | _1879_;
	assign _0316_ = _0315_ & ~_1821_;
	assign _0317_ = _0316_ ^ _1822_;
	assign _0318_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1996_ : _0317_);
	assign _0319_ = (_1150_ ? _1996_ : _0318_);
	assign _0320_ = (_1102_ ? _1996_ : _0319_);
	assign _0321_ = _0320_ ^ _0253_;
	assign _0322_ = _0312_ & ~_0217_;
	assign _0323_ = ~(_0322_ | _0231_);
	assign _0324_ = _0323_ ^ _0221_;
	assign _0325_ = ~(_0324_ ^ _0321_);
	assign _0326_ = _0325_ | ~_0314_;
	assign _0327_ = _0326_ | ~_0305_;
	assign _0328_ = ~_0313_;
	assign _0329_ = _0310_ & ~_0328_;
	assign _0330_ = _0329_ & ~_0325_;
	assign _0331_ = _0324_ & _0321_;
	assign _0332_ = _0331_ | _0330_;
	assign _0333_ = _0327_ & ~_0332_;
	assign _0334_ = ~(_0274_ ^ _0273_);
	assign _0335_ = ~(_0334_ | _0276_);
	assign _0336_ = ~(_0335_ & _0252_);
	assign _0337_ = ~(_0336_ | _0333_);
	assign _0338_ = _0280_ & ~_0337_;
	assign _0339_ = ~(_1988_ | _1989_);
	assign _0340_ = _1874_ & ~_0339_;
	assign _0341_ = ~(_0340_ ^ _1865_);
	assign _0342_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0317_ : _0341_);
	assign _0343_ = (_1150_ ? _1996_ : _0342_);
	assign _0344_ = (_1102_ ? _1996_ : _0343_);
	assign _0345_ = _0344_ ^ _0253_;
	assign _0346_ = ~(_0202_ | _0161_);
	assign _0347_ = _0157_ & ~_0346_;
	assign _0348_ = ~(_0347_ | _0143_);
	assign _0349_ = _0140_ & ~_0348_;
	assign _0350_ = _0349_ ^ _0134_;
	assign _0351_ = _0350_ & _0345_;
	assign _0352_ = _0350_ ^ _0345_;
	assign _0353_ = _1988_ ^ _1989_;
	assign _0354_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0306_ : _0353_);
	assign _0355_ = (_1150_ ? _1996_ : _0354_);
	assign _0356_ = (_1102_ ? _1996_ : _0355_);
	assign _0357_ = ~(_0356_ ^ _0253_);
	assign _0358_ = _0347_ ^ _0143_;
	assign _0359_ = _0357_ | ~_0358_;
	assign _0360_ = _0352_ & ~_0359_;
	assign _0361_ = _0360_ | _0351_;
	assign _0362_ = ~(_0358_ ^ _0357_);
	assign _0363_ = ~_0362_;
	assign _0364_ = _0352_ & ~_0363_;
	assign _0365_ = ~(_1986_ | _1936_);
	assign _0366_ = _1932_ & ~_0365_;
	assign _0367_ = ~(_0366_ | _1910_);
	assign _0368_ = _1907_ & ~_0367_;
	assign _0369_ = _0368_ ^ _1895_;
	assign _0370_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0285_ : _0369_);
	assign _0371_ = (_1150_ ? _0261_ : _0370_);
	assign _0372_ = (_1102_ ? _1996_ : _0371_);
	assign _0373_ = ~(_0372_ ^ _0253_);
	assign _0374_ = _0202_ | _0160_;
	assign _0375_ = _0374_ & ~_0154_;
	assign _0376_ = _0375_ ^ _0155_;
	assign _0377_ = _0373_ | ~_0376_;
	assign _0378_ = ~(_0376_ ^ _0373_);
	assign _0379_ = _0366_ ^ _1910_;
	assign _0380_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0296_ : _0379_);
	assign _0381_ = (_1150_ ? _0270_ : _0380_);
	assign _0382_ = (_1102_ ? _1996_ : _0381_);
	assign _0383_ = ~(_0382_ ^ _0253_);
	assign _0384_ = _0202_ ^ _0160_;
	assign _0385_ = _0383_ | ~_0384_;
	assign _0386_ = _0378_ & ~_0385_;
	assign _0387_ = _0377_ & ~_0386_;
	assign _0388_ = _0364_ & ~_0387_;
	assign _0389_ = _0388_ | _0361_;
	assign _0390_ = _0384_ ^ _0383_;
	assign _0391_ = _0390_ | ~_0378_;
	assign _0392_ = _0364_ & ~_0391_;
	assign _0393_ = ~(_1986_ | _1935_);
	assign _0394_ = _0393_ | ~_1930_;
	assign _0395_ = _0394_ ^ _1921_;
	assign _0396_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0341_ : _0395_);
	assign _0397_ = (_1150_ ? _0318_ : _0396_);
	assign _0398_ = (_1102_ ? _1996_ : _0397_);
	assign _0399_ = ~(_0398_ ^ _0253_);
	assign _0400_ = ~(_0200_ | _0178_);
	assign _0401_ = _0400_ | ~_0175_;
	assign _0402_ = _0401_ ^ _0169_;
	assign _0403_ = _0399_ | ~_0402_;
	assign _0404_ = ~(_0402_ ^ _0399_);
	assign _0405_ = _1986_ ^ _1935_;
	assign _0406_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0353_ : _0405_);
	assign _0407_ = (_1150_ ? _0307_ : _0406_);
	assign _0408_ = (_1102_ ? _1996_ : _0407_);
	assign _0409_ = ~(_0408_ ^ _0253_);
	assign _0410_ = _0200_ ^ _0178_;
	assign _0411_ = _0409_ | ~_0410_;
	assign _0412_ = _0404_ & ~_0411_;
	assign _0413_ = _0403_ & ~_0412_;
	assign _0414_ = ~(_0410_ ^ _0409_);
	assign _0415_ = ~_0414_;
	assign _0416_ = _0404_ & ~_0415_;
	assign _0417_ = ~(_0198_ ^ _0186_);
	assign _0418_ = ~(_1984_ | _1959_);
	assign _0419_ = _1956_ & ~_0418_;
	assign _0420_ = ~(_0419_ ^ _1947_);
	assign _0421_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0369_ : _0420_);
	assign _0422_ = (_1150_ ? _0286_ : _0421_);
	assign _0423_ = (_1102_ ? _1996_ : _0422_);
	assign _0424_ = _0423_ ^ _0253_;
	assign _0425_ = ~(_0424_ & _0417_);
	assign _0426_ = _0424_ ^ _0417_;
	assign _0427_ = _0197_ ^ _1783_;
	assign _0428_ = _0427_ ^ _0190_;
	assign _0429_ = _0428_ ^ _1783_;
	assign _0430_ = ~_0429_;
	assign _0431_ = _1984_ ^ _1959_;
	assign _0432_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0379_ : _0431_);
	assign _0433_ = ~_0432_;
	assign _0434_ = (_1150_ ? _0298_ : _0433_);
	assign _0435_ = (_1102_ ? _1997_ : _0434_);
	assign _0436_ = (_0435_ ? _2122_ : _0430_);
	assign _0437_ = _0426_ & ~_0436_;
	assign _0438_ = _0425_ & ~_0437_;
	assign _0439_ = _0416_ & ~_0438_;
	assign _0440_ = _0413_ & ~_0439_;
	assign _0441_ = _0392_ & ~_0440_;
	assign _0442_ = _0441_ | _0389_;
	assign _0443_ = ~(_0302_ ^ _0301_);
	assign _0444_ = ~_0443_;
	assign _0445_ = _0444_ | _0294_;
	assign _0446_ = _0326_ | _0445_;
	assign _0447_ = _0446_ | _0336_;
	assign _0448_ = _0442_ & ~_0447_;
	assign _0449_ = _0338_ & ~_0448_;
	assign _0450_ = _0242_ & _1793_;
	assign _0451_ = _0243_ & _2128_;
	assign _0452_ = ~(_0451_ | _0450_);
	assign _0453_ = ~(_0243_ & _0238_);
	assign _0454_ = _0126_ & ~_0453_;
	assign _0455_ = _0452_ & ~_0454_;
	assign _0456_ = _0453_ | ~_0128_;
	assign _0457_ = _0234_ & ~_0456_;
	assign _0458_ = _0455_ & ~_0457_;
	assign _0459_ = _0456_ | _0223_;
	assign _0460_ = _0204_ & ~_0459_;
	assign _0461_ = _0458_ & ~_0460_;
	assign _0462_ = ~(_0242_ ^ _1655_);
	assign _0463_ = _0462_ ^ _0461_;
	assign _0464_ = _0463_ ^ _2123_;
	assign _0465_ = _0464_ ^ _0449_;
	assign _0466_ = _0442_ & ~_0445_;
	assign _0467_ = _0466_ | _0305_;
	assign _0468_ = _0314_ ^ _0467_;
	assign _0469_ = ~(_0440_ | _0391_);
	assign _0470_ = _0387_ & ~_0469_;
	assign _0471_ = _0470_ ^ _0363_;
	assign _0472_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0468_ : _0471_);
	assign _0473_ = _0442_ & ~_0446_;
	assign _0474_ = _0333_ & ~_0473_;
	assign _0475_ = _0335_ & ~_0474_;
	assign _0476_ = _0278_ & ~_0475_;
	assign _0477_ = _0476_ ^ _0251_;
	assign _0478_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0465_ : _0477_);
	assign _0479_ = (_1150_ ? _0478_ : _0472_);
	assign _0480_ = (_1102_ ? _0465_ : _0479_);
	assign _0481_ = _2060_ & ~_2117_;
	assign _0482_ = _2055_ & ~_0481_;
	assign _0483_ = _2028_ & ~_0482_;
	assign _0484_ = _2024_ & ~_0483_;
	assign _0485_ = _2012_ & ~_0484_;
	assign _0486_ = _2009_ & ~_0485_;
	assign _0487_ = _0486_ ^ _2007_;
	assign _0488_ = _0487_ & ~_2122_;
	assign _0489_ = _0487_ ^ _2122_;
	assign _0490_ = ~(_0484_ ^ _2012_);
	assign _0491_ = _2122_ | ~_0490_;
	assign _0492_ = ~(_0491_ | _0489_);
	assign _0493_ = ~(_0492_ | _0488_);
	assign _0494_ = ~(_0490_ ^ _2122_);
	assign _0495_ = _0494_ & ~_0489_;
	assign _0496_ = _0482_ | _2027_;
	assign _0497_ = _0496_ & ~_2021_;
	assign _0498_ = ~(_0497_ ^ _2022_);
	assign _0499_ = _2122_ | ~_0498_;
	assign _0500_ = ~(_0498_ ^ _2122_);
	assign _0501_ = ~(_0482_ ^ _2027_);
	assign _0502_ = _2122_ ^ _1660_;
	assign _0503_ = _0501_ | ~_0502_;
	assign _0504_ = _0500_ & ~_0503_;
	assign _0505_ = _0499_ & ~_0504_;
	assign _0506_ = _0495_ & ~_0505_;
	assign _0507_ = _0493_ & ~_0506_;
	assign _0508_ = _0502_ ^ _0501_;
	assign _0509_ = _0500_ & ~_0508_;
	assign _0510_ = _0509_ & _0495_;
	assign _0511_ = ~(_2117_ | _2059_);
	assign _0512_ = _2053_ & ~_0511_;
	assign _0513_ = _0512_ | _2043_;
	assign _0514_ = _0513_ & ~_2039_;
	assign _0515_ = ~(_0514_ ^ _2040_);
	assign _0516_ = ~(_0515_ & _0502_);
	assign _0517_ = _0512_ ^ _2043_;
	assign _0518_ = _0517_ & _0502_;
	assign _0519_ = _0515_ ^ _0502_;
	assign _0520_ = _0519_ & _0518_;
	assign _0521_ = _0516_ & ~_0520_;
	assign _0522_ = ~(_0517_ ^ _0502_);
	assign _0523_ = _0519_ & ~_0522_;
	assign _0524_ = _2117_ | _2058_;
	assign _0525_ = _0524_ & ~_2050_;
	assign _0526_ = _0525_ ^ _2051_;
	assign _0527_ = ~(_2122_ ^ _1688_);
	assign _0528_ = _0526_ | ~_0527_;
	assign _0529_ = _2117_ ^ _2058_;
	assign _0530_ = _0529_ & _0502_;
	assign _0531_ = ~(_0527_ ^ _0526_);
	assign _0532_ = _0531_ & _0530_;
	assign _0533_ = _0528_ & ~_0532_;
	assign _0534_ = _0523_ & ~_0533_;
	assign _0535_ = _0521_ & ~_0534_;
	assign _0536_ = _0510_ & ~_0535_;
	assign _0537_ = _0507_ & ~_0536_;
	assign _0538_ = ~(_0529_ ^ _0502_);
	assign _0539_ = _0538_ | ~_0531_;
	assign _0540_ = _0523_ & ~_0539_;
	assign _0541_ = _0540_ & _0510_;
	assign _0542_ = _2090_ & ~_2115_;
	assign _0543_ = _2086_ & ~_0542_;
	assign _0544_ = _2076_ & ~_0543_;
	assign _0545_ = _2073_ & ~_0544_;
	assign _0546_ = _0545_ ^ _2068_;
	assign _0547_ = _2122_ | ~_0546_;
	assign _0548_ = _0546_ ^ _2122_;
	assign _0549_ = ~(_0543_ ^ _2076_);
	assign _0550_ = ~(_0549_ & _0502_);
	assign _0551_ = ~(_0550_ | _0548_);
	assign _0552_ = _0547_ & ~_0551_;
	assign _0553_ = _0549_ ^ _0502_;
	assign _0554_ = _0553_ & ~_0548_;
	assign _0555_ = ~(_2115_ | _2089_);
	assign _0556_ = _2084_ & ~_0555_;
	assign _0557_ = ~(_0556_ ^ _2082_);
	assign _0558_ = _1715_ & _1697_;
	assign _0559_ = ~(_0558_ ^ _2122_);
	assign _0560_ = ~(_0559_ & _0557_);
	assign _0561_ = _2115_ ^ _2089_;
	assign _0562_ = _0561_ & _0502_;
	assign _0563_ = _0559_ ^ _0557_;
	assign _0564_ = _0563_ & _0562_;
	assign _0565_ = _0560_ & ~_0564_;
	assign _0566_ = _0554_ & ~_0565_;
	assign _0567_ = _0552_ & ~_0566_;
	assign _0568_ = ~(_0561_ ^ _0502_);
	assign _0569_ = _0563_ & ~_0568_;
	assign _0570_ = _0569_ & _0554_;
	assign _0571_ = _2104_ & ~_2113_;
	assign _0572_ = _2101_ & ~_0571_;
	assign _0573_ = _0572_ ^ _2097_;
	assign _0574_ = ~(_0573_ & _0502_);
	assign _0575_ = ~(_0573_ ^ _0502_);
	assign _0576_ = ~(_2113_ ^ _2104_);
	assign _0577_ = _2122_ | ~_0576_;
	assign _0578_ = ~(_0577_ | _0575_);
	assign _0579_ = _0574_ & ~_0578_;
	assign _0580_ = ~(_0576_ ^ _2122_);
	assign _0581_ = _0580_ & ~_0575_;
	assign _0582_ = ~(_2111_ ^ _2108_);
	assign _0583_ = _1660_ & _0001_;
	assign _0584_ = _0583_ ^ _2122_;
	assign _0585_ = ~(_0584_ & _0582_);
	assign _0586_ = ~(_0584_ ^ _0582_);
	assign _0587_ = _2110_ ^ _2018_;
	assign _0588_ = _0587_ ^ _1783_;
	assign _0589_ = (_1660_ ? _0253_ : _0588_);
	assign _0590_ = _0589_ & ~_0586_;
	assign _0591_ = _0585_ & ~_0590_;
	assign _0592_ = _0581_ & ~_0591_;
	assign _0593_ = _0579_ & ~_0592_;
	assign _0594_ = _0570_ & ~_0593_;
	assign _0595_ = _0567_ & ~_0594_;
	assign _0596_ = _0541_ & ~_0595_;
	assign _0597_ = _0537_ & ~_0596_;
	assign _0598_ = ~(_2122_ ^ _2121_);
	assign _0599_ = ~(_0598_ ^ _0597_);
	assign _0600_ = ~_0599_;
	assign _0601_ = _0463_ ^ _2122_;
	assign _0602_ = _0601_ & _0260_;
	assign _0603_ = ~(_0601_ ^ _0260_);
	assign _0604_ = ~(_0601_ & _0269_);
	assign _0605_ = ~(_0604_ | _0603_);
	assign _0606_ = ~(_0605_ | _0602_);
	assign _0607_ = _0601_ ^ _0269_;
	assign _0608_ = _0607_ & ~_0603_;
	assign _0609_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0463_ : _0244_);
	assign _0610_ = (_1150_ ? _0463_ : _0609_);
	assign _0611_ = (_1102_ ? _0463_ : _0610_);
	assign _0612_ = ~(_0611_ ^ _0253_);
	assign _0613_ = ~(_0612_ & _0317_);
	assign _0614_ = _0612_ ^ _0317_;
	assign _0615_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0463_ : _0246_);
	assign _0616_ = (_1150_ ? _0463_ : _0615_);
	assign _0617_ = (_1102_ ? _0463_ : _0616_);
	assign _0618_ = ~(_0617_ ^ _0253_);
	assign _0619_ = ~(_0618_ & _0306_);
	assign _0620_ = _0614_ & ~_0619_;
	assign _0621_ = _0613_ & ~_0620_;
	assign _0622_ = _0608_ & ~_0621_;
	assign _0623_ = _0606_ & ~_0622_;
	assign _0624_ = ~(_0618_ ^ _0306_);
	assign _0625_ = _0614_ & ~_0624_;
	assign _0626_ = _0625_ & _0608_;
	assign _0627_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0463_ : _0267_);
	assign _0628_ = (_1150_ ? _0463_ : _0627_);
	assign _0629_ = (_1102_ ? _0463_ : _0628_);
	assign _0630_ = ~(_0629_ ^ _0253_);
	assign _0631_ = ~(_0630_ & _0285_);
	assign _0632_ = _0630_ ^ _0285_;
	assign _0633_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0463_ : _0274_);
	assign _0634_ = (_1150_ ? _0463_ : _0633_);
	assign _0635_ = (_1102_ ? _0463_ : _0634_);
	assign _0636_ = ~(_0635_ ^ _0253_);
	assign _0637_ = ~(_0636_ & _0296_);
	assign _0638_ = _0632_ & ~_0637_;
	assign _0639_ = _0631_ & ~_0638_;
	assign _0640_ = _0636_ ^ _0297_;
	assign _0641_ = _0632_ & ~_0640_;
	assign _0642_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0244_ : _0324_);
	assign _0643_ = (_1150_ ? _0463_ : _0642_);
	assign _0644_ = (_1102_ ? _0463_ : _0643_);
	assign _0645_ = ~(_0644_ ^ _0253_);
	assign _0646_ = ~(_0645_ & _0341_);
	assign _0647_ = _0645_ ^ _0341_;
	assign _0648_ = ~_0463_;
	assign _0649_ = ~_0246_;
	assign _0650_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0649_ : _0328_);
	assign _0651_ = (_1150_ ? _0648_ : _0650_);
	assign _0652_ = (_1102_ ? _0648_ : _0651_);
	assign _0653_ = _0652_ ^ _0253_;
	assign _0654_ = ~(_0653_ & _0353_);
	assign _0655_ = _0647_ & ~_0654_;
	assign _0656_ = _0646_ & ~_0655_;
	assign _0657_ = _0641_ & ~_0656_;
	assign _0658_ = _0639_ & ~_0657_;
	assign _0659_ = _0626_ & ~_0658_;
	assign _0660_ = _0659_ | ~_0623_;
	assign _0661_ = ~(_0653_ ^ _0353_);
	assign _0662_ = _0661_ | ~_0647_;
	assign _0663_ = _0641_ & ~_0662_;
	assign _0664_ = _0663_ & _0626_;
	assign _0665_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0267_ : _0292_);
	assign _0666_ = (_1150_ ? _0463_ : _0665_);
	assign _0667_ = (_1102_ ? _0463_ : _0666_);
	assign _0668_ = ~(_0667_ ^ _0253_);
	assign _0669_ = ~(_0668_ & _0369_);
	assign _0670_ = _0668_ ^ _0369_;
	assign _0671_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0274_ : _0302_);
	assign _0672_ = (_1150_ ? _0463_ : _0671_);
	assign _0673_ = (_1102_ ? _0463_ : _0672_);
	assign _0674_ = ~(_0673_ ^ _0253_);
	assign _0675_ = ~(_0674_ & _0379_);
	assign _0676_ = _0670_ & ~_0675_;
	assign _0677_ = _0669_ & ~_0676_;
	assign _0678_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0324_ : _0350_);
	assign _0679_ = (_1150_ ? _0609_ : _0678_);
	assign _0680_ = (_1102_ ? _0463_ : _0679_);
	assign _0681_ = _0680_ ^ _0253_;
	assign _0682_ = ~(_0681_ ^ _0395_);
	assign _0683_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0313_ : _0358_);
	assign _0684_ = (_1150_ ? _0615_ : _0683_);
	assign _0685_ = (_1102_ ? _0463_ : _0684_);
	assign _0686_ = ~(_0685_ ^ _0253_);
	assign _0687_ = ~(_0686_ & _0405_);
	assign _0688_ = _0682_ & ~_0687_;
	assign _0689_ = _0395_ & ~_0681_;
	assign _0690_ = _0689_ | _0688_;
	assign _0691_ = ~(_0674_ ^ _0379_);
	assign _0692_ = _0670_ & ~_0691_;
	assign _0693_ = _0692_ & _0690_;
	assign _0694_ = _0677_ & ~_0693_;
	assign _0695_ = ~(_0686_ ^ _0405_);
	assign _0696_ = _0695_ | ~_0682_;
	assign _0697_ = _0692_ & ~_0696_;
	assign _0698_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0292_ : _0376_);
	assign _0699_ = (_1150_ ? _0627_ : _0698_);
	assign _0700_ = (_1102_ ? _0463_ : _0699_);
	assign _0701_ = ~(_0700_ ^ _0253_);
	assign _0702_ = ~(_0701_ & _0420_);
	assign _0703_ = _0701_ ^ _0420_;
	assign _0704_ = ~_0431_;
	assign _0705_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0302_ : _0384_);
	assign _0706_ = (_1150_ ? _0633_ : _0705_);
	assign _0707_ = (_1102_ ? _0463_ : _0706_);
	assign _0708_ = ~(_0707_ ^ _0253_);
	assign _0709_ = _0704_ | ~_0708_;
	assign _0710_ = _0703_ & ~_0709_;
	assign _0711_ = _0702_ & ~_0710_;
	assign _0712_ = ~(_0708_ ^ _0704_);
	assign _0713_ = ~_0712_;
	assign _0714_ = _0703_ & ~_0713_;
	assign _0715_ = ~(_1982_ ^ _1969_);
	assign _0716_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0350_ : _0402_);
	assign _0717_ = (_1150_ ? _0642_ : _0716_);
	assign _0718_ = (_1102_ ? _0463_ : _0717_);
	assign _0719_ = ~(_0718_ ^ _0253_);
	assign _0720_ = ~(_0719_ & _0715_);
	assign _0721_ = _0719_ ^ _0715_;
	assign _0722_ = _1981_ ^ _1998_;
	assign _0723_ = _0722_ ^ _1973_;
	assign _0724_ = _0723_ ^ _1998_;
	assign _0725_ = ~_0724_;
	assign _0726_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0358_ : _0410_);
	assign _0727_ = ~_0726_;
	assign _0728_ = (_1150_ ? _0650_ : _0727_);
	assign _0729_ = (_1102_ ? _0648_ : _0728_);
	assign _0730_ = (_0729_ ? _0253_ : _0725_);
	assign _0731_ = _0721_ & ~_0730_;
	assign _0732_ = _0720_ & ~_0731_;
	assign _0733_ = _0714_ & ~_0732_;
	assign _0734_ = _0711_ & ~_0733_;
	assign _0735_ = _0697_ & ~_0734_;
	assign _0736_ = _0694_ & ~_0735_;
	assign _0737_ = _0664_ & ~_0736_;
	assign _0738_ = _0737_ | _0660_;
	assign _0739_ = _0601_ ^ _1996_;
	assign _0740_ = _0739_ ^ _0738_;
	assign _0741_ = (io_in[10] ? _0740_ : _0600_);
	assign _0742_ = ~(_0741_ ^ _0480_);
	assign _0743_ = _0712_ & ~_0732_;
	assign _0744_ = _0709_ & ~_0743_;
	assign _0745_ = ~(_0744_ ^ _0703_);
	assign _0746_ = ~_0745_;
	assign _0747_ = _0742_ & ~_0746_;
	assign _0748_ = _0745_ ^ _0742_;
	assign _0749_ = _0442_ & ~_0444_;
	assign _0750_ = _0303_ & ~_0749_;
	assign _0751_ = _0750_ ^ _0294_;
	assign _0752_ = ~(_0440_ | _0390_);
	assign _0753_ = _0385_ & ~_0752_;
	assign _0754_ = ~(_0753_ ^ _0378_);
	assign _0755_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0751_ : _0754_);
	assign _0756_ = _0474_ | _0334_;
	assign _0757_ = _0756_ & ~_0275_;
	assign _0758_ = _0757_ ^ _0276_;
	assign _0759_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0465_ : _0758_);
	assign _0760_ = (_1150_ ? _0759_ : _0755_);
	assign _0761_ = (_1102_ ? _0465_ : _0760_);
	assign _0762_ = _0761_ ^ _0741_;
	assign _0763_ = _0732_ ^ _0713_;
	assign _0764_ = _0762_ | ~_0763_;
	assign _0765_ = _0748_ & ~_0764_;
	assign _0766_ = _0765_ | _0747_;
	assign _0767_ = _0763_ ^ _0762_;
	assign _0768_ = _0748_ & ~_0767_;
	assign _0769_ = _0443_ ^ _0442_;
	assign _0770_ = _0440_ ^ _0390_;
	assign _0771_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0769_ : _0770_);
	assign _0772_ = _0474_ ^ _0334_;
	assign _0773_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0465_ : _0772_);
	assign _0774_ = (_1150_ ? _0773_ : _0771_);
	assign _0775_ = (_1102_ ? _0465_ : _0774_);
	assign _0776_ = _0775_ ^ _0741_;
	assign _0777_ = ~(_0730_ ^ _0721_);
	assign _0778_ = _0776_ | ~_0777_;
	assign _0779_ = ~(_0777_ ^ _0776_);
	assign _0780_ = _0729_ ^ _2122_;
	assign _0781_ = _0780_ ^ _0725_;
	assign _0782_ = _0781_ ^ _2122_;
	assign _0783_ = ~_0782_;
	assign _0784_ = ~_0465_;
	assign _0785_ = _0362_ & ~_0470_;
	assign _0786_ = _0359_ & ~_0785_;
	assign _0787_ = ~(_0786_ ^ _0352_);
	assign _0788_ = ~_0787_;
	assign _0789_ = _0414_ & ~_0438_;
	assign _0790_ = _0411_ & ~_0789_;
	assign _0791_ = ~(_0790_ ^ _0404_);
	assign _0792_ = ~_0791_;
	assign _0793_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0788_ : _0792_);
	assign _0794_ = _0476_ | _0251_;
	assign _0795_ = _0794_ & ~_0247_;
	assign _0796_ = ~(_0795_ ^ _0248_);
	assign _0797_ = ~(_0314_ & _0467_);
	assign _0798_ = _0797_ & ~_0329_;
	assign _0799_ = _0798_ ^ _0325_;
	assign _0800_ = ~_0799_;
	assign _0801_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0796_ : _0800_);
	assign _0802_ = (_1150_ ? _0801_ : _0793_);
	assign _0803_ = (_1102_ ? _0784_ : _0802_);
	assign _0804_ = (_0803_ ? _0741_ : _0783_);
	assign _0805_ = _0779_ & ~_0804_;
	assign _0806_ = _0778_ & ~_0805_;
	assign _0807_ = _0768_ & ~_0806_;
	assign _0808_ = _0807_ | _0766_;
	assign _0809_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0799_ : _0787_);
	assign _0810_ = _0795_ ^ _0248_;
	assign _0811_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0465_ : _0810_);
	assign _0812_ = (_1150_ ? _0811_ : _0809_);
	assign _0813_ = (_1102_ ? _0465_ : _0812_);
	assign _0814_ = _0813_ ^ _0741_;
	assign _0815_ = _0734_ ^ _0695_;
	assign _0816_ = _0815_ ^ _0814_;
	assign _0817_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0772_ : _0769_);
	assign _0818_ = (_1150_ ? _0465_ : _0817_);
	assign _0819_ = (_1102_ ? _0465_ : _0818_);
	assign _0820_ = ~(_0819_ ^ _0741_);
	assign _0821_ = ~(_0734_ | _0695_);
	assign _0822_ = _0821_ | ~_0687_;
	assign _0823_ = _0822_ ^ _0682_;
	assign _0824_ = ~(_0823_ ^ _0820_);
	assign _0825_ = _0824_ | _0816_;
	assign _0826_ = _0808_ & ~_0825_;
	assign _0827_ = _0815_ & ~_0814_;
	assign _0828_ = _0827_ & ~_0824_;
	assign _0829_ = _0823_ & _0820_;
	assign _0830_ = _0829_ | _0828_;
	assign _0831_ = _0830_ | _0826_;
	assign _0832_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0758_ : _0751_);
	assign _0833_ = (_1150_ ? _0465_ : _0832_);
	assign _0834_ = (_1102_ ? _0465_ : _0833_);
	assign _0835_ = _0834_ ^ _0741_;
	assign _0836_ = _0734_ | _0696_;
	assign _0837_ = _0836_ & ~_0690_;
	assign _0838_ = _0837_ ^ _0691_;
	assign _0839_ = _0838_ ^ _0835_;
	assign _0840_ = _0839_ ^ _0831_;
	assign _0841_ = ~_0840_;
	assign _0842_ = _0593_ | _0568_;
	assign _0843_ = _0842_ & ~_0562_;
	assign _0844_ = ~(_0843_ ^ _0563_);
	assign _0845_ = _0741_ ^ _2017_;
	assign _0846_ = ~(_0845_ & _0844_);
	assign _0847_ = _0593_ ^ _0568_;
	assign _0848_ = _0741_ ^ _0558_;
	assign _0849_ = _0848_ & _0847_;
	assign _0850_ = _0845_ ^ _0844_;
	assign _0851_ = ~(_0850_ & _0849_);
	assign _0852_ = ~(_0851_ & _0846_);
	assign _0853_ = _0848_ ^ _0847_;
	assign _0854_ = _0853_ & _0850_;
	assign _0855_ = _0580_ & ~_0591_;
	assign _0856_ = _0577_ & ~_0855_;
	assign _0857_ = _0856_ ^ _0575_;
	assign _0858_ = ~(_0857_ & _0845_);
	assign _0859_ = _0857_ ^ _0845_;
	assign _0860_ = ~(_0591_ ^ _0580_);
	assign _0861_ = ~(_0860_ & _0741_);
	assign _0862_ = _0859_ & ~_0861_;
	assign _0863_ = _0858_ & ~_0862_;
	assign _0864_ = _0860_ ^ _0741_;
	assign _0865_ = _0864_ & _0859_;
	assign _0866_ = ~(_0589_ ^ _0586_);
	assign _0867_ = ~(_0866_ & _0845_);
	assign _0868_ = ~(_0866_ ^ _0845_);
	assign _0869_ = _0588_ ^ _0502_;
	assign _0870_ = _0869_ ^ _0253_;
	assign _0871_ = (_0583_ ? _0741_ : _0870_);
	assign _0872_ = _0871_ & ~_0868_;
	assign _0873_ = _0867_ & ~_0872_;
	assign _0874_ = _0865_ & ~_0873_;
	assign _0875_ = _0863_ & ~_0874_;
	assign _0876_ = _0854_ & ~_0875_;
	assign _0877_ = _0876_ | _0852_;
	assign _0878_ = _0569_ & ~_0593_;
	assign _0879_ = _0565_ & ~_0878_;
	assign _0880_ = ~(_0879_ ^ _0553_);
	assign _0881_ = _0880_ ^ _0845_;
	assign _0882_ = ~_0881_;
	assign _0883_ = _0882_ ^ _0877_;
	assign _0884_ = ~_0883_;
	assign _0060_ = (io_in[10] ? _0884_ : _0841_);
	assign _0885_ = _0838_ & ~_0835_;
	assign _0886_ = _0831_ & ~_0839_;
	assign _0887_ = ~(_0886_ | _0885_);
	assign _0888_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0477_ : _0468_);
	assign _0889_ = (_1150_ ? _0465_ : _0888_);
	assign _0890_ = (_1102_ ? _0465_ : _0889_);
	assign _0891_ = ~(_0890_ ^ _0741_);
	assign _0892_ = ~(_0837_ | _0691_);
	assign _0893_ = _0675_ & ~_0892_;
	assign _0894_ = ~(_0893_ ^ _0670_);
	assign _0895_ = ~(_0894_ ^ _0891_);
	assign _0896_ = _0895_ ^ _0887_;
	assign _0897_ = _0880_ & _0845_;
	assign _0898_ = _0877_ & ~_0882_;
	assign _0899_ = ~(_0898_ | _0897_);
	assign _0900_ = _0553_ & ~_0879_;
	assign _0901_ = _0550_ & ~_0900_;
	assign _0902_ = _0901_ ^ _0548_;
	assign _0903_ = _0902_ ^ _0845_;
	assign _0904_ = _0903_ ^ _0899_;
	assign _0905_ = ~_0904_;
	assign _0061_ = (io_in[10] ? _0905_ : _0896_);
	assign _0906_ = _0895_ | _0839_;
	assign _0907_ = _0906_ | _0825_;
	assign _0908_ = _0808_ & ~_0907_;
	assign _0909_ = _0830_ & ~_0906_;
	assign _0910_ = _0894_ & _0891_;
	assign _0911_ = _0885_ & ~_0895_;
	assign _0912_ = _0911_ | _0910_;
	assign _0913_ = _0912_ | _0909_;
	assign _0914_ = _0913_ | _0908_;
	assign _0915_ = ~_0741_;
	assign _0916_ = (_1150_ ? _0784_ : _0801_);
	assign _0917_ = (_1102_ ? _0784_ : _0916_);
	assign _0918_ = _0917_ ^ _0915_;
	assign _0919_ = _0736_ ^ _0661_;
	assign _0920_ = _0919_ ^ _0918_;
	assign _0921_ = _0920_ ^ _0914_;
	assign _0922_ = ~_0921_;
	assign _0923_ = ~(_0903_ & _0881_);
	assign _0924_ = _0923_ | ~_0854_;
	assign _0925_ = ~(_0924_ | _0875_);
	assign _0926_ = _0902_ & _0845_;
	assign _0927_ = _0903_ & _0897_;
	assign _0928_ = _0927_ | _0926_;
	assign _0929_ = _0852_ & ~_0923_;
	assign _0930_ = _0929_ | _0928_;
	assign _0931_ = _0930_ | _0925_;
	assign _0932_ = _0595_ ^ _0538_;
	assign _0933_ = _0741_ ^ _1688_;
	assign _0934_ = _0933_ ^ _0932_;
	assign _0935_ = _0934_ ^ _0931_;
	assign _0062_ = (io_in[10] ? _0935_ : _0922_);
	assign _0937_ = _0919_ & ~_0918_;
	assign _0938_ = _0914_ & ~_0920_;
	assign _0939_ = ~(_0938_ | _0937_);
	assign _0940_ = (_1150_ ? _0465_ : _0773_);
	assign _0941_ = (_1102_ ? _0465_ : _0940_);
	assign _0942_ = ~(_0941_ ^ _0741_);
	assign _0943_ = ~(_0736_ | _0661_);
	assign _0944_ = _0943_ | ~_0654_;
	assign _0945_ = _0944_ ^ _0647_;
	assign _0947_ = _0945_ ^ _0942_;
	assign _0948_ = ~_0947_;
	assign _0949_ = _0948_ ^ _0939_;
	assign _0950_ = _0933_ & _0932_;
	assign _0951_ = _0934_ & _0931_;
	assign _0952_ = _0951_ | _0950_;
	assign _0953_ = _0595_ | _0538_;
	assign _0954_ = _0953_ & ~_0530_;
	assign _0955_ = ~(_0954_ ^ _0531_);
	assign _0956_ = _0955_ ^ _0845_;
	assign _0958_ = _0956_ ^ _0952_;
	assign _0063_ = (io_in[10] ? _0958_ : _0949_);
	assign _0959_ = _0948_ | _0920_;
	assign _0960_ = _0914_ & ~_0959_;
	assign _0961_ = _0945_ & _0942_;
	assign _0962_ = _0937_ & ~_0948_;
	assign _0963_ = _0962_ | _0961_;
	assign _0964_ = _0963_ | _0960_;
	assign _0965_ = (_1150_ ? _0465_ : _0759_);
	assign _0966_ = (_1102_ ? _0465_ : _0965_);
	assign _0967_ = ~(_0966_ ^ _0741_);
	assign _0968_ = ~(_0736_ | _0662_);
	assign _0969_ = _0656_ & ~_0968_;
	assign _0970_ = _0969_ ^ _0640_;
	assign _0971_ = ~(_0970_ ^ _0967_);
	assign _0972_ = ~(_0971_ ^ _0964_);
	assign _0973_ = _0955_ & _0845_;
	assign _0974_ = _0956_ & _0950_;
	assign _0975_ = _0974_ | _0973_;
	assign _0976_ = ~(_0956_ & _0934_);
	assign _0977_ = _0931_ & ~_0976_;
	assign _0978_ = _0977_ | _0975_;
	assign _0979_ = ~(_0595_ | _0539_);
	assign _0980_ = _0533_ & ~_0979_;
	assign _0981_ = _0980_ ^ _0522_;
	assign _0982_ = _0981_ ^ _0845_;
	assign _0983_ = _0982_ ^ _0978_;
	assign _0053_ = (io_in[10] ? _0983_ : _0972_);
	assign _0984_ = _0970_ & _0967_;
	assign _0985_ = _0964_ & ~_0971_;
	assign _0986_ = _0985_ | _0984_;
	assign _0987_ = (_1150_ ? _0465_ : _0478_);
	assign _0988_ = (_1102_ ? _0465_ : _0987_);
	assign _0989_ = ~(_0988_ ^ _0741_);
	assign _0990_ = ~(_0969_ | _0640_);
	assign _0991_ = _0637_ & ~_0990_;
	assign _0992_ = ~(_0991_ ^ _0632_);
	assign _0993_ = _0992_ ^ _0989_;
	assign _0994_ = _0993_ ^ _0986_;
	assign _0995_ = _0981_ & _0845_;
	assign _0996_ = _0982_ & _0978_;
	assign _0997_ = _0996_ | _0995_;
	assign _0998_ = _0980_ | _0522_;
	assign _0999_ = _0998_ & ~_0518_;
	assign _1000_ = ~(_0999_ ^ _0519_);
	assign _1001_ = _1000_ ^ _0845_;
	assign _1002_ = _1001_ ^ _0997_;
	assign _0054_ = (io_in[10] ? _1002_ : _0994_);
	assign _1003_ = _0971_ | ~_0993_;
	assign _1004_ = _1003_ | _0959_;
	assign _1005_ = _0914_ & ~_1004_;
	assign _1006_ = _0963_ & ~_1003_;
	assign _1007_ = _0992_ & _0989_;
	assign _1008_ = _0993_ & _0984_;
	assign _1009_ = _1008_ | _1007_;
	assign _1010_ = _1009_ | _1006_;
	assign _1011_ = _1010_ | _1005_;
	assign _1012_ = (_1150_ ? _0465_ : _0811_);
	assign _1013_ = (_1102_ ? _0465_ : _1012_);
	assign _1014_ = ~(_1013_ ^ _0741_);
	assign _1015_ = _0663_ & ~_0736_;
	assign _1016_ = _0658_ & ~_1015_;
	assign _1017_ = _1016_ ^ _0624_;
	assign _1018_ = ~(_1017_ ^ _1014_);
	assign _1019_ = ~(_1018_ ^ _1011_);
	assign _1020_ = ~(_1001_ & _0982_);
	assign _1021_ = _1020_ | _0976_;
	assign _1022_ = _0931_ & ~_1021_;
	assign _1023_ = _0975_ & ~_1020_;
	assign _1024_ = _1000_ & _0845_;
	assign _1025_ = _1001_ & _0995_;
	assign _1026_ = _1025_ | _1024_;
	assign _1027_ = _1026_ | _1023_;
	assign _1028_ = _1027_ | _1022_;
	assign _1029_ = _0540_ & ~_0595_;
	assign _1030_ = _0535_ & ~_1029_;
	assign _1031_ = _1030_ ^ _0508_;
	assign _1032_ = _1031_ ^ _0741_;
	assign _1033_ = _1032_ ^ _1028_;
	assign _0055_ = (io_in[10] ? _1033_ : _1019_);
	assign _1034_ = _1017_ & _1014_;
	assign _1035_ = _1011_ & ~_1018_;
	assign _1036_ = _1035_ | _1034_;
	assign _1037_ = ~(_0741_ ^ _0465_);
	assign _1038_ = ~(_1016_ | _0624_);
	assign _1039_ = _0619_ & ~_1038_;
	assign _1040_ = ~(_1039_ ^ _0614_);
	assign _1041_ = _1040_ ^ _1037_;
	assign _1042_ = _1041_ ^ _1036_;
	assign _1043_ = _1031_ & _0741_;
	assign _1044_ = _1032_ & _1028_;
	assign _1045_ = _1044_ | _1043_;
	assign _1046_ = ~(_1030_ | _0508_);
	assign _1047_ = _0503_ & ~_1046_;
	assign _1048_ = ~(_1047_ ^ _0500_);
	assign _1049_ = _1048_ ^ _0741_;
	assign _1050_ = _1049_ ^ _1045_;
	assign _0056_ = (io_in[10] ? _1050_ : _1042_);
	assign _1051_ = _1040_ & _1037_;
	assign _1052_ = ~_1041_;
	assign _1053_ = _1034_ & ~_1052_;
	assign _1054_ = _1053_ | _1051_;
	assign _1055_ = _1052_ | _1018_;
	assign _1056_ = _1011_ & ~_1055_;
	assign _1057_ = _1056_ | _1054_;
	assign _1058_ = _0625_ & ~_1016_;
	assign _1059_ = _0621_ & ~_1058_;
	assign _1060_ = ~(_1059_ ^ _0607_);
	assign _1061_ = _1060_ ^ _1037_;
	assign _1062_ = _1061_ ^ _1057_;
	assign _1063_ = _1048_ & _0741_;
	assign _1064_ = _1049_ & _1043_;
	assign _1065_ = _1064_ | _1063_;
	assign _1066_ = ~(_1049_ & _1032_);
	assign _1067_ = _1028_ & ~_1066_;
	assign _1068_ = _1067_ | _1065_;
	assign _1069_ = _0509_ & ~_1030_;
	assign _1070_ = _0505_ & ~_1069_;
	assign _1071_ = ~(_1070_ ^ _0494_);
	assign _1072_ = _1071_ ^ _0741_;
	assign _1073_ = _1072_ ^ _1068_;
	assign _0057_ = (io_in[10] ? _1073_ : _1062_);
	assign _1074_ = _1060_ & _1037_;
	assign _1075_ = _1061_ & _1057_;
	assign _1076_ = _1075_ | _1074_;
	assign _1077_ = _0607_ & ~_1059_;
	assign _1078_ = _0604_ & ~_1077_;
	assign _1079_ = _1078_ ^ _0603_;
	assign _1080_ = _1079_ ^ _1037_;
	assign _1081_ = _1080_ ^ _1076_;
	assign _1082_ = _1071_ & _0741_;
	assign _1083_ = _1072_ & _1068_;
	assign _1084_ = _1083_ | _1082_;
	assign _1085_ = _0494_ & ~_1070_;
	assign _1086_ = _0491_ & ~_1085_;
	assign _1087_ = _1086_ ^ _0489_;
	assign _1088_ = _1087_ ^ _0741_;
	assign _1089_ = _1088_ ^ _1084_;
	assign _0058_ = (io_in[10] ? _1089_ : _1081_);
	assign _1090_ = _1079_ & _1037_;
	assign _1092_ = _1080_ & _1074_;
	assign _1093_ = ~(_1092_ | _1090_);
	assign _1094_ = ~(_1080_ & _1061_);
	assign _1095_ = _1054_ & ~_1094_;
	assign _1096_ = _1093_ & ~_1095_;
	assign _1097_ = _1094_ | _1055_;
	assign _1098_ = _1010_ & ~_1097_;
	assign _1099_ = _1096_ & ~_1098_;
	assign _1100_ = _1097_ | _1004_;
	assign _1101_ = _0914_ & ~_1100_;
	assign _1103_ = _1099_ & ~_1101_;
	assign _1104_ = _1037_ ^ _0740_;
	assign _1105_ = ~(_1104_ ^ _1103_);
	assign _1106_ = _1087_ & _0741_;
	assign _1107_ = _1088_ & _1082_;
	assign _1108_ = _1107_ | _1106_;
	assign _1109_ = ~(_1088_ & _1072_);
	assign _1110_ = _1065_ & ~_1109_;
	assign _1111_ = _1110_ | _1108_;
	assign _1112_ = _1109_ | _1066_;
	assign _1114_ = _1027_ & ~_1112_;
	assign _1115_ = _1114_ | _1111_;
	assign _1116_ = _1112_ | _1021_;
	assign _1117_ = _0931_ & ~_1116_;
	assign _1118_ = _1117_ | _1115_;
	assign _1119_ = _0741_ ^ _0599_;
	assign _1120_ = _1119_ ^ _1118_;
	assign _0059_ = (io_in[10] ? _1120_ : _1105_);
	assign _1121_ = _0946_ & ~_0957_;
	assign _1122_ = ~_1121_;
	assign _1124_ = ~(_0741_ ^ _0583_);
	assign _1125_ = _1124_ ^ _0870_;
	assign _1126_ = _1125_ ^ _0915_;
	assign _0036_ = _1122_ & ~_1126_;
	assign _1127_ = _0871_ ^ _0868_;
	assign _0044_ = _1122_ & ~_1127_;
	assign _1128_ = _0873_ ^ _0864_;
	assign _0045_ = _1122_ & ~_1128_;
	assign _1129_ = _0864_ & ~_0873_;
	assign _1130_ = _0861_ & ~_1129_;
	assign _1132_ = _1130_ ^ _0859_;
	assign _0046_ = _1122_ & ~_1132_;
	assign _1133_ = _0875_ ^ _0853_;
	assign _0047_ = _1122_ & ~_1133_;
	assign _1134_ = _0875_ | ~_0853_;
	assign _1135_ = _1134_ & ~_0849_;
	assign _1136_ = _1135_ ^ _0850_;
	assign _0048_ = _1122_ & ~_1136_;
	assign _0049_ = _1122_ & ~_0883_;
	assign _0050_ = _1122_ & ~_0904_;
	assign _1138_ = io_in[0] & ~io_in[10];
	assign _0051_ = (_1121_ ? _1138_ : _0935_);
	assign _1139_ = io_in[1] & ~io_in[10];
	assign _0052_ = (_1121_ ? _1139_ : _0958_);
	assign _1140_ = io_in[2] & ~io_in[10];
	assign _0037_ = (_1121_ ? _1140_ : _0983_);
	assign _1141_ = io_in[3] & ~io_in[10];
	assign _0038_ = (_1121_ ? _1141_ : _1002_);
	assign _1142_ = io_in[4] & ~io_in[10];
	assign _0039_ = (_1121_ ? _1142_ : _1033_);
	assign _1144_ = io_in[5] & ~io_in[10];
	assign _0040_ = (_1121_ ? _1144_ : _1050_);
	assign _1145_ = io_in[6] & ~io_in[10];
	assign _0041_ = (_1121_ ? _1145_ : _1073_);
	assign _1146_ = io_in[7] & ~io_in[10];
	assign _0042_ = (_1121_ ? _1146_ : _1089_);
	assign _1147_ = io_in[8] & ~io_in[10];
	assign _0043_ = (_1121_ ? _1147_ : _1120_);
	assign _1148_ = _0803_ ^ _0915_;
	assign _1149_ = _1148_ ^ _0783_;
	assign _1151_ = _1149_ ^ _0741_;
	assign _0002_ = _1122_ & ~_1151_;
	assign _1152_ = _0804_ ^ _0779_;
	assign _0010_ = _1122_ & ~_1152_;
	assign _1153_ = ~_0767_;
	assign _1154_ = _0806_ ^ _1153_;
	assign _0011_ = _1122_ & ~_1154_;
	assign _1155_ = _1153_ & ~_0806_;
	assign _1156_ = _0764_ & ~_1155_;
	assign _1157_ = _1156_ ^ _0748_;
	assign _0012_ = _1122_ & ~_1157_;
	assign _1159_ = _0816_ ^ _0808_;
	assign _0013_ = _1122_ & ~_1159_;
	assign _1160_ = _0808_ & ~_0816_;
	assign _1161_ = _1160_ | _0827_;
	assign _1162_ = _1161_ ^ _0824_;
	assign _0014_ = _1122_ & ~_1162_;
	assign _0015_ = _1122_ & ~_0840_;
	assign _0016_ = _0896_ & ~_1121_;
	assign _0017_ = _1122_ & ~_0921_;
	assign _0018_ = _0949_ & ~_1121_;
	assign _1164_ = io_in[0] & io_in[10];
	assign _0003_ = (_1121_ ? _1164_ : _0972_);
	assign _1165_ = io_in[1] & io_in[10];
	assign _0004_ = (_1121_ ? _1165_ : _0994_);
	assign _1166_ = io_in[2] & io_in[10];
	assign _0005_ = (_1121_ ? _1166_ : _1019_);
	assign _1167_ = io_in[3] & io_in[10];
	assign _0006_ = (_1121_ ? _1167_ : _1042_);
	assign _1168_ = io_in[4] & io_in[10];
	assign _0007_ = (_1121_ ? _1168_ : _1062_);
	assign _0008_ = _1081_ & ~_1121_;
	assign _0009_ = _1105_ & ~_1121_;
	assign _1170_ = ~_0740_;
	assign _1171_ = ~_0894_;
	assign _1172_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1171_ : _0746_);
	assign _1173_ = ~_0992_;
	assign _1174_ = ~(_1078_ ^ _0603_);
	assign _1175_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1174_ : _1173_);
	assign _1176_ = (_1150_ ? _1175_ : _1172_);
	assign _1178_ = (_1102_ ? _1170_ : _1176_);
	assign _1179_ = _1178_ ^ _0915_;
	assign _1180_ = _0435_ ^ _0253_;
	assign _1181_ = _1180_ ^ _0430_;
	assign _1182_ = _1181_ ^ _0253_;
	assign _1183_ = _1182_ ^ _1179_;
	assign _1184_ = _1183_ ^ _0915_;
	assign _0019_ = _1122_ & ~_1184_;
	assign _1185_ = (_1178_ ? _0741_ : _1182_);
	assign _1186_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0919_ : _0815_);
	assign _1188_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0740_ : _1017_);
	assign _1189_ = (_1150_ ? _1188_ : _1186_);
	assign _1190_ = (_1102_ ? _0740_ : _1189_);
	assign _1191_ = _1190_ ^ _0741_;
	assign _1192_ = ~(_0436_ ^ _0426_);
	assign _1193_ = ~_1192_;
	assign _1194_ = _1193_ ^ _1191_;
	assign _1195_ = ~(_1194_ ^ _1185_);
	assign _0027_ = (_1121_ ? _1091_ : _1195_);
	assign _1196_ = _1185_ & ~_1194_;
	assign _1198_ = _1191_ & ~_1193_;
	assign _1199_ = _1198_ | _1196_;
	assign _1200_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0945_ : _0823_);
	assign _1201_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0740_ : _1040_);
	assign _1202_ = (_1150_ ? _1201_ : _1200_);
	assign _1203_ = (_1102_ ? _0740_ : _1202_);
	assign _1204_ = _1203_ ^ _0741_;
	assign _1205_ = _0438_ ^ _0415_;
	assign _1206_ = ~(_1205_ ^ _1204_);
	assign _1207_ = _1206_ ^ _1199_;
	assign _0028_ = _1122_ & ~_1207_;
	assign _1209_ = _1205_ & _1204_;
	assign _1210_ = _1199_ & ~_1206_;
	assign _1211_ = ~(_1210_ | _1209_);
	assign _1212_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0970_ : _0838_);
	assign _1213_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0740_ : _1060_);
	assign _1214_ = (_1150_ ? _1213_ : _1212_);
	assign _1215_ = (_1102_ ? _0740_ : _1214_);
	assign _1216_ = _1215_ ^ _0741_;
	assign _1217_ = ~(_1216_ ^ _0791_);
	assign _1219_ = _1217_ ^ _1211_;
	assign _0029_ = (_1121_ ? _1091_ : _1219_);
	assign _1220_ = _1217_ | _1206_;
	assign _1221_ = _1199_ & ~_1220_;
	assign _1222_ = _1216_ & _0791_;
	assign _1223_ = _1209_ & ~_1217_;
	assign _1224_ = _1223_ | _1222_;
	assign _1225_ = _1224_ | _1221_;
	assign _1226_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0992_ : _0894_);
	assign _1227_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _0740_ : _1079_);
	assign _1229_ = (_1150_ ? _1227_ : _1226_);
	assign _1230_ = (_1102_ ? _0740_ : _1229_);
	assign _1231_ = ~(_1230_ ^ _0741_);
	assign _1232_ = _1231_ ^ _0770_;
	assign _1233_ = ~(_1232_ ^ _1225_);
	assign _0030_ = (_1121_ ? _1091_ : _1233_);
	assign _1234_ = _0770_ & ~_1231_;
	assign _1235_ = _1232_ | ~_1225_;
	assign _1236_ = _1235_ & ~_1234_;
	assign _1237_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1017_ : _0919_);
	assign _1239_ = (_1150_ ? _0740_ : _1237_);
	assign _1240_ = (_1102_ ? _0740_ : _1239_);
	assign _1241_ = _1240_ ^ _0741_;
	assign _1242_ = ~(_1241_ ^ _0754_);
	assign _1243_ = _1242_ ^ _1236_;
	assign _0031_ = (_1121_ ? _1091_ : _1243_);
	assign _1244_ = _1242_ | _1232_;
	assign _1245_ = _1225_ & ~_1244_;
	assign _1246_ = _1234_ & ~_1242_;
	assign _1247_ = _1241_ & _0754_;
	assign _1249_ = _1247_ | _1246_;
	assign _1250_ = _1249_ | _1245_;
	assign _1251_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1040_ : _0945_);
	assign _1252_ = (_1150_ ? _0740_ : _1251_);
	assign _1253_ = (_1102_ ? _0740_ : _1252_);
	assign _1254_ = _1253_ ^ _0741_;
	assign _1255_ = ~(_1254_ ^ _0471_);
	assign \mchip.cordic_module.next_x [6] = ~(_1255_ ^ _1250_);
	assign _0032_ = \mchip.cordic_module.next_x [6] & ~_1121_;
	assign _1256_ = _1254_ & _0471_;
	assign _1258_ = _1250_ & ~_1255_;
	assign _1259_ = ~(_1258_ | _1256_);
	assign _1260_ = (\mchip.cordic_module.fstage_0.stage_0.step_ctr [2] ? _1060_ : _0970_);
	assign _1261_ = (_1150_ ? _0740_ : _1260_);
	assign _1262_ = (_1102_ ? _0740_ : _1261_);
	assign _1263_ = _1262_ ^ _0741_;
	assign _1264_ = ~(_1263_ ^ _0787_);
	assign \mchip.cordic_module.next_x [7] = _1264_ ^ _1259_;
	assign _0033_ = (_1121_ ? _1091_ : \mchip.cordic_module.next_x [7]);
	assign _1265_ = _1264_ | _1255_;
	assign _1267_ = _1265_ | _1244_;
	assign _1268_ = _1225_ & ~_1267_;
	assign _1269_ = _1249_ & ~_1265_;
	assign _1270_ = _1263_ & _0787_;
	assign _1271_ = _1256_ & ~_1264_;
	assign _1272_ = _1271_ | _1270_;
	assign _1273_ = _1272_ | _1269_;
	assign _1274_ = _1273_ | _1268_;
	assign _1275_ = (_1150_ ? _1170_ : _1175_);
	assign _1276_ = (_1102_ ? _1170_ : _1275_);
	assign _1278_ = _1276_ ^ _0741_;
	assign _1279_ = _1278_ ^ _0769_;
	assign \mchip.cordic_module.next_x [8] = ~(_1279_ ^ _1274_);
	assign _0034_ = (_1121_ ? _1091_ : \mchip.cordic_module.next_x [8]);
	assign _1280_ = _0769_ & ~_1278_;
	assign _1281_ = _1274_ & ~_1279_;
	assign _1282_ = ~(_1281_ | _1280_);
	assign _1283_ = (_1150_ ? _0740_ : _1188_);
	assign _1284_ = (_1102_ ? _0740_ : _1283_);
	assign _1285_ = _1284_ ^ _0741_;
	assign _1287_ = _1285_ ^ _0751_;
	assign _1288_ = _1287_ ^ _1282_;
	assign \mchip.cordic_module.next_x [9] = ~_1288_;
	assign _0035_ = _1122_ & ~_1288_;
	assign _1289_ = ~_1287_;
	assign _1290_ = _1289_ | _1279_;
	assign _1291_ = _1274_ & ~_1290_;
	assign _1292_ = _1285_ & _0751_;
	assign _1293_ = _1280_ & ~_1289_;
	assign _1294_ = _1293_ | _1292_;
	assign _1296_ = _1294_ | _1291_;
	assign _1297_ = (_1150_ ? _0740_ : _1201_);
	assign _1298_ = (_1102_ ? _0740_ : _1297_);
	assign _1299_ = _1298_ ^ _0741_;
	assign _1300_ = _1299_ ^ _0468_;
	assign \mchip.cordic_module.next_x [10] = _1300_ ^ _1296_;
	assign _1301_ = io_in[5] | ~io_in[10];
	assign _0020_ = (_1121_ ? _1301_ : \mchip.cordic_module.next_x [10]);
	assign _1302_ = _1299_ & _0468_;
	assign _1303_ = _1300_ & _1296_;
	assign _1305_ = _1303_ | _1302_;
	assign _1306_ = (_1150_ ? _0740_ : _1213_);
	assign _1307_ = (_1102_ ? _0740_ : _1306_);
	assign _1308_ = _1307_ ^ _0741_;
	assign _1309_ = _1308_ ^ _0799_;
	assign \mchip.cordic_module.next_x [11] = _1309_ ^ _1305_;
	assign _1310_ = io_in[6] | ~io_in[10];
	assign _0021_ = (_1121_ ? _1310_ : \mchip.cordic_module.next_x [11]);
	assign _1311_ = ~(_1309_ & _1300_);
	assign _1312_ = _1311_ | _1290_;
	assign _1314_ = _1274_ & ~_1312_;
	assign _1315_ = _1294_ & ~_1311_;
	assign _1316_ = _1308_ & _0799_;
	assign _1317_ = _1309_ & _1302_;
	assign _1318_ = _1317_ | _1316_;
	assign _1319_ = _1318_ | _1315_;
	assign _1320_ = _1319_ | _1314_;
	assign _1321_ = (_1150_ ? _0740_ : _1227_);
	assign _1322_ = (_1102_ ? _0740_ : _1321_);
	assign _1323_ = _1322_ ^ _0741_;
	assign _1325_ = _1323_ ^ _0772_;
	assign \mchip.cordic_module.next_x [12] = _1325_ ^ _1320_;
	assign _1326_ = io_in[7] & io_in[10];
	assign _0022_ = (_1121_ ? _1326_ : \mchip.cordic_module.next_x [12]);
	assign _1327_ = _1323_ & _0772_;
	assign _1328_ = _1325_ & _1320_;
	assign _1329_ = _1328_ | _1327_;
	assign _1330_ = _0741_ ^ _0740_;
	assign _1331_ = _1330_ ^ _0758_;
	assign \mchip.cordic_module.next_x [13] = _1331_ ^ _1329_;
	assign _1333_ = io_in[8] & io_in[10];
	assign _0023_ = (_1121_ ? _1333_ : \mchip.cordic_module.next_x [13]);
	assign _1334_ = _1330_ & _0758_;
	assign _1335_ = _1331_ & _1327_;
	assign _1336_ = _1335_ | _1334_;
	assign _1337_ = ~(_1331_ & _1325_);
	assign _1338_ = _1320_ & ~_1337_;
	assign _1339_ = _1338_ | _1336_;
	assign _1340_ = _1330_ ^ _0477_;
	assign \mchip.cordic_module.next_x [14] = _1340_ ^ _1339_;
	assign _1342_ = io_in[9] | ~io_in[10];
	assign _0024_ = (_1121_ ? _1342_ : \mchip.cordic_module.next_x [14]);
	assign _1343_ = _1330_ & _0477_;
	assign _1344_ = _1340_ & _1339_;
	assign _1345_ = _1344_ | _1343_;
	assign _1346_ = _1330_ ^ _0810_;
	assign \mchip.cordic_module.next_x [15] = _1346_ ^ _1345_;
	assign _0025_ = \mchip.cordic_module.next_x [15] & ~_1121_;
	assign _1347_ = _1330_ & _0810_;
	assign _1348_ = _1346_ & _1343_;
	assign _1350_ = ~(_1348_ | _1347_);
	assign _1351_ = ~(_1346_ & _1340_);
	assign _1352_ = _1336_ & ~_1351_;
	assign _1353_ = _1350_ & ~_1352_;
	assign _1354_ = _1351_ | _1337_;
	assign _1355_ = _1319_ & ~_1354_;
	assign _1356_ = _1353_ & ~_1355_;
	assign _1357_ = _1354_ | _1312_;
	assign _1358_ = _1274_ & ~_1357_;
	assign _1359_ = _1356_ & ~_1358_;
	assign _1361_ = _1330_ ^ _0465_;
	assign _1362_ = _1361_ ^ _1359_;
	assign \mchip.cordic_module.next_x [16] = ~_1362_;
	assign _0026_ = _1122_ & ~_1362_;
	assign _2134_[1] = ~(_1684_ & _1659_);
	assign _2134_[2] = _1686_ ^ _0957_;
	assign \mchip.cordic_module.done  = _0098_ & ~io_in[13];
	always @(posedge io_in[12])
		if (io_in[13])
			_0064_ <= 1'h0;
		else if (_0001_)
			_0064_ <= _0036_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0065_ <= 1'h0;
		else if (_0001_)
			_0065_ <= _0044_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0066_ <= 1'h0;
		else if (_0001_)
			_0066_ <= _0045_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0067_ <= 1'h0;
		else if (_0001_)
			_0067_ <= _0046_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0068_ <= 1'h0;
		else if (_0001_)
			_0068_ <= _0047_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0069_ <= 1'h0;
		else if (_0001_)
			_0069_ <= _0048_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0070_ <= 1'h0;
		else if (_0001_)
			_0070_ <= _0049_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0071_ <= 1'h0;
		else if (_0001_)
			_0071_ <= _0050_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0072_ <= 1'h0;
		else if (_0001_)
			_0072_ <= _0051_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0073_ <= 1'h0;
		else if (_0001_)
			_0073_ <= _0052_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0074_ <= 1'h0;
		else if (_0001_)
			_0074_ <= _0037_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0075_ <= 1'h0;
		else if (_0001_)
			_0075_ <= _0038_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0076_ <= 1'h0;
		else if (_0001_)
			_0076_ <= _0039_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0077_ <= 1'h0;
		else if (_0001_)
			_0077_ <= _0040_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0078_ <= 1'h0;
		else if (_0001_)
			_0078_ <= _0041_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0079_ <= 1'h0;
		else if (_0001_)
			_0079_ <= _0042_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0080_ <= 1'h0;
		else if (_0001_)
			_0080_ <= _0043_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0081_ <= 1'h0;
		else if (_0001_)
			_0081_ <= _0002_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0082_ <= 1'h0;
		else if (_0001_)
			_0082_ <= _0010_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0083_ <= 1'h0;
		else if (_0001_)
			_0083_ <= _0011_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0084_ <= 1'h0;
		else if (_0001_)
			_0084_ <= _0012_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0085_ <= 1'h0;
		else if (_0001_)
			_0085_ <= _0013_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0086_ <= 1'h0;
		else if (_0001_)
			_0086_ <= _0014_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0087_ <= 1'h0;
		else if (_0001_)
			_0087_ <= _0015_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0088_ <= 1'h0;
		else if (_0001_)
			_0088_ <= _0016_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0089_ <= 1'h0;
		else if (_0001_)
			_0089_ <= _0017_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0090_ <= 1'h0;
		else if (_0001_)
			_0090_ <= _0018_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0091_ <= 1'h0;
		else if (_0001_)
			_0091_ <= _0003_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0092_ <= 1'h0;
		else if (_0001_)
			_0092_ <= _0004_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0093_ <= 1'h0;
		else if (_0001_)
			_0093_ <= _0005_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0094_ <= 1'h0;
		else if (_0001_)
			_0094_ <= _0006_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0095_ <= 1'h0;
		else if (_0001_)
			_0095_ <= _0007_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0096_ <= 1'h0;
		else if (_0001_)
			_0096_ <= _0008_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0097_ <= 1'h0;
		else if (_0001_)
			_0097_ <= _0009_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0098_ <= 1'h0;
		else if (!_0001_)
			_0098_ <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			_0099_ <= 1'h0;
		else if (!\mchip.cordic_module.done )
			_0099_ <= \mchip.cordic_module.fstage_0.stage_0.step_ctr [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0100_ <= 1'h0;
		else if (!\mchip.cordic_module.done )
			_0100_ <= _2134_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0101_ <= 1'h0;
		else if (!\mchip.cordic_module.done )
			_0101_ <= _2134_[2];
	reg \mchip.cordic_module.out1_reg[6] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[6]  <= _0060_;
	assign \mchip.cordic_module.out1 [6] = \mchip.cordic_module.out1_reg[6] ;
	reg \mchip.cordic_module.out1_reg[7] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[7]  <= _0061_;
	assign \mchip.cordic_module.out1 [7] = \mchip.cordic_module.out1_reg[7] ;
	reg \mchip.cordic_module.out1_reg[8] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[8]  <= _0062_;
	assign \mchip.cordic_module.out1 [8] = \mchip.cordic_module.out1_reg[8] ;
	reg \mchip.cordic_module.out1_reg[9] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[9]  <= _0063_;
	assign \mchip.cordic_module.out1 [9] = \mchip.cordic_module.out1_reg[9] ;
	reg \mchip.cordic_module.out1_reg[10] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[10]  <= _0053_;
	assign \mchip.cordic_module.out1 [10] = \mchip.cordic_module.out1_reg[10] ;
	reg \mchip.cordic_module.out1_reg[11] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[11]  <= _0054_;
	assign \mchip.cordic_module.out1 [11] = \mchip.cordic_module.out1_reg[11] ;
	reg \mchip.cordic_module.out1_reg[12] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[12]  <= _0055_;
	assign \mchip.cordic_module.out1 [12] = \mchip.cordic_module.out1_reg[12] ;
	reg \mchip.cordic_module.out1_reg[13] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[13]  <= _0056_;
	assign \mchip.cordic_module.out1 [13] = \mchip.cordic_module.out1_reg[13] ;
	reg \mchip.cordic_module.out1_reg[14] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[14]  <= _0057_;
	assign \mchip.cordic_module.out1 [14] = \mchip.cordic_module.out1_reg[14] ;
	reg \mchip.cordic_module.out1_reg[15] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[15]  <= _0058_;
	assign \mchip.cordic_module.out1 [15] = \mchip.cordic_module.out1_reg[15] ;
	reg \mchip.cordic_module.out1_reg[16] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out1_reg[16]  <= _0059_;
	assign \mchip.cordic_module.out1 [16] = \mchip.cordic_module.out1_reg[16] ;
	reg \mchip.cordic_module.out2_reg[6] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[6]  <= \mchip.cordic_module.next_x [6];
	assign \mchip.cordic_module.out2 [6] = \mchip.cordic_module.out2_reg[6] ;
	reg \mchip.cordic_module.out2_reg[7] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[7]  <= \mchip.cordic_module.next_x [7];
	assign \mchip.cordic_module.out2 [7] = \mchip.cordic_module.out2_reg[7] ;
	reg \mchip.cordic_module.out2_reg[8] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[8]  <= \mchip.cordic_module.next_x [8];
	assign \mchip.cordic_module.out2 [8] = \mchip.cordic_module.out2_reg[8] ;
	reg \mchip.cordic_module.out2_reg[9] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[9]  <= \mchip.cordic_module.next_x [9];
	assign \mchip.cordic_module.out2 [9] = \mchip.cordic_module.out2_reg[9] ;
	reg \mchip.cordic_module.out2_reg[10] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[10]  <= \mchip.cordic_module.next_x [10];
	assign \mchip.cordic_module.out2 [10] = \mchip.cordic_module.out2_reg[10] ;
	reg \mchip.cordic_module.out2_reg[11] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[11]  <= \mchip.cordic_module.next_x [11];
	assign \mchip.cordic_module.out2 [11] = \mchip.cordic_module.out2_reg[11] ;
	reg \mchip.cordic_module.out2_reg[12] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[12]  <= \mchip.cordic_module.next_x [12];
	assign \mchip.cordic_module.out2 [12] = \mchip.cordic_module.out2_reg[12] ;
	reg \mchip.cordic_module.out2_reg[13] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[13]  <= \mchip.cordic_module.next_x [13];
	assign \mchip.cordic_module.out2 [13] = \mchip.cordic_module.out2_reg[13] ;
	reg \mchip.cordic_module.out2_reg[14] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[14]  <= \mchip.cordic_module.next_x [14];
	assign \mchip.cordic_module.out2 [14] = \mchip.cordic_module.out2_reg[14] ;
	reg \mchip.cordic_module.out2_reg[15] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[15]  <= \mchip.cordic_module.next_x [15];
	assign \mchip.cordic_module.out2 [15] = \mchip.cordic_module.out2_reg[15] ;
	reg \mchip.cordic_module.out2_reg[16] ;
	always @(posedge io_in[12])
		if (_0000_)
			\mchip.cordic_module.out2_reg[16]  <= \mchip.cordic_module.next_x [16];
	assign \mchip.cordic_module.out2 [16] = \mchip.cordic_module.out2_reg[16] ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0102_ <= 1'h0;
		else if (_0001_)
			_0102_ <= _0019_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0103_ <= 1'h0;
		else if (_0001_)
			_0103_ <= _0027_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0104_ <= 1'h0;
		else if (_0001_)
			_0104_ <= _0028_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0105_ <= 1'h0;
		else if (_0001_)
			_0105_ <= _0029_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0106_ <= 1'h0;
		else if (_0001_)
			_0106_ <= _0030_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0107_ <= 1'h0;
		else if (_0001_)
			_0107_ <= _0031_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0108_ <= 1'h0;
		else if (_0001_)
			_0108_ <= _0032_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0109_ <= 1'h0;
		else if (_0001_)
			_0109_ <= _0033_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0110_ <= 1'h0;
		else if (_0001_)
			_0110_ <= _0034_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0111_ <= 1'h0;
		else if (_0001_)
			_0111_ <= _0035_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0112_ <= 1'h0;
		else if (_0001_)
			_0112_ <= _0020_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0113_ <= 1'h0;
		else if (_0001_)
			_0113_ <= _0021_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0114_ <= 1'h0;
		else if (_0001_)
			_0114_ <= _0022_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0115_ <= 1'h0;
		else if (_0001_)
			_0115_ <= _0023_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0116_ <= 1'h0;
		else if (_0001_)
			_0116_ <= _0024_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0117_ <= 1'h0;
		else if (_0001_)
			_0117_ <= _0025_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0118_ <= 1'h0;
		else if (_0001_)
			_0118_ <= _0026_;
	assign _2134_[0] = \mchip.cordic_module.fstage_0.stage_0.step_ctr [2];
	assign io_out[13:11] = {2'h0, \mchip.cordic_module.done };
	assign \mchip.clock  = io_in[12];
	assign \mchip.cordic_module.clk  = io_in[12];
	assign \mchip.cordic_module.fstage_0.clk  = io_in[12];
	assign \mchip.cordic_module.fstage_0.mode  = io_in[10];
	assign \mchip.cordic_module.fstage_0.out_x  = {\mchip.cordic_module.next_x [16:6], 6'h00};
	assign \mchip.cordic_module.fstage_0.reset  = io_in[13];
	assign \mchip.cordic_module.fstage_0.stage_0.clk  = io_in[12];
	assign \mchip.cordic_module.fstage_0.stage_0.mode  = io_in[10];
	assign \mchip.cordic_module.fstage_0.stage_0.reset  = io_in[13];
	assign {\mchip.cordic_module.fstage_0.stage_0.step_ctr [4:3], \mchip.cordic_module.fstage_0.stage_0.step_ctr [1:0]} = 4'h0;
	assign \mchip.cordic_module.fstage_0.stage_0.subx.in_b [15:0] = 16'h0000;
	assign \mchip.cordic_module.fstage_0.stage_0.suby.in_b [15:0] = 16'h0000;
	assign \mchip.cordic_module.fstage_0.stage_0.subz.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_0.subz.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_0.subz.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_0.x_coeff [15:0] = 16'h0000;
	assign \mchip.cordic_module.fstage_0.stage_0.y_coeff [15:0] = 16'h0000;
	assign \mchip.cordic_module.fstage_0.stage_0.z_coeff  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_1.clk  = io_in[12];
	assign \mchip.cordic_module.fstage_0.stage_1.mode  = io_in[10];
	assign \mchip.cordic_module.fstage_0.stage_1.reset  = io_in[13];
	assign \mchip.cordic_module.fstage_0.stage_1.step_ctr  = {2'h0, \mchip.cordic_module.fstage_0.stage_0.step_ctr [2], 2'h1};
	assign \mchip.cordic_module.fstage_0.stage_1.subx.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_1.subx.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_1.suby.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_1.suby.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_1.subz.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_1.subz.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_1.subz.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_1.z_coeff  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_2.clk  = io_in[12];
	assign \mchip.cordic_module.fstage_0.stage_2.mode  = io_in[10];
	assign \mchip.cordic_module.fstage_0.stage_2.reset  = io_in[13];
	assign \mchip.cordic_module.fstage_0.stage_2.step_ctr  = {2'h0, \mchip.cordic_module.fstage_0.stage_0.step_ctr [2], 2'h2};
	assign \mchip.cordic_module.fstage_0.stage_2.subx.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_2.subx.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_2.suby.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_2.suby.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_2.subz.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_2.subz.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_2.subz.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_2.z_coeff  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_3.clk  = io_in[12];
	assign \mchip.cordic_module.fstage_0.stage_3.mode  = io_in[10];
	assign \mchip.cordic_module.fstage_0.stage_3.out_x  = {\mchip.cordic_module.next_x [16:6], 6'h00};
	assign \mchip.cordic_module.fstage_0.stage_3.reset  = io_in[13];
	assign \mchip.cordic_module.fstage_0.stage_3.step_ctr  = {2'h0, \mchip.cordic_module.fstage_0.stage_0.step_ctr [2], 2'h3};
	assign \mchip.cordic_module.fstage_0.stage_3.subx.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_3.subx.inside_add.out  = {\mchip.cordic_module.next_x [16:6], 6'h00};
	assign \mchip.cordic_module.fstage_0.stage_3.subx.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_3.subx.out  = {\mchip.cordic_module.next_x [16:6], 6'h00};
	assign \mchip.cordic_module.fstage_0.stage_3.suby.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_3.suby.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_3.subz.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_3.subz.inside_add.in_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_3.subz.modified_b  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.stage_3.z_coeff  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.step_ctr  = {2'h0, \mchip.cordic_module.fstage_0.stage_0.step_ctr [2], 2'h0};
	assign \mchip.cordic_module.fstage_0.z_coeff_0  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.z_coeff_1  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.z_coeff_2  = 17'h00000;
	assign \mchip.cordic_module.fstage_0.z_coeff_3  = 17'h00000;
	assign \mchip.cordic_module.in_val  = io_in[9:0];
	assign \mchip.cordic_module.in_val_32768  = {io_in[8:0], 8'h00};
	assign \mchip.cordic_module.in_x_32768  = {2'h0, io_in[9:5], 10'h000};
	assign \mchip.cordic_module.in_y_32768  = {2'h0, io_in[4:0], 10'h000};
	assign \mchip.cordic_module.init_x  = 17'h00000;
	assign \mchip.cordic_module.init_y  = 17'h00000;
	assign \mchip.cordic_module.init_z  = 17'h00000;
	assign \mchip.cordic_module.mode_toggle  = io_in[10];
	assign \mchip.cordic_module.next_x [5:0] = 6'h00;
	assign \mchip.cordic_module.out1 [5:0] = 6'h00;
	assign \mchip.cordic_module.out2 [5:0] = 6'h00;
	assign \mchip.cordic_module.out_toggle  = io_in[11];
	assign \mchip.cordic_module.rst  = io_in[13];
	assign \mchip.cordic_module.step_ctr_4  = {2'h0, \mchip.cordic_module.fstage_0.stage_0.step_ctr [2], 2'h0};
	assign \mchip.cordic_module.val  = io_out[10:0];
	assign \mchip.cordic_module.z_coeff[0]  = 17'h06488;
	assign \mchip.cordic_module.z_coeff[10]  = 17'h00020;
	assign \mchip.cordic_module.z_coeff[11]  = 17'h00010;
	assign \mchip.cordic_module.z_coeff[12]  = 17'h00008;
	assign \mchip.cordic_module.z_coeff[13]  = 17'h00004;
	assign \mchip.cordic_module.z_coeff[14]  = 17'h00002;
	assign \mchip.cordic_module.z_coeff[15]  = 17'h00001;
	assign \mchip.cordic_module.z_coeff[1]  = 17'h03b59;
	assign \mchip.cordic_module.z_coeff[2]  = 17'h01f5b;
	assign \mchip.cordic_module.z_coeff[3]  = 17'h00feb;
	assign \mchip.cordic_module.z_coeff[4]  = 17'h007fd;
	assign \mchip.cordic_module.z_coeff[5]  = 17'h00400;
	assign \mchip.cordic_module.z_coeff[6]  = 17'h00200;
	assign \mchip.cordic_module.z_coeff[7]  = 17'h00100;
	assign \mchip.cordic_module.z_coeff[8]  = 17'h00080;
	assign \mchip.cordic_module.z_coeff[9]  = 17'h00040;
	assign \mchip.cordic_module.z_coeff_group[0]  = 17'h00000;
	assign \mchip.cordic_module.z_coeff_group[1]  = 17'h00000;
	assign \mchip.cordic_module.z_coeff_group[2]  = 17'h00000;
	assign \mchip.cordic_module.z_coeff_group[3]  = 17'h00000;
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.cordic_module.done , io_out[10:0]};
	assign \mchip.reset  = io_in[13];
endmodule
module d14_siyuanl4_matrixcalc (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire [4:0] _2025_;
	wire [4:0] _2026_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [7:0] \mchip.data_in ;
	wire [4:0] \mchip.data_out ;
	wire \mchip.enter ;
	wire \mchip.error ;
	wire \mchip.finish ;
	wire [3:0] \mchip.index ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.matrix_calculator.add_finish ;
	wire [4:0] \mchip.matrix_calculator.add_logic.add1.S ;
	wire [4:0] \mchip.matrix_calculator.add_logic.add1_out ;
	wire [4:0] \mchip.matrix_calculator.add_logic.add2.S ;
	wire [4:0] \mchip.matrix_calculator.add_logic.add2_out ;
	wire \mchip.matrix_calculator.add_logic.clk ;
	wire \mchip.matrix_calculator.add_logic.finish ;
	wire \mchip.matrix_calculator.add_logic.fsm.clk ;
	reg [9:0] \mchip.matrix_calculator.add_logic.fsm.cur_state ;
	wire \mchip.matrix_calculator.add_logic.fsm.finish ;
	wire [63:0] \mchip.matrix_calculator.add_logic.fsm.mat_A ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_1 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_10 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_11 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_12 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_13 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_14 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_15 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_16 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_2 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_3 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_4 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_5 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_6 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_7 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_8 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_A_9 ;
	wire [63:0] \mchip.matrix_calculator.add_logic.fsm.mat_B ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_1 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_10 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_11 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_12 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_13 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_14 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_15 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_16 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_2 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_3 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_4 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_5 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_6 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_7 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_8 ;
	wire [3:0] \mchip.matrix_calculator.add_logic.fsm.mat_B_9 ;
	wire \mchip.matrix_calculator.add_logic.fsm.rst ;
	wire \mchip.matrix_calculator.add_logic.fsm.shift_en ;
	wire [63:0] \mchip.matrix_calculator.add_logic.mat_A ;
	wire [63:0] \mchip.matrix_calculator.add_logic.mat_B ;
	wire [159:0] \mchip.matrix_calculator.add_logic.mat_out ;
	wire \mchip.matrix_calculator.add_logic.rst ;
	wire [159:0] \mchip.matrix_calculator.add_logic.shift1.Q ;
	wire \mchip.matrix_calculator.add_logic.shift1.clock ;
	wire [19:0] \mchip.matrix_calculator.add_logic.shift1.data_in ;
	wire \mchip.matrix_calculator.add_logic.shift1.en ;
	wire \mchip.matrix_calculator.add_logic.shift1.rst ;
	wire \mchip.matrix_calculator.add_logic.shift_en ;
	wire [19:0] \mchip.matrix_calculator.add_logic.shift_in ;
	wire \mchip.matrix_calculator.add_logic.sign ;
	wire [159:0] \mchip.matrix_calculator.add_output ;
	wire \mchip.matrix_calculator.clk ;
	wire [7:0] \mchip.matrix_calculator.data_in ;
	wire [4:0] \mchip.matrix_calculator.data_out ;
	wire \mchip.matrix_calculator.ed_de.clk ;
	wire \mchip.matrix_calculator.ed_de.signal ;
	reg \mchip.matrix_calculator.ed_de.tmp1 ;
	wire \mchip.matrix_calculator.enter ;
	wire \mchip.matrix_calculator.error ;
	wire \mchip.matrix_calculator.finish ;
	wire \mchip.matrix_calculator.fsm.add_finish ;
	wire \mchip.matrix_calculator.fsm.clk ;
	reg [20:0] \mchip.matrix_calculator.fsm.cur_state ;
	wire \mchip.matrix_calculator.fsm.error ;
	wire \mchip.matrix_calculator.fsm.finish ;
	wire [1:0] \mchip.matrix_calculator.fsm.input_op ;
	wire \mchip.matrix_calculator.fsm.mul_finish ;
	wire \mchip.matrix_calculator.fsm.rst ;
	wire [3:0] \mchip.matrix_calculator.index ;
	wire [4:0] \mchip.matrix_calculator.index_count ;
	reg [4:0] \mchip.matrix_calculator.index_counter.Q ;
	wire \mchip.matrix_calculator.index_counter.clear ;
	wire \mchip.matrix_calculator.index_counter.clock ;
	wire \mchip.matrix_calculator.index_counter.en ;
	wire [127:0] \mchip.matrix_calculator.input_matrix ;
	wire [63:0] \mchip.matrix_calculator.input_matrix_A ;
	wire [63:0] \mchip.matrix_calculator.input_matrix_B ;
	wire [1:0] \mchip.matrix_calculator.input_op ;
	wire \mchip.matrix_calculator.mul_finish ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.add_in1 ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.add_in2 ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.add_in3 ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.add_in4 ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.add_in5 ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.add_in6 ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.add_in7 ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.add_in8 ;
	wire [9:0] \mchip.matrix_calculator.mul_logic.add_out ;
	wire [9:0] \mchip.matrix_calculator.mul_logic.add_out2 ;
	wire \mchip.matrix_calculator.mul_logic.clk ;
	wire \mchip.matrix_calculator.mul_logic.finish ;
	wire \mchip.matrix_calculator.mul_logic.fsm.clk ;
	reg [10:0] \mchip.matrix_calculator.mul_logic.fsm.cur_state ;
	wire \mchip.matrix_calculator.mul_logic.fsm.finish ;
	wire \mchip.matrix_calculator.mul_logic.fsm.layer_2_en ;
	wire [63:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_1 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_10 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_11 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_12 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_13 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_14 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_15 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_16 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_2 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_3 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_4 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_5 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_6 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_7 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_8 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_A_9 ;
	wire [63:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_1 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_10 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_11 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_12 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_13 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_14 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_15 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_16 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_2 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_3 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_4 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_5 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_6 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_7 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_8 ;
	wire [3:0] \mchip.matrix_calculator.mul_logic.fsm.mat_B_9 ;
	wire \mchip.matrix_calculator.mul_logic.fsm.rst ;
	wire [31:0] \mchip.matrix_calculator.mul_logic.layer_1_2_reg.D ;
	reg [31:0] \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q ;
	wire \mchip.matrix_calculator.mul_logic.layer_1_2_reg.clear ;
	wire \mchip.matrix_calculator.mul_logic.layer_1_2_reg.clock ;
	wire [31:0] \mchip.matrix_calculator.mul_logic.layer_1_reg.D ;
	reg [31:0] \mchip.matrix_calculator.mul_logic.layer_1_reg.Q ;
	wire \mchip.matrix_calculator.mul_logic.layer_1_reg.clear ;
	wire \mchip.matrix_calculator.mul_logic.layer_1_reg.clock ;
	wire \mchip.matrix_calculator.mul_logic.layer_2_en ;
	wire [63:0] \mchip.matrix_calculator.mul_logic.mat_A ;
	wire [63:0] \mchip.matrix_calculator.mul_logic.mat_B ;
	wire [159:0] \mchip.matrix_calculator.mul_logic.mat_out ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult1.S ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult1_out ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult2.S ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult2_out ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult3.S ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult3_out ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult4.S ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult4_out ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult5.S ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult5_out ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult6.S ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult6_out ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult7.S ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult7_out ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult8.S ;
	wire [7:0] \mchip.matrix_calculator.mul_logic.mult8_out ;
	wire \mchip.matrix_calculator.mul_logic.rst ;
	reg [159:0] \mchip.matrix_calculator.mul_logic.shift_register.Q ;
	wire \mchip.matrix_calculator.mul_logic.shift_register.clock ;
	wire [19:0] \mchip.matrix_calculator.mul_logic.shift_register.data_in ;
	wire \mchip.matrix_calculator.mul_logic.shift_register.en ;
	wire \mchip.matrix_calculator.mul_logic.shift_register.rst ;
	wire [159:0] \mchip.matrix_calculator.mul_output ;
	wire [1:0] \mchip.matrix_calculator.op_reg.D ;
	reg [1:0] \mchip.matrix_calculator.op_reg.Q ;
	wire \mchip.matrix_calculator.op_reg.clear ;
	wire \mchip.matrix_calculator.op_reg.clock ;
	wire \mchip.matrix_calculator.op_reg.en ;
	wire [1:0] \mchip.matrix_calculator.operation ;
	wire [159:0] \mchip.matrix_calculator.output_mux.I0 ;
	wire [159:0] \mchip.matrix_calculator.output_mux.I1 ;
	wire \mchip.matrix_calculator.output_mux.S ;
	wire \mchip.matrix_calculator.rst ;
	reg [127:0] \mchip.matrix_calculator.shift_register.Q ;
	wire \mchip.matrix_calculator.shift_register.clock ;
	wire [7:0] \mchip.matrix_calculator.shift_register.data_in ;
	wire \mchip.matrix_calculator.shift_register.en ;
	wire \mchip.matrix_calculator.shift_register.rst ;
	wire \mchip.matrix_calculator.sw ;
	wire \mchip.matrix_calculator.sw_de.clk ;
	wire \mchip.matrix_calculator.sw_de.signal ;
	reg \mchip.matrix_calculator.sw_de.tmp1 ;
	wire [1:0] \mchip.operation ;
	wire \mchip.reset ;
	wire \mchip.rst ;
	wire \mchip.sw ;
	wire \mchip.sync1.async ;
	wire \mchip.sync1.clock ;
	reg \mchip.sync1.sync ;
	reg \mchip.sync1.tmp1 ;
	wire \mchip.sync1.tmp2 ;
	wire \mchip.sync10.async ;
	wire \mchip.sync10.clock ;
	reg \mchip.sync10.sync ;
	reg \mchip.sync10.tmp1 ;
	wire \mchip.sync10.tmp2 ;
	wire \mchip.sync11.async ;
	wire \mchip.sync11.clock ;
	reg \mchip.sync11.sync ;
	reg \mchip.sync11.tmp1 ;
	wire \mchip.sync11.tmp2 ;
	wire \mchip.sync12.async ;
	wire \mchip.sync12.clock ;
	reg \mchip.sync12.sync ;
	reg \mchip.sync12.tmp1 ;
	wire \mchip.sync12.tmp2 ;
	wire \mchip.sync13.async ;
	wire \mchip.sync13.clock ;
	reg \mchip.sync13.sync ;
	reg \mchip.sync13.tmp1 ;
	wire \mchip.sync13.tmp2 ;
	wire \mchip.sync2.async ;
	wire \mchip.sync2.clock ;
	reg \mchip.sync2.sync ;
	reg \mchip.sync2.tmp1 ;
	wire \mchip.sync2.tmp2 ;
	wire \mchip.sync3.async ;
	wire \mchip.sync3.clock ;
	reg \mchip.sync3.sync ;
	reg \mchip.sync3.tmp1 ;
	wire \mchip.sync3.tmp2 ;
	wire \mchip.sync4.async ;
	wire \mchip.sync4.clock ;
	reg \mchip.sync4.sync ;
	reg \mchip.sync4.tmp1 ;
	wire \mchip.sync4.tmp2 ;
	wire \mchip.sync5.async ;
	wire \mchip.sync5.clock ;
	reg \mchip.sync5.sync ;
	reg \mchip.sync5.tmp1 ;
	wire \mchip.sync5.tmp2 ;
	wire \mchip.sync6.async ;
	wire \mchip.sync6.clock ;
	reg \mchip.sync6.sync ;
	reg \mchip.sync6.tmp1 ;
	wire \mchip.sync6.tmp2 ;
	wire \mchip.sync7.async ;
	wire \mchip.sync7.clock ;
	reg \mchip.sync7.sync ;
	reg \mchip.sync7.tmp1 ;
	wire \mchip.sync7.tmp2 ;
	wire \mchip.sync8.async ;
	wire \mchip.sync8.clock ;
	reg \mchip.sync8.sync ;
	reg \mchip.sync8.tmp1 ;
	wire \mchip.sync8.tmp2 ;
	wire \mchip.sync9.async ;
	wire \mchip.sync9.clock ;
	reg \mchip.sync9.sync ;
	reg \mchip.sync9.tmp1 ;
	wire \mchip.sync9.tmp2 ;
	assign _0605_ = (\mchip.matrix_calculator.op_reg.Q [0] ? _0603_ : _0604_);
	assign _0606_ = ~(\mchip.matrix_calculator.shift_register.Q [69] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0607_ = \mchip.matrix_calculator.shift_register.Q [77] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0608_ = _0606_ & ~_0607_;
	assign _0609_ = \mchip.matrix_calculator.shift_register.Q [93] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0610_ = \mchip.matrix_calculator.shift_register.Q [85] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0611_ = _0610_ | _0609_;
	assign _0612_ = _0608_ & ~_0611_;
	assign _0613_ = \mchip.matrix_calculator.shift_register.Q [125] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0614_ = \mchip.matrix_calculator.shift_register.Q [117] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0615_ = _0614_ | _0613_;
	assign _0616_ = \mchip.matrix_calculator.shift_register.Q [109] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0617_ = \mchip.matrix_calculator.shift_register.Q [101] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0618_ = _0617_ | _0616_;
	assign _0619_ = _0618_ | _0615_;
	assign _0620_ = _0612_ & ~_0619_;
	assign _0621_ = _1718_ & ~_0620_;
	assign _0622_ = _0621_ ^ _0605_;
	assign \mchip.matrix_calculator.add_logic.add1.S [1] = _0622_ ^ _0586_;
	assign _0623_ = _0621_ & _0605_;
	assign _0624_ = _0622_ & _0586_;
	assign _0625_ = _0624_ | _0623_;
	assign _0626_ = ~(\mchip.matrix_calculator.shift_register.Q [6] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0627_ = \mchip.matrix_calculator.shift_register.Q [14] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0628_ = _0626_ & ~_0627_;
	assign _0629_ = \mchip.matrix_calculator.shift_register.Q [30] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0630_ = \mchip.matrix_calculator.shift_register.Q [22] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0631_ = _0630_ | _0629_;
	assign _0632_ = _0628_ & ~_0631_;
	assign _0633_ = \mchip.matrix_calculator.shift_register.Q [62] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0634_ = \mchip.matrix_calculator.shift_register.Q [54] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0635_ = _0634_ | _0633_;
	assign _0636_ = \mchip.matrix_calculator.shift_register.Q [46] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0637_ = \mchip.matrix_calculator.shift_register.Q [38] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0638_ = _0637_ | _0636_;
	assign _0639_ = _0638_ | _0635_;
	assign _0640_ = _0632_ & ~_0639_;
	assign _0641_ = _1718_ & ~_0640_;
	assign _0642_ = ~_0641_;
	assign _0643_ = ~(_0602_ | _1751_);
	assign _0644_ = _0641_ ^ _0643_;
	assign _0645_ = (\mchip.matrix_calculator.op_reg.Q [0] ? _0642_ : _0644_);
	assign _0646_ = ~(\mchip.matrix_calculator.shift_register.Q [70] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0647_ = \mchip.matrix_calculator.shift_register.Q [78] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0648_ = _0646_ & ~_0647_;
	assign _0649_ = \mchip.matrix_calculator.shift_register.Q [94] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0650_ = \mchip.matrix_calculator.shift_register.Q [86] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0651_ = _0650_ | _0649_;
	assign _0652_ = _0648_ & ~_0651_;
	assign _0653_ = \mchip.matrix_calculator.shift_register.Q [126] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0654_ = \mchip.matrix_calculator.shift_register.Q [118] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0655_ = _0654_ | _0653_;
	assign _0656_ = \mchip.matrix_calculator.shift_register.Q [110] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0657_ = \mchip.matrix_calculator.shift_register.Q [102] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0658_ = _0657_ | _0656_;
	assign _0659_ = _0658_ | _0655_;
	assign _0660_ = _0652_ & ~_0659_;
	assign _0661_ = _1718_ & ~_0660_;
	assign _0662_ = _0661_ ^ _0645_;
	assign \mchip.matrix_calculator.add_logic.add1.S [2] = _0662_ ^ _0625_;
	assign _0663_ = _0661_ & _0645_;
	assign _0664_ = _0662_ & _0625_;
	assign _0665_ = _0664_ | _0663_;
	assign _0666_ = ~(\mchip.matrix_calculator.shift_register.Q [7] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0667_ = \mchip.matrix_calculator.shift_register.Q [15] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0668_ = _0666_ & ~_0667_;
	assign _0669_ = \mchip.matrix_calculator.shift_register.Q [31] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0670_ = \mchip.matrix_calculator.shift_register.Q [23] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0671_ = _0670_ | _0669_;
	assign _0672_ = _0668_ & ~_0671_;
	assign _0673_ = \mchip.matrix_calculator.shift_register.Q [63] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0674_ = \mchip.matrix_calculator.shift_register.Q [55] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0675_ = _0674_ | _0673_;
	assign _0676_ = \mchip.matrix_calculator.shift_register.Q [47] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0677_ = \mchip.matrix_calculator.shift_register.Q [39] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0678_ = _0677_ | _0676_;
	assign _0679_ = _0678_ | _0675_;
	assign _0680_ = _0672_ & ~_0679_;
	assign _0681_ = _1718_ & ~_0680_;
	assign _0682_ = _0641_ | ~_0643_;
	assign _0683_ = _0681_ ^ _0682_;
	assign _0684_ = (\mchip.matrix_calculator.op_reg.Q [0] ? _0681_ : _0683_);
	assign _0685_ = ~(\mchip.matrix_calculator.shift_register.Q [71] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0686_ = \mchip.matrix_calculator.shift_register.Q [79] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0687_ = _0685_ & ~_0686_;
	assign _0688_ = \mchip.matrix_calculator.shift_register.Q [95] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0689_ = \mchip.matrix_calculator.shift_register.Q [87] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0690_ = _0689_ | _0688_;
	assign _0691_ = _0687_ & ~_0690_;
	assign _0692_ = \mchip.matrix_calculator.shift_register.Q [127] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0693_ = \mchip.matrix_calculator.shift_register.Q [119] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0694_ = _0693_ | _0692_;
	assign _0695_ = \mchip.matrix_calculator.shift_register.Q [111] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0696_ = \mchip.matrix_calculator.shift_register.Q [103] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0697_ = _0696_ | _0695_;
	assign _0698_ = _0697_ | _0694_;
	assign _0699_ = _0691_ & ~_0698_;
	assign _0700_ = _1718_ & ~_0699_;
	assign _0701_ = ~(_0700_ ^ _0684_);
	assign \mchip.matrix_calculator.add_logic.add1.S [3] = _0701_ ^ _0665_;
	assign _0702_ = _0684_ | ~_0700_;
	assign _0703_ = _0701_ & _0663_;
	assign _0704_ = _0702_ & ~_0703_;
	assign _0705_ = ~(_0701_ & _0662_);
	assign _0706_ = _0625_ & ~_0705_;
	assign _0707_ = _0704_ & ~_0706_;
	assign _0708_ = _0681_ | _0641_;
	assign _0709_ = _0643_ & ~_0708_;
	assign _0710_ = _0582_ & ~_0709_;
	assign \mchip.matrix_calculator.add_logic.add1.S [4] = _0710_ ^ _0707_;
	assign _0711_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [72];
	assign _0712_ = \mchip.matrix_calculator.shift_register.Q [88] & ~_0445_;
	assign _0713_ = _0711_ & ~_0712_;
	assign _0714_ = \mchip.matrix_calculator.shift_register.Q [120] & ~_0440_;
	assign _0715_ = \mchip.matrix_calculator.shift_register.Q [104] & ~_0442_;
	assign _0716_ = _0715_ | _0714_;
	assign _0717_ = _0713_ & ~_0716_;
	assign _0718_ = ~(_0717_ | _0453_);
	assign _0719_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [36];
	assign _0720_ = \mchip.matrix_calculator.shift_register.Q [44] & ~_1815_;
	assign _0721_ = _0719_ & ~_0720_;
	assign _0722_ = _0721_ | _0042_;
	assign \mchip.matrix_calculator.mul_logic.mult2.S [0] = _0718_ & ~_0722_;
	assign _0723_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [68];
	assign _0724_ = \mchip.matrix_calculator.shift_register.Q [84] & ~_0445_;
	assign _0725_ = _0723_ & ~_0724_;
	assign _0726_ = \mchip.matrix_calculator.shift_register.Q [116] & ~_0440_;
	assign _0727_ = \mchip.matrix_calculator.shift_register.Q [100] & ~_0442_;
	assign _0728_ = _0727_ | _0726_;
	assign _0729_ = _0725_ & ~_0728_;
	assign _0730_ = ~(_0729_ | _0453_);
	assign _0731_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [16];
	assign _0732_ = \mchip.matrix_calculator.shift_register.Q [24] & ~_1815_;
	assign _0733_ = _0731_ & ~_0732_;
	assign _0734_ = _0733_ | _0042_;
	assign \mchip.matrix_calculator.mul_logic.mult7.S [0] = _0730_ & ~_0734_;
	assign _0735_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [64];
	assign _0736_ = \mchip.matrix_calculator.shift_register.Q [80] & ~_0445_;
	assign _0737_ = _0735_ & ~_0736_;
	assign _0738_ = \mchip.matrix_calculator.shift_register.Q [112] & ~_0440_;
	assign _0739_ = \mchip.matrix_calculator.shift_register.Q [96] & ~_0442_;
	assign _0740_ = _0739_ | _0738_;
	assign _0741_ = _0737_ & ~_0740_;
	assign _0742_ = ~(_0741_ | _0453_);
	assign _0743_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [0];
	assign _0744_ = \mchip.matrix_calculator.shift_register.Q [8] & ~_1815_;
	assign _0745_ = _0743_ & ~_0744_;
	assign _0746_ = _0745_ | _0042_;
	assign \mchip.matrix_calculator.mul_logic.mult8.S [0] = _0742_ & ~_0746_;
	assign _0747_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [32];
	assign _0748_ = \mchip.matrix_calculator.shift_register.Q [40] & ~_1815_;
	assign _0749_ = _0747_ & ~_0748_;
	assign _0750_ = _0749_ | _0042_;
	assign \mchip.matrix_calculator.mul_logic.mult6.S [0] = _0718_ & ~_0750_;
	assign _0751_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [48];
	assign _0752_ = \mchip.matrix_calculator.shift_register.Q [56] & ~_1815_;
	assign _0753_ = _0751_ & ~_0752_;
	assign _0754_ = _0753_ | _0042_;
	assign \mchip.matrix_calculator.mul_logic.mult5.S [0] = _0454_ & ~_0754_;
	assign _0755_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [4];
	assign _0756_ = \mchip.matrix_calculator.shift_register.Q [12] & ~_1815_;
	assign _0757_ = _0755_ & ~_0756_;
	assign _0758_ = _0757_ | _0042_;
	assign \mchip.matrix_calculator.mul_logic.mult4.S [0] = _0742_ & ~_0758_;
	assign _0759_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [20];
	assign _0760_ = \mchip.matrix_calculator.shift_register.Q [28] & ~_1815_;
	assign _0761_ = _0759_ & ~_0760_;
	assign _0762_ = _0761_ | _0042_;
	assign \mchip.matrix_calculator.mul_logic.mult3.S [0] = _0730_ & ~_0762_;
	assign _0763_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [24] ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [16];
	assign _0764_ = ~(_0763_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [0]);
	assign _0765_ = _0763_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [0];
	assign _0766_ = ~(_0765_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [8]);
	assign _0767_ = ~(_0766_ & _0764_);
	assign _0768_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [24] & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [16];
	assign _0769_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [25] ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [17]);
	assign _0770_ = ~(_0769_ ^ _0768_);
	assign _0771_ = _0770_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [1];
	assign _0772_ = _0771_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [9];
	assign _0773_ = _0772_ & _0767_;
	assign _0774_ = ~(_0770_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [1]);
	assign _0775_ = ~(_0771_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [9]);
	assign _0776_ = ~(_0775_ & _0774_);
	assign _0777_ = _0768_ & ~_0769_;
	assign _0778_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [25] & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [17];
	assign _0779_ = _0778_ | _0777_;
	assign _0780_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [26] ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [18]);
	assign _0781_ = ~(_0780_ ^ _0779_);
	assign _0782_ = _0781_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [2];
	assign _0783_ = _0782_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [10];
	assign _0784_ = ~(_0783_ ^ _0776_);
	assign \mchip.matrix_calculator.mul_logic.add_out [2] = ~(_0784_ ^ _0773_);
	assign _0785_ = _0783_ & _0776_;
	assign _0786_ = _0773_ & ~_0784_;
	assign _0787_ = ~(_0786_ | _0785_);
	assign _0788_ = _0781_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [2];
	assign _0789_ = _0782_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [10];
	assign _0790_ = _0789_ | _0788_;
	assign _0791_ = ~\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [3];
	assign _0792_ = _0780_ | ~_0779_;
	assign _0793_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [26] & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [18];
	assign _0794_ = _0792_ & ~_0793_;
	assign _0795_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [27] ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [19]);
	assign _0796_ = _0795_ ^ _0794_;
	assign _0797_ = _0796_ ^ _0791_;
	assign _0798_ = _0797_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [11];
	assign _0799_ = _0798_ ^ _0790_;
	assign \mchip.matrix_calculator.mul_logic.add_out [3] = _0799_ ^ _0787_;
	assign _0800_ = _0790_ & ~_0798_;
	assign _0801_ = _0785_ & ~_0799_;
	assign _0802_ = _0801_ | _0800_;
	assign _0803_ = _0799_ | _0784_;
	assign _0804_ = _0773_ & ~_0803_;
	assign _0805_ = _0804_ | _0802_;
	assign _0806_ = _0796_ & ~_0791_;
	assign _0807_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [11] & ~_0797_;
	assign _0808_ = _0807_ | _0806_;
	assign _0809_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [27] & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [19];
	assign _0810_ = _0793_ & ~_0795_;
	assign _0811_ = _0810_ | _0809_;
	assign _0812_ = _0795_ | _0780_;
	assign _0813_ = _0779_ & ~_0812_;
	assign _0814_ = _0813_ | _0811_;
	assign _0815_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [28] ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [20]);
	assign _0816_ = ~(_0815_ ^ _0814_);
	assign _0817_ = _0816_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [4];
	assign _0818_ = _0817_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [12];
	assign _0819_ = ~(_0818_ ^ _0808_);
	assign \mchip.matrix_calculator.mul_logic.add_out [4] = ~(_0819_ ^ _0805_);
	assign _0820_ = _0818_ & _0808_;
	assign _0821_ = _0805_ & ~_0819_;
	assign _0822_ = ~(_0821_ | _0820_);
	assign _0823_ = _0816_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [4];
	assign _0824_ = _0817_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [12];
	assign _0825_ = _0824_ | _0823_;
	assign _0826_ = ~\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [5];
	assign _0827_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [28] & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [20];
	assign _0828_ = _0814_ & ~_0815_;
	assign _0829_ = ~(_0828_ | _0827_);
	assign _0830_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [29] ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [21]);
	assign _0831_ = _0830_ ^ _0829_;
	assign _0832_ = _0831_ ^ _0826_;
	assign _0833_ = _0832_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [13];
	assign _0834_ = _0833_ ^ _0825_;
	assign \mchip.matrix_calculator.mul_logic.add_out [5] = _0834_ ^ _0822_;
	assign _0835_ = _0834_ | _0819_;
	assign _0836_ = _0805_ & ~_0835_;
	assign _0837_ = _0825_ & ~_0833_;
	assign _0838_ = _0820_ & ~_0834_;
	assign _0839_ = _0838_ | _0837_;
	assign _0840_ = _0839_ | _0836_;
	assign _0841_ = _0831_ & ~_0826_;
	assign _0842_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [13] & ~_0832_;
	assign _0843_ = _0842_ | _0841_;
	assign _0844_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [29] & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [21];
	assign _0845_ = _0827_ & ~_0830_;
	assign _0846_ = _0845_ | _0844_;
	assign _0847_ = _0830_ | _0815_;
	assign _0848_ = _0814_ & ~_0847_;
	assign _0849_ = _0848_ | _0846_;
	assign _0850_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [30] ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [22];
	assign _0851_ = _0850_ ^ _0849_;
	assign _0852_ = _0851_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [6];
	assign _0853_ = _0852_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [14];
	assign _0854_ = ~(_0853_ ^ _0843_);
	assign \mchip.matrix_calculator.mul_logic.add_out [6] = ~(_0854_ ^ _0840_);
	assign _0855_ = _0853_ & _0843_;
	assign _0856_ = _0840_ & ~_0854_;
	assign _0857_ = ~(_0856_ | _0855_);
	assign _0858_ = ~(_0851_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [6]);
	assign _0859_ = _0852_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [14];
	assign _0860_ = _0858_ & ~_0859_;
	assign _0861_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [30] & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [22];
	assign _0862_ = _0850_ & _0849_;
	assign _0863_ = _0862_ | _0861_;
	assign _0864_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [31] ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [23];
	assign _0865_ = _0864_ ^ _0863_;
	assign _0866_ = _0865_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [7];
	assign _0867_ = _0866_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [15];
	assign _0868_ = _0867_ ^ _0860_;
	assign \mchip.matrix_calculator.mul_logic.add_out [7] = _0868_ ^ _0857_;
	assign _0869_ = _0860_ | ~_0867_;
	assign _0870_ = _0855_ & ~_0868_;
	assign _0871_ = _0869_ & ~_0870_;
	assign _0872_ = _0868_ | _0854_;
	assign _0873_ = _0839_ & ~_0872_;
	assign _0874_ = _0871_ & ~_0873_;
	assign _0875_ = _0872_ | _0835_;
	assign _0876_ = _0805_ & ~_0875_;
	assign _0877_ = _0876_ | ~_0874_;
	assign _0878_ = ~(_0865_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [7]);
	assign _0879_ = ~(_0866_ & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [15]);
	assign _0880_ = ~(_0879_ & _0878_);
	assign _0881_ = ~(_0864_ & _0850_);
	assign _0882_ = _0881_ | _0847_;
	assign _0883_ = _0882_ | ~_0814_;
	assign _0884_ = _0846_ & ~_0881_;
	assign _0885_ = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [31] & \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [23];
	assign _0886_ = _0864_ & _0861_;
	assign _0887_ = _0886_ | _0885_;
	assign _0888_ = _0887_ | _0884_;
	assign _0889_ = _0883_ & ~_0888_;
	assign _0890_ = _0889_ ^ _0880_;
	assign \mchip.matrix_calculator.mul_logic.add_out [8] = ~(_0890_ ^ _0877_);
	assign \mchip.matrix_calculator.mul_logic.add_out [1] = _0772_ ^ _0767_;
	assign _0891_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [24] ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [16];
	assign _0892_ = ~(_0891_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [0]);
	assign _0893_ = _0891_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [0];
	assign _0894_ = ~(_0893_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [8]);
	assign _0895_ = ~(_0894_ & _0892_);
	assign _0896_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [24] & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [16];
	assign _0897_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [25] ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [17]);
	assign _0898_ = ~(_0897_ ^ _0896_);
	assign _0899_ = _0898_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [1];
	assign _0900_ = _0899_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [9];
	assign \mchip.matrix_calculator.mul_logic.add_out2 [1] = _0900_ ^ _0895_;
	assign _0901_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [21];
	assign _0902_ = \mchip.matrix_calculator.shift_register.Q [29] & ~_1815_;
	assign _0903_ = _0901_ & ~_0902_;
	assign _0904_ = _0903_ | _0042_;
	assign _0905_ = _0730_ & ~_0904_;
	assign _0906_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [69];
	assign _0907_ = \mchip.matrix_calculator.shift_register.Q [85] & ~_0445_;
	assign _0908_ = _0906_ & ~_0907_;
	assign _0909_ = \mchip.matrix_calculator.shift_register.Q [117] & ~_0440_;
	assign _0910_ = \mchip.matrix_calculator.shift_register.Q [101] & ~_0442_;
	assign _0911_ = _0910_ | _0909_;
	assign _0912_ = _0908_ & ~_0911_;
	assign _0913_ = _0912_ | _0453_;
	assign _0914_ = _0913_ | _0762_;
	assign \mchip.matrix_calculator.mul_logic.mult3.S [1] = ~(_0914_ ^ _0905_);
	assign _0915_ = _0905_ & ~_0914_;
	assign _0916_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [22];
	assign _0917_ = \mchip.matrix_calculator.shift_register.Q [30] & ~_1815_;
	assign _0918_ = _0916_ & ~_0917_;
	assign _0919_ = _0918_ | _0042_;
	assign _0920_ = _0919_ | ~_0730_;
	assign _0921_ = ~(_0913_ | _0904_);
	assign _0922_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [70];
	assign _0923_ = \mchip.matrix_calculator.shift_register.Q [86] & ~_0445_;
	assign _0924_ = _0922_ & ~_0923_;
	assign _0925_ = \mchip.matrix_calculator.shift_register.Q [118] & ~_0440_;
	assign _0926_ = \mchip.matrix_calculator.shift_register.Q [102] & ~_0442_;
	assign _0927_ = _0926_ | _0925_;
	assign _0928_ = _0924_ & ~_0927_;
	assign _0929_ = _0928_ | _0453_;
	assign _0930_ = _0929_ | _0762_;
	assign _0931_ = _0930_ ^ _0921_;
	assign _0932_ = ~(_0931_ ^ _0920_);
	assign \mchip.matrix_calculator.mul_logic.mult3.S [2] = ~(_0932_ ^ _0915_);
	assign _0933_ = _0915_ & ~_0932_;
	assign _0934_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [23];
	assign _0935_ = \mchip.matrix_calculator.shift_register.Q [31] & ~_1815_;
	assign _0936_ = _0934_ & ~_0935_;
	assign _0937_ = _0936_ | _0042_;
	assign _0938_ = _0730_ & ~_0937_;
	assign _0939_ = _0931_ | _0920_;
	assign _0940_ = _0921_ & ~_0930_;
	assign _0941_ = _0939_ & ~_0940_;
	assign _0942_ = ~(_0919_ | _0913_);
	assign _0943_ = ~(_0929_ | _0904_);
	assign _0944_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [71];
	assign _0945_ = \mchip.matrix_calculator.shift_register.Q [87] & ~_0445_;
	assign _0946_ = _0944_ & ~_0945_;
	assign _0947_ = \mchip.matrix_calculator.shift_register.Q [119] & ~_0440_;
	assign _0948_ = \mchip.matrix_calculator.shift_register.Q [103] & ~_0442_;
	assign _0949_ = _0948_ | _0947_;
	assign _0950_ = _0946_ & ~_0949_;
	assign _0951_ = _0950_ | _0453_;
	assign _0952_ = _0951_ | _0762_;
	assign _0953_ = _0952_ ^ _0943_;
	assign _0954_ = _0953_ ^ _0942_;
	assign _0955_ = ~(_0954_ ^ _0941_);
	assign _0956_ = _0955_ ^ _0938_;
	assign \mchip.matrix_calculator.mul_logic.mult3.S [3] = ~(_0956_ ^ _0933_);
	assign _0957_ = _0933_ & ~_0956_;
	assign _0958_ = ~(_0954_ | _0941_);
	assign _0959_ = _0938_ & ~_0955_;
	assign _0960_ = _0959_ | _0958_;
	assign _0961_ = ~(_0937_ | _0913_);
	assign _0962_ = _0953_ | ~_0942_;
	assign _0963_ = _0943_ & ~_0952_;
	assign _0964_ = _0963_ | ~_0962_;
	assign _0965_ = _0929_ | _0919_;
	assign _0966_ = ~(_0951_ | _0904_);
	assign _0967_ = _0966_ ^ _0965_;
	assign _0968_ = _0967_ ^ _0964_;
	assign _0969_ = ~(_0968_ ^ _0961_);
	assign _0970_ = ~(_0969_ ^ _0960_);
	assign \mchip.matrix_calculator.mul_logic.mult3.S [4] = ~(_0970_ ^ _0957_);
	assign _0971_ = _0969_ & _0960_;
	assign _0972_ = _0957_ & ~_0970_;
	assign _0973_ = ~(_0972_ | _0971_);
	assign _0974_ = _0961_ & ~_0968_;
	assign _0975_ = _0964_ & ~_0967_;
	assign _0976_ = _0975_ | _0974_;
	assign _0977_ = ~(_0937_ | _0929_);
	assign _0978_ = _0965_ | ~_0966_;
	assign _0979_ = ~(_0951_ | _0919_);
	assign _0980_ = _0979_ ^ _0978_;
	assign _0981_ = ~(_0980_ ^ _0977_);
	assign _0982_ = ~(_0981_ ^ _0976_);
	assign \mchip.matrix_calculator.mul_logic.mult3.S [5] = _0982_ ^ _0973_;
	assign _0983_ = _0981_ & _0976_;
	assign _0984_ = _0971_ & ~_0982_;
	assign _0985_ = _0984_ | _0983_;
	assign _0986_ = _0982_ | _0970_;
	assign _0987_ = _0957_ & ~_0986_;
	assign _0988_ = _0987_ | _0985_;
	assign _0989_ = _0977_ & ~_0980_;
	assign _0990_ = _0979_ & ~_0978_;
	assign _0991_ = _0990_ | _0989_;
	assign _0992_ = ~(_0951_ | _0937_);
	assign _0993_ = _0992_ ^ _0991_;
	assign \mchip.matrix_calculator.mul_logic.mult3.S [6] = _0993_ ^ _0988_;
	assign _0994_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [73];
	assign _0995_ = \mchip.matrix_calculator.shift_register.Q [89] & ~_0445_;
	assign _0996_ = _0994_ & ~_0995_;
	assign _0997_ = \mchip.matrix_calculator.shift_register.Q [121] & ~_0440_;
	assign _0998_ = \mchip.matrix_calculator.shift_register.Q [105] & ~_0442_;
	assign _0999_ = _0998_ | _0997_;
	assign _1000_ = _0996_ & ~_0999_;
	assign _1001_ = _1000_ | _0453_;
	assign _1002_ = ~(_1001_ | _0750_);
	assign _1003_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [33];
	assign _1004_ = \mchip.matrix_calculator.shift_register.Q [41] & ~_1815_;
	assign _1005_ = _1003_ & ~_1004_;
	assign _1006_ = _1005_ | _0042_;
	assign _1007_ = _1006_ | ~_0718_;
	assign _1008_ = _1002_ & ~_1007_;
	assign _1009_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [34];
	assign _1010_ = \mchip.matrix_calculator.shift_register.Q [42] & ~_1815_;
	assign _1011_ = _1009_ & ~_1010_;
	assign _1012_ = _1011_ | _0042_;
	assign _1013_ = _0718_ & ~_1012_;
	assign _1014_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [74];
	assign _1015_ = \mchip.matrix_calculator.shift_register.Q [90] & ~_0445_;
	assign _1016_ = _1014_ & ~_1015_;
	assign _1017_ = \mchip.matrix_calculator.shift_register.Q [122] & ~_0440_;
	assign _1018_ = \mchip.matrix_calculator.shift_register.Q [106] & ~_0442_;
	assign _1019_ = _1018_ | _1017_;
	assign _1020_ = _1016_ & ~_1019_;
	assign _1021_ = _1020_ | _0453_;
	assign _1022_ = ~(_1021_ | _0750_);
	assign _1023_ = _1022_ ^ _1013_;
	assign _1024_ = ~(_1006_ | _1001_);
	assign _1025_ = ~(_1024_ ^ _1023_);
	assign _1026_ = _1008_ & ~_1025_;
	assign _1027_ = _1024_ & _1023_;
	assign _1028_ = ~(_1021_ | _1006_);
	assign _1029_ = _1022_ & _1013_;
	assign _1030_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [75];
	assign _1031_ = \mchip.matrix_calculator.shift_register.Q [91] & ~_0445_;
	assign _1032_ = _1030_ & ~_1031_;
	assign _1033_ = \mchip.matrix_calculator.shift_register.Q [123] & ~_0440_;
	assign _1034_ = \mchip.matrix_calculator.shift_register.Q [107] & ~_0442_;
	assign _1035_ = _1034_ | _1033_;
	assign _1036_ = _1032_ & ~_1035_;
	assign _1037_ = _1036_ | _0453_;
	assign _1038_ = _1037_ | _0750_;
	assign _1039_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [35];
	assign _1040_ = \mchip.matrix_calculator.shift_register.Q [43] & ~_1815_;
	assign _1041_ = _1039_ & ~_1040_;
	assign _1042_ = _1041_ | _0042_;
	assign _1043_ = _0718_ & ~_1042_;
	assign _1044_ = _1012_ | _1001_;
	assign _1045_ = _1044_ ^ _1043_;
	assign _1046_ = ~(_1045_ ^ _1038_);
	assign _1047_ = _1046_ ^ _1029_;
	assign _1048_ = _1047_ ^ _1028_;
	assign _1049_ = _1048_ ^ _1027_;
	assign \mchip.matrix_calculator.mul_logic.mult6.S [3] = ~(_1049_ ^ _1026_);
	assign _1050_ = _1026_ & ~_1049_;
	assign _1051_ = _1027_ & ~_1048_;
	assign _1052_ = _1051_ | _1050_;
	assign _1053_ = _1028_ & ~_1047_;
	assign _1054_ = _1029_ & ~_1046_;
	assign _1055_ = _1054_ | _1053_;
	assign _1056_ = ~(_1037_ | _1006_);
	assign _1057_ = _1045_ | _1038_;
	assign _1058_ = _1043_ & ~_1044_;
	assign _1059_ = _1058_ | ~_1057_;
	assign _1060_ = ~(_1042_ | _1001_);
	assign _1061_ = _1021_ | _1012_;
	assign _1062_ = _1061_ ^ _1060_;
	assign _1063_ = _1062_ ^ _1059_;
	assign _1064_ = ~(_1063_ ^ _1056_);
	assign _1065_ = ~(_1064_ ^ _1055_);
	assign \mchip.matrix_calculator.mul_logic.mult6.S [4] = ~(_1065_ ^ _1052_);
	assign _1066_ = _1064_ & _1055_;
	assign _1067_ = _1052_ & ~_1065_;
	assign _1068_ = ~(_1067_ | _1066_);
	assign _1069_ = _1056_ & ~_1063_;
	assign _1070_ = _1059_ & ~_1062_;
	assign _1071_ = _1070_ | _1069_;
	assign _1072_ = _1060_ & ~_1061_;
	assign _1073_ = ~(_1042_ | _1021_);
	assign _1074_ = ~(_1037_ | _1012_);
	assign _1075_ = _1074_ ^ _1073_;
	assign _1076_ = _1075_ ^ _1072_;
	assign _1077_ = ~(_1076_ ^ _1071_);
	assign \mchip.matrix_calculator.mul_logic.mult6.S [5] = _1077_ ^ _1068_;
	assign _1078_ = _1076_ & _1071_;
	assign _1079_ = _1066_ & ~_1077_;
	assign _1080_ = _1079_ | _1078_;
	assign _1081_ = _1077_ | _1065_;
	assign _1082_ = _1052_ & ~_1081_;
	assign _1083_ = _1082_ | _1080_;
	assign _1084_ = ~(_1075_ & _1072_);
	assign _1085_ = ~(_1074_ & _1073_);
	assign _1086_ = ~(_1042_ | _1037_);
	assign _1087_ = ~(_1086_ ^ _1085_);
	assign _1088_ = ~(_1087_ ^ _1084_);
	assign \mchip.matrix_calculator.mul_logic.mult6.S [6] = _1088_ ^ _1083_;
	assign _1089_ = _1085_ | ~_1086_;
	assign _1090_ = _1084_ | ~_1087_;
	assign _1091_ = _1088_ & _1083_;
	assign _1092_ = _1090_ & ~_1091_;
	assign \mchip.matrix_calculator.mul_logic.mult6.S [7] = _1092_ ^ _1089_;
	assign \mchip.matrix_calculator.mul_logic.mult6.S [2] = ~(_1025_ ^ _1008_);
	assign \mchip.matrix_calculator.mul_logic.mult6.S [1] = ~(_1007_ ^ _1002_);
	assign \mchip.matrix_calculator.mul_logic.add_out [0] = _0765_ ^ \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [8];
	assign _1093_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [1];
	assign _1094_ = \mchip.matrix_calculator.shift_register.Q [9] & ~_1815_;
	assign _1095_ = _1093_ & ~_1094_;
	assign _1096_ = _1095_ | _0042_;
	assign _1097_ = _0742_ & ~_1096_;
	assign _1098_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [65];
	assign _1099_ = \mchip.matrix_calculator.shift_register.Q [81] & ~_0445_;
	assign _1100_ = _1098_ & ~_1099_;
	assign _1101_ = \mchip.matrix_calculator.shift_register.Q [113] & ~_0440_;
	assign _1102_ = \mchip.matrix_calculator.shift_register.Q [97] & ~_0442_;
	assign _1103_ = _1102_ | _1101_;
	assign _1104_ = _1100_ & ~_1103_;
	assign _1105_ = _1104_ | _0453_;
	assign _1106_ = _1105_ | _0746_;
	assign \mchip.matrix_calculator.mul_logic.mult8.S [1] = ~(_1106_ ^ _1097_);
	assign _1107_ = _1097_ & ~_1106_;
	assign _1108_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [2];
	assign _1109_ = \mchip.matrix_calculator.shift_register.Q [10] & ~_1815_;
	assign _1110_ = _1108_ & ~_1109_;
	assign _1111_ = _1110_ | _0042_;
	assign _1112_ = _0742_ & ~_1111_;
	assign _1113_ = ~(_1105_ | _1096_);
	assign _1114_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [66];
	assign _1115_ = \mchip.matrix_calculator.shift_register.Q [82] & ~_0445_;
	assign _1116_ = _1114_ & ~_1115_;
	assign _1117_ = \mchip.matrix_calculator.shift_register.Q [114] & ~_0440_;
	assign _1118_ = \mchip.matrix_calculator.shift_register.Q [98] & ~_0442_;
	assign _1119_ = _1118_ | _1117_;
	assign _1120_ = _1116_ & ~_1119_;
	assign _1121_ = _1120_ | _0453_;
	assign _1122_ = _1121_ | _0746_;
	assign _1123_ = _1122_ ^ _1113_;
	assign _1124_ = _1123_ ^ _1112_;
	assign \mchip.matrix_calculator.mul_logic.mult8.S [2] = ~(_1124_ ^ _1107_);
	assign _1125_ = _1107_ & ~_1124_;
	assign _1126_ = _1123_ | ~_1112_;
	assign _1127_ = _1113_ & ~_1122_;
	assign _1128_ = _1127_ | ~_1126_;
	assign _1129_ = ~(_1121_ | _1096_);
	assign _1130_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [67];
	assign _1131_ = \mchip.matrix_calculator.shift_register.Q [83] & ~_0445_;
	assign _1132_ = _1130_ & ~_1131_;
	assign _1133_ = \mchip.matrix_calculator.shift_register.Q [115] & ~_0440_;
	assign _1134_ = \mchip.matrix_calculator.shift_register.Q [99] & ~_0442_;
	assign _1135_ = _1134_ | _1133_;
	assign _1136_ = _1132_ & ~_1135_;
	assign _1137_ = _1136_ | _0453_;
	assign _1138_ = ~(_1137_ | _0746_);
	assign _1139_ = _1138_ ^ _1129_;
	assign _1140_ = _1111_ | _1105_;
	assign _1141_ = _1140_ ^ _1139_;
	assign _1142_ = ~(_1141_ ^ _1128_);
	assign _1143_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [3];
	assign _1144_ = \mchip.matrix_calculator.shift_register.Q [11] & ~_1815_;
	assign _1145_ = _1143_ & ~_1144_;
	assign _1146_ = _1145_ | _0042_;
	assign _1147_ = _0742_ & ~_1146_;
	assign _1148_ = ~_1147_;
	assign _1149_ = _1148_ ^ _1142_;
	assign _1150_ = _1125_ & ~_1149_;
	assign _1151_ = _1128_ & ~_1141_;
	assign _1152_ = _1142_ & ~_1148_;
	assign _1153_ = _1152_ | _1151_;
	assign _1154_ = ~(_1146_ | _1105_);
	assign _1155_ = ~(_1138_ & _1129_);
	assign _1156_ = _1139_ & ~_1140_;
	assign _1157_ = _1156_ | ~_1155_;
	assign _1158_ = _1121_ | _1111_;
	assign _1159_ = ~(_1137_ | _1096_);
	assign _1160_ = _1159_ ^ _1158_;
	assign _1161_ = _1160_ ^ _1157_;
	assign _1162_ = ~(_1161_ ^ _1154_);
	assign _1163_ = ~(_1162_ ^ _1153_);
	assign \mchip.matrix_calculator.mul_logic.mult8.S [4] = ~(_1163_ ^ _1150_);
	assign _1164_ = _1162_ & _1153_;
	assign _1165_ = _1150_ & ~_1163_;
	assign _1166_ = ~(_1165_ | _1164_);
	assign _1167_ = _1154_ & ~_1161_;
	assign _1168_ = _1157_ & ~_1160_;
	assign _1169_ = _1168_ | _1167_;
	assign _1170_ = ~(_1146_ | _1121_);
	assign _1171_ = _1158_ | ~_1159_;
	assign _1172_ = ~(_1137_ | _1111_);
	assign _1173_ = _1172_ ^ _1171_;
	assign _1174_ = ~(_1173_ ^ _1170_);
	assign _1175_ = ~(_1174_ ^ _1169_);
	assign \mchip.matrix_calculator.mul_logic.mult8.S [5] = _1175_ ^ _1166_;
	assign _1176_ = _1174_ & _1169_;
	assign _1177_ = _1164_ & ~_1175_;
	assign _1178_ = _1177_ | _1176_;
	assign _1179_ = _1175_ | _1163_;
	assign _1180_ = _1150_ & ~_1179_;
	assign _1181_ = _1180_ | _1178_;
	assign _1182_ = _1170_ & ~_1173_;
	assign _1183_ = _1172_ & ~_1171_;
	assign _1184_ = _1183_ | _1182_;
	assign _1185_ = ~(_1146_ | _1137_);
	assign _1186_ = _1185_ ^ _1184_;
	assign \mchip.matrix_calculator.mul_logic.mult8.S [6] = _1186_ ^ _1181_;
	assign \mchip.matrix_calculator.mul_logic.mult8.S [3] = ~(_1149_ ^ _1125_);
	assign _1187_ = _0900_ & _0895_;
	assign _1188_ = ~(_0898_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [1]);
	assign _1189_ = ~(_0899_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [9]);
	assign _1190_ = ~(_1189_ & _1188_);
	assign _1191_ = _0896_ & ~_0897_;
	assign _1192_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [25] & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [17];
	assign _1193_ = _1192_ | _1191_;
	assign _1194_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [26] ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [18]);
	assign _1195_ = ~(_1194_ ^ _1193_);
	assign _1196_ = _1195_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [2];
	assign _1197_ = _1196_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [10];
	assign _1198_ = ~(_1197_ ^ _1190_);
	assign \mchip.matrix_calculator.mul_logic.add_out2 [2] = ~(_1198_ ^ _1187_);
	assign _1199_ = _1197_ & _1190_;
	assign _1200_ = _1187_ & ~_1198_;
	assign _1201_ = ~(_1200_ | _1199_);
	assign _1202_ = _1195_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [2];
	assign _1203_ = _1196_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [10];
	assign _1204_ = _1203_ | _1202_;
	assign _1205_ = ~\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [3];
	assign _1206_ = _1194_ | ~_1193_;
	assign _1207_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [26] & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [18];
	assign _1208_ = _1206_ & ~_1207_;
	assign _1209_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [27] ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [19]);
	assign _1210_ = _1209_ ^ _1208_;
	assign _1211_ = _1210_ ^ _1205_;
	assign _1212_ = _1211_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [11];
	assign _1213_ = _1212_ ^ _1204_;
	assign \mchip.matrix_calculator.mul_logic.add_out2 [3] = _1213_ ^ _1201_;
	assign _1214_ = _1204_ & ~_1212_;
	assign _1215_ = _1199_ & ~_1213_;
	assign _1216_ = _1215_ | _1214_;
	assign _1217_ = _1213_ | _1198_;
	assign _1218_ = _1187_ & ~_1217_;
	assign _1219_ = _1218_ | _1216_;
	assign _1220_ = _1210_ & ~_1205_;
	assign _1221_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [11] & ~_1211_;
	assign _1222_ = _1221_ | _1220_;
	assign _1223_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [27] & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [19];
	assign _1224_ = _1207_ & ~_1209_;
	assign _1225_ = _1224_ | _1223_;
	assign _1226_ = _1209_ | _1194_;
	assign _1227_ = _1193_ & ~_1226_;
	assign _1228_ = _1227_ | _1225_;
	assign _1229_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [28] ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [20]);
	assign _1230_ = ~(_1229_ ^ _1228_);
	assign _1231_ = _1230_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [4];
	assign _1232_ = _1231_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [12];
	assign _1233_ = ~(_1232_ ^ _1222_);
	assign \mchip.matrix_calculator.mul_logic.add_out2 [4] = ~(_1233_ ^ _1219_);
	assign _1234_ = _1232_ & _1222_;
	assign _1235_ = _1219_ & ~_1233_;
	assign _1236_ = ~(_1235_ | _1234_);
	assign _1237_ = _1230_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [4];
	assign _1238_ = _1231_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [12];
	assign _1239_ = _1238_ | _1237_;
	assign _1240_ = ~\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [5];
	assign _1241_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [28] & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [20];
	assign _1242_ = _1228_ & ~_1229_;
	assign _1243_ = ~(_1242_ | _1241_);
	assign _1244_ = ~(\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [29] ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [21]);
	assign _1245_ = _1244_ ^ _1243_;
	assign _1246_ = _1245_ ^ _1240_;
	assign _1247_ = _1246_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [13];
	assign _1248_ = _1247_ ^ _1239_;
	assign \mchip.matrix_calculator.mul_logic.add_out2 [5] = _1248_ ^ _1236_;
	assign _1249_ = _1248_ | _1233_;
	assign _1250_ = _1219_ & ~_1249_;
	assign _1251_ = _1239_ & ~_1247_;
	assign _1252_ = _1234_ & ~_1248_;
	assign _1253_ = _1252_ | _1251_;
	assign _1254_ = _1253_ | _1250_;
	assign _1255_ = _1245_ & ~_1240_;
	assign _1256_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [13] & ~_1246_;
	assign _1257_ = _1256_ | _1255_;
	assign _1258_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [29] & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [21];
	assign _1259_ = _1241_ & ~_1244_;
	assign _1260_ = _1259_ | _1258_;
	assign _1261_ = _1244_ | _1229_;
	assign _1262_ = _1228_ & ~_1261_;
	assign _1263_ = _1262_ | _1260_;
	assign _1264_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [30] ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [22];
	assign _1265_ = _1264_ ^ _1263_;
	assign _1266_ = _1265_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [6];
	assign _1267_ = _1266_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [14];
	assign _1268_ = ~(_1267_ ^ _1257_);
	assign \mchip.matrix_calculator.mul_logic.add_out2 [6] = ~(_1268_ ^ _1254_);
	assign _1269_ = _1267_ & _1257_;
	assign _1270_ = _1254_ & ~_1268_;
	assign _1271_ = ~(_1270_ | _1269_);
	assign _1272_ = ~(_1265_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [6]);
	assign _1273_ = _1266_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [14];
	assign _1274_ = _1272_ & ~_1273_;
	assign _1275_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [30] & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [22];
	assign _1276_ = _1264_ & _1263_;
	assign _1277_ = _1276_ | _1275_;
	assign _1278_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [31] ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [23];
	assign _1279_ = _1278_ ^ _1277_;
	assign _1280_ = _1279_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [7];
	assign _1281_ = _1280_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [15];
	assign _1282_ = _1281_ ^ _1274_;
	assign \mchip.matrix_calculator.mul_logic.add_out2 [7] = _1282_ ^ _1271_;
	assign _1283_ = _1274_ | ~_1281_;
	assign _1284_ = _1269_ & ~_1282_;
	assign _1285_ = _1283_ & ~_1284_;
	assign _1286_ = _1282_ | _1268_;
	assign _1287_ = _1253_ & ~_1286_;
	assign _1288_ = _1285_ & ~_1287_;
	assign _1289_ = _1286_ | _1249_;
	assign _1290_ = _1219_ & ~_1289_;
	assign _1291_ = _1290_ | ~_1288_;
	assign _1292_ = ~(_1279_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [7]);
	assign _1293_ = ~(_1280_ & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [15]);
	assign _1294_ = ~(_1293_ & _1292_);
	assign _1295_ = ~(_1278_ & _1264_);
	assign _1296_ = _1295_ | _1261_;
	assign _1297_ = _1296_ | ~_1228_;
	assign _1298_ = _1260_ & ~_1295_;
	assign _1299_ = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [31] & \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [23];
	assign _1300_ = _1278_ & _1275_;
	assign _1301_ = _1300_ | _1299_;
	assign _1302_ = _1301_ | _1298_;
	assign _1303_ = _1297_ & ~_1302_;
	assign _1304_ = _1303_ ^ _1294_;
	assign \mchip.matrix_calculator.mul_logic.add_out2 [8] = ~(_1304_ ^ _1291_);
	assign _1305_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [53];
	assign _1306_ = \mchip.matrix_calculator.shift_register.Q [61] & ~_1815_;
	assign _1307_ = _1305_ & ~_1306_;
	assign _1308_ = _1307_ | _0042_;
	assign _1309_ = _0454_ & ~_1308_;
	assign _1310_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [77];
	assign _1311_ = \mchip.matrix_calculator.shift_register.Q [93] & ~_0445_;
	assign _1312_ = _1310_ & ~_1311_;
	assign _1313_ = \mchip.matrix_calculator.shift_register.Q [125] & ~_0440_;
	assign _1314_ = \mchip.matrix_calculator.shift_register.Q [109] & ~_0442_;
	assign _1315_ = _1314_ | _1313_;
	assign _1316_ = _1312_ & ~_1315_;
	assign _1317_ = _1316_ | _0453_;
	assign _1318_ = _1317_ | _0458_;
	assign \mchip.matrix_calculator.mul_logic.mult1.S [1] = ~(_1318_ ^ _1309_);
	assign _1319_ = _1309_ & ~_1318_;
	assign _1320_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [54];
	assign _1321_ = \mchip.matrix_calculator.shift_register.Q [62] & ~_1815_;
	assign _1322_ = _1320_ & ~_1321_;
	assign _1323_ = _1322_ | _0042_;
	assign _1324_ = _1323_ | ~_0454_;
	assign _1325_ = ~(_1317_ | _1308_);
	assign _1326_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [78];
	assign _1327_ = \mchip.matrix_calculator.shift_register.Q [94] & ~_0445_;
	assign _1328_ = _1326_ & ~_1327_;
	assign _1329_ = \mchip.matrix_calculator.shift_register.Q [126] & ~_0440_;
	assign _1330_ = \mchip.matrix_calculator.shift_register.Q [110] & ~_0442_;
	assign _1331_ = _1330_ | _1329_;
	assign _1332_ = _1328_ & ~_1331_;
	assign _1333_ = _1332_ | _0453_;
	assign _1334_ = _1333_ | _0458_;
	assign _1335_ = _1334_ ^ _1325_;
	assign _1336_ = _1335_ ^ _1324_;
	assign \mchip.matrix_calculator.mul_logic.mult1.S [2] = _1336_ ^ _1319_;
	assign _1337_ = _1336_ & _1319_;
	assign _1338_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [55];
	assign _1339_ = \mchip.matrix_calculator.shift_register.Q [63] & ~_1815_;
	assign _1340_ = _1338_ & ~_1339_;
	assign _1341_ = _1340_ | _0042_;
	assign _1342_ = _0454_ & ~_1341_;
	assign _1343_ = _1335_ | _1324_;
	assign _1344_ = _1325_ & ~_1334_;
	assign _1345_ = _1343_ & ~_1344_;
	assign _1346_ = ~(_1323_ | _1317_);
	assign _1347_ = ~(_1333_ | _1308_);
	assign _1348_ = _0447_ | ~\mchip.matrix_calculator.shift_register.Q [79];
	assign _1349_ = \mchip.matrix_calculator.shift_register.Q [95] & ~_0445_;
	assign _1350_ = _1348_ & ~_1349_;
	assign _1351_ = \mchip.matrix_calculator.shift_register.Q [127] & ~_0440_;
	assign _1352_ = \mchip.matrix_calculator.shift_register.Q [111] & ~_0442_;
	assign _1353_ = _1352_ | _1351_;
	assign _1354_ = _1350_ & ~_1353_;
	assign _1355_ = _1354_ | _0453_;
	assign _1356_ = _1355_ | _0458_;
	assign _1357_ = _1356_ ^ _1347_;
	assign _1358_ = _1357_ ^ _1346_;
	assign _1359_ = ~(_1358_ ^ _1345_);
	assign _1360_ = _1359_ ^ _1342_;
	assign \mchip.matrix_calculator.mul_logic.mult1.S [3] = ~(_1360_ ^ _1337_);
	assign _1361_ = _1337_ & ~_1360_;
	assign _1362_ = ~(_1358_ | _1345_);
	assign _1363_ = _1342_ & ~_1359_;
	assign _1364_ = _1363_ | _1362_;
	assign _1365_ = ~(_1341_ | _1317_);
	assign _1366_ = _1357_ | ~_1346_;
	assign _1367_ = _1347_ & ~_1356_;
	assign _1368_ = _1367_ | ~_1366_;
	assign _1369_ = _1333_ | _1323_;
	assign _1370_ = ~(_1355_ | _1308_);
	assign _1371_ = _1370_ ^ _1369_;
	assign _1372_ = _1371_ ^ _1368_;
	assign _1373_ = ~(_1372_ ^ _1365_);
	assign _1374_ = ~(_1373_ ^ _1364_);
	assign \mchip.matrix_calculator.mul_logic.mult1.S [4] = ~(_1374_ ^ _1361_);
	assign _1375_ = _1373_ & _1364_;
	assign _1376_ = _1361_ & ~_1374_;
	assign _1377_ = ~(_1376_ | _1375_);
	assign _1378_ = _1365_ & ~_1372_;
	assign _1379_ = _1368_ & ~_1371_;
	assign _1380_ = _1379_ | _1378_;
	assign _1381_ = ~(_1341_ | _1333_);
	assign _1382_ = _1369_ | ~_1370_;
	assign _1383_ = ~(_1355_ | _1323_);
	assign _1384_ = _1383_ ^ _1382_;
	assign _1385_ = ~(_1384_ ^ _1381_);
	assign _1386_ = ~(_1385_ ^ _1380_);
	assign \mchip.matrix_calculator.mul_logic.mult1.S [5] = _1386_ ^ _1377_;
	assign _1387_ = _1385_ & _1380_;
	assign _1388_ = _1375_ & ~_1386_;
	assign _1389_ = _1388_ | _1387_;
	assign _1390_ = _1386_ | _1374_;
	assign _1391_ = _1361_ & ~_1390_;
	assign _1392_ = _1391_ | _1389_;
	assign _1393_ = _1381_ & ~_1384_;
	assign _1394_ = _1383_ & ~_1382_;
	assign _1395_ = _1394_ | _1393_;
	assign _1396_ = ~(_1355_ | _1341_);
	assign _1397_ = _1396_ ^ _1395_;
	assign \mchip.matrix_calculator.mul_logic.mult1.S [6] = _1397_ ^ _1392_;
	assign \mchip.matrix_calculator.mul_logic.add_out2 [0] = _0893_ ^ \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [8];
	assign _1398_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [49];
	assign _1399_ = \mchip.matrix_calculator.shift_register.Q [57] & ~_1815_;
	assign _1400_ = _1398_ & ~_1399_;
	assign _1401_ = _1400_ | _0042_;
	assign _1402_ = _0454_ & ~_1401_;
	assign _1403_ = _1317_ | _0754_;
	assign \mchip.matrix_calculator.mul_logic.mult5.S [1] = ~(_1403_ ^ _1402_);
	assign _1404_ = _1402_ & ~_1403_;
	assign _1405_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [50];
	assign _1406_ = \mchip.matrix_calculator.shift_register.Q [58] & ~_1815_;
	assign _1407_ = _1405_ & ~_1406_;
	assign _1408_ = _1407_ | _0042_;
	assign _1409_ = _1408_ | ~_0454_;
	assign _1410_ = ~(_1401_ | _1317_);
	assign _1411_ = _1333_ | _0754_;
	assign _1412_ = _1411_ ^ _1410_;
	assign _1413_ = _1412_ ^ _1409_;
	assign \mchip.matrix_calculator.mul_logic.mult5.S [2] = _1413_ ^ _1404_;
	assign _1414_ = _1413_ & _1404_;
	assign _1415_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [51];
	assign _1416_ = \mchip.matrix_calculator.shift_register.Q [59] & ~_1815_;
	assign _1417_ = _1415_ & ~_1416_;
	assign _1418_ = _1417_ | _0042_;
	assign _1419_ = _0454_ & ~_1418_;
	assign _1420_ = _1412_ | _1409_;
	assign _1421_ = _1410_ & ~_1411_;
	assign _1422_ = _1420_ & ~_1421_;
	assign _1423_ = ~(_1408_ | _1317_);
	assign _1424_ = ~(_1401_ | _1333_);
	assign _1425_ = _1355_ | _0754_;
	assign _1426_ = _1425_ ^ _1424_;
	assign _1427_ = _1426_ ^ _1423_;
	assign _1428_ = ~(_1427_ ^ _1422_);
	assign _1429_ = _1428_ ^ _1419_;
	assign \mchip.matrix_calculator.mul_logic.mult5.S [3] = ~(_1429_ ^ _1414_);
	assign _1430_ = _1414_ & ~_1429_;
	assign _1431_ = ~(_1427_ | _1422_);
	assign _1432_ = _1419_ & ~_1428_;
	assign _1433_ = _1432_ | _1431_;
	assign _1434_ = ~(_1418_ | _1317_);
	assign _1435_ = _1426_ | ~_1423_;
	assign _1436_ = _1424_ & ~_1425_;
	assign _1437_ = _1436_ | ~_1435_;
	assign _1438_ = _1408_ | _1333_;
	assign _1439_ = ~(_1401_ | _1355_);
	assign _1440_ = _1439_ ^ _1438_;
	assign _1441_ = _1440_ ^ _1437_;
	assign _1442_ = ~(_1441_ ^ _1434_);
	assign _1443_ = ~(_1442_ ^ _1433_);
	assign \mchip.matrix_calculator.mul_logic.mult5.S [4] = ~(_1443_ ^ _1430_);
	assign _1444_ = _1442_ & _1433_;
	assign _1445_ = _1430_ & ~_1443_;
	assign _1446_ = ~(_1445_ | _1444_);
	assign _1447_ = _1434_ & ~_1441_;
	assign _1448_ = _1437_ & ~_1440_;
	assign _1449_ = _1448_ | _1447_;
	assign _1450_ = ~(_1418_ | _1333_);
	assign _1451_ = _1438_ | ~_1439_;
	assign _1452_ = ~(_1408_ | _1355_);
	assign _1453_ = _1452_ ^ _1451_;
	assign _1454_ = ~(_1453_ ^ _1450_);
	assign _1455_ = ~(_1454_ ^ _1449_);
	assign \mchip.matrix_calculator.mul_logic.mult5.S [5] = _1455_ ^ _1446_;
	assign _1456_ = _1454_ & _1449_;
	assign _1457_ = _1444_ & ~_1455_;
	assign _1458_ = _1457_ | _1456_;
	assign _1459_ = _1455_ | _1443_;
	assign _1460_ = _1430_ & ~_1459_;
	assign _1461_ = _1460_ | _1458_;
	assign _1462_ = _1450_ & ~_1453_;
	assign _1463_ = _1452_ & ~_1451_;
	assign _1464_ = _1463_ | _1462_;
	assign _1465_ = ~(_1418_ | _1355_);
	assign _1466_ = _1465_ ^ _1464_;
	assign \mchip.matrix_calculator.mul_logic.mult5.S [6] = _1466_ ^ _1461_;
	assign _1467_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [5];
	assign _1468_ = \mchip.matrix_calculator.shift_register.Q [13] & ~_1815_;
	assign _1469_ = _1467_ & ~_1468_;
	assign _1470_ = _1469_ | _0042_;
	assign _1471_ = _0742_ & ~_1470_;
	assign _1472_ = _1105_ | _0758_;
	assign \mchip.matrix_calculator.mul_logic.mult4.S [1] = ~(_1472_ ^ _1471_);
	assign _1473_ = _1471_ & ~_1472_;
	assign _1474_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [6];
	assign _1475_ = \mchip.matrix_calculator.shift_register.Q [14] & ~_1815_;
	assign _1476_ = _1474_ & ~_1475_;
	assign _1477_ = _1476_ | _0042_;
	assign _1478_ = _1477_ | ~_0742_;
	assign _1479_ = ~(_1470_ | _1105_);
	assign _1480_ = _1121_ | _0758_;
	assign _1481_ = _1480_ ^ _1479_;
	assign _1482_ = ~(_1481_ ^ _1478_);
	assign \mchip.matrix_calculator.mul_logic.mult4.S [2] = ~(_1482_ ^ _1473_);
	assign _1483_ = _1473_ & ~_1482_;
	assign _1484_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [7];
	assign _1485_ = \mchip.matrix_calculator.shift_register.Q [15] & ~_1815_;
	assign _1486_ = _1484_ & ~_1485_;
	assign _1487_ = _1486_ | _0042_;
	assign _1488_ = _0742_ & ~_1487_;
	assign _1489_ = _1481_ | _1478_;
	assign _1490_ = _1479_ & ~_1480_;
	assign _1491_ = _1489_ & ~_1490_;
	assign _1492_ = ~(_1477_ | _1105_);
	assign _1493_ = ~(_1470_ | _1121_);
	assign _1494_ = _1137_ | _0758_;
	assign _1495_ = _1494_ ^ _1493_;
	assign _1496_ = _1495_ ^ _1492_;
	assign _1497_ = ~(_1496_ ^ _1491_);
	assign _1498_ = _1497_ ^ _1488_;
	assign \mchip.matrix_calculator.mul_logic.mult4.S [3] = ~(_1498_ ^ _1483_);
	assign _1499_ = _1483_ & ~_1498_;
	assign _1500_ = ~(_1496_ | _1491_);
	assign _1501_ = _1488_ & ~_1497_;
	assign _1502_ = _1501_ | _1500_;
	assign _1503_ = ~(_1487_ | _1105_);
	assign _1504_ = _1495_ | ~_1492_;
	assign _1505_ = _1493_ & ~_1494_;
	assign _1506_ = _1505_ | ~_1504_;
	assign _1507_ = _1477_ | _1121_;
	assign _1508_ = ~(_1470_ | _1137_);
	assign _1509_ = _1508_ ^ _1507_;
	assign _1510_ = _1509_ ^ _1506_;
	assign _1511_ = ~(_1510_ ^ _1503_);
	assign _1512_ = ~(_1511_ ^ _1502_);
	assign \mchip.matrix_calculator.mul_logic.mult4.S [4] = ~(_1512_ ^ _1499_);
	assign _1513_ = _1511_ & _1502_;
	assign _1514_ = _1499_ & ~_1512_;
	assign _1515_ = ~(_1514_ | _1513_);
	assign _1516_ = _1503_ & ~_1510_;
	assign _1517_ = _1506_ & ~_1509_;
	assign _1518_ = _1517_ | _1516_;
	assign _1519_ = ~(_1487_ | _1121_);
	assign _1520_ = _1507_ | ~_1508_;
	assign _1521_ = ~(_1477_ | _1137_);
	assign _1522_ = _1521_ ^ _1520_;
	assign _1523_ = ~(_1522_ ^ _1519_);
	assign _1524_ = ~(_1523_ ^ _1518_);
	assign \mchip.matrix_calculator.mul_logic.mult4.S [5] = _1524_ ^ _1515_;
	assign _1525_ = _1523_ & _1518_;
	assign _1526_ = _1513_ & ~_1524_;
	assign _1527_ = _1526_ | _1525_;
	assign _1528_ = _1524_ | _1512_;
	assign _1529_ = _1499_ & ~_1528_;
	assign _1530_ = _1529_ | _1527_;
	assign _1531_ = _1519_ & ~_1522_;
	assign _1532_ = _1521_ & ~_1520_;
	assign _1533_ = _1532_ | _1531_;
	assign _1534_ = ~(_1487_ | _1137_);
	assign _1535_ = _1534_ ^ _1533_;
	assign \mchip.matrix_calculator.mul_logic.mult4.S [6] = _1535_ ^ _1530_;
	assign _1536_ = ~(_0913_ | _0734_);
	assign _1537_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [17];
	assign _1538_ = \mchip.matrix_calculator.shift_register.Q [25] & ~_1815_;
	assign _1539_ = _1537_ & ~_1538_;
	assign _1540_ = _1539_ | _0042_;
	assign _1541_ = _1540_ | ~_0730_;
	assign \mchip.matrix_calculator.mul_logic.mult7.S [1] = ~(_1541_ ^ _1536_);
	assign _1542_ = _1536_ & ~_1541_;
	assign _1543_ = _0929_ | _0734_;
	assign _1544_ = ~(_1540_ | _0913_);
	assign _1545_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [18];
	assign _1546_ = \mchip.matrix_calculator.shift_register.Q [26] & ~_1815_;
	assign _1547_ = _1545_ & ~_1546_;
	assign _1548_ = _1547_ | _0042_;
	assign _1549_ = _0730_ & ~_1548_;
	assign _1550_ = _1549_ ^ _1544_;
	assign _1551_ = _1550_ ^ _1543_;
	assign \mchip.matrix_calculator.mul_logic.mult7.S [2] = ~(_1551_ ^ _1542_);
	assign _1552_ = _1542_ & ~_1551_;
	assign _1553_ = _1550_ & ~_1543_;
	assign _1554_ = ~(_0951_ | _0734_);
	assign _1555_ = _1549_ & _1544_;
	assign _1556_ = ~(_1540_ | _0929_);
	assign _1557_ = ~(_1548_ | _0913_);
	assign _1558_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [19];
	assign _1559_ = \mchip.matrix_calculator.shift_register.Q [27] & ~_1815_;
	assign _1560_ = _1558_ & ~_1559_;
	assign _1561_ = _1560_ | _0042_;
	assign _1562_ = _1561_ | ~_0730_;
	assign _1563_ = _1562_ ^ _1557_;
	assign _1564_ = _1563_ ^ _1556_;
	assign _1565_ = _1564_ ^ _1555_;
	assign _1566_ = _1565_ ^ _1554_;
	assign _1567_ = _1566_ ^ _1553_;
	assign \mchip.matrix_calculator.mul_logic.mult7.S [3] = ~(_1567_ ^ _1552_);
	assign _1568_ = _1552_ & ~_1567_;
	assign _1569_ = _1553_ & ~_1566_;
	assign _1570_ = _1569_ | _1568_;
	assign _1571_ = _1554_ & ~_1565_;
	assign _1572_ = _1555_ & ~_1564_;
	assign _1573_ = _1572_ | _1571_;
	assign _1574_ = _1563_ | ~_1556_;
	assign _1575_ = _1557_ & ~_1562_;
	assign _1576_ = _1574_ & ~_1575_;
	assign _1577_ = ~(_1540_ | _0951_);
	assign _1578_ = _1548_ | _0929_;
	assign _1579_ = _1561_ | _0913_;
	assign _1580_ = ~(_1579_ ^ _1578_);
	assign _1581_ = _1580_ ^ _1577_;
	assign _1582_ = _1581_ ^ _1576_;
	assign _1583_ = ~(_1582_ ^ _1573_);
	assign \mchip.matrix_calculator.mul_logic.mult7.S [4] = ~(_1583_ ^ _1570_);
	assign _1584_ = _1582_ & _1573_;
	assign _1585_ = _1570_ & ~_1583_;
	assign _1586_ = ~(_1585_ | _1584_);
	assign _1587_ = ~(_1581_ | _1576_);
	assign _1588_ = _1579_ | _1578_;
	assign _1589_ = _1577_ & ~_1580_;
	assign _1590_ = _1588_ & ~_1589_;
	assign _1591_ = _1548_ | _0951_;
	assign _1592_ = _1561_ | _0929_;
	assign _1593_ = ~(_1592_ ^ _1591_);
	assign _1594_ = _1593_ ^ _1590_;
	assign _1595_ = ~(_1594_ ^ _1587_);
	assign \mchip.matrix_calculator.mul_logic.mult7.S [5] = _1595_ ^ _1586_;
	assign _1596_ = _1594_ & _1587_;
	assign _1597_ = _1584_ & ~_1595_;
	assign _1598_ = _1597_ | _1596_;
	assign _1599_ = _1595_ | _1583_;
	assign _1600_ = _1570_ & ~_1599_;
	assign _1601_ = _1600_ | _1598_;
	assign _1602_ = _1593_ | _1590_;
	assign _1603_ = _1592_ | _1591_;
	assign _1604_ = ~(_1561_ | _0951_);
	assign _1605_ = ~(_1604_ ^ _1603_);
	assign _1606_ = ~(_1605_ ^ _1602_);
	assign \mchip.matrix_calculator.mul_logic.mult7.S [6] = _1606_ ^ _1601_;
	assign _1607_ = _1603_ | ~_1604_;
	assign _1608_ = _1602_ | ~_1605_;
	assign _1609_ = _1606_ & _1601_;
	assign _1610_ = _1608_ & ~_1609_;
	assign \mchip.matrix_calculator.mul_logic.mult7.S [7] = _1610_ ^ _1607_;
	assign _1611_ = ~(_1001_ | _0722_);
	assign _1612_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [37];
	assign _1613_ = \mchip.matrix_calculator.shift_register.Q [45] & ~_1815_;
	assign _1614_ = _1612_ & ~_1613_;
	assign _1615_ = _1614_ | _0042_;
	assign _1616_ = _1615_ | ~_0718_;
	assign \mchip.matrix_calculator.mul_logic.mult2.S [1] = ~(_1616_ ^ _1611_);
	assign _1617_ = _1611_ & ~_1616_;
	assign _1618_ = _1021_ | _0722_;
	assign _1619_ = ~(_1615_ | _1001_);
	assign _1620_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [38];
	assign _1621_ = \mchip.matrix_calculator.shift_register.Q [46] & ~_1815_;
	assign _1622_ = _1620_ & ~_1621_;
	assign _1623_ = _1622_ | _0042_;
	assign _1624_ = _1623_ | ~_0718_;
	assign _1625_ = _1624_ ^ _1619_;
	assign _1626_ = ~(_1625_ ^ _1618_);
	assign \mchip.matrix_calculator.mul_logic.mult2.S [2] = ~(_1626_ ^ _1617_);
	assign _1627_ = _1617_ & ~_1626_;
	assign _1628_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [39];
	assign _1629_ = \mchip.matrix_calculator.shift_register.Q [47] & ~_1815_;
	assign _1630_ = _1628_ & ~_1629_;
	assign _1631_ = _1630_ | _0042_;
	assign _1632_ = _0718_ & ~_1631_;
	assign _1633_ = _1625_ | _1618_;
	assign _1634_ = _1619_ & ~_1624_;
	assign _1635_ = _1633_ & ~_1634_;
	assign _1636_ = ~(_1037_ | _0722_);
	assign _1637_ = ~(_1615_ | _1021_);
	assign _1638_ = _1623_ | _1001_;
	assign _1639_ = _1638_ ^ _1637_;
	assign _1640_ = _1639_ ^ _1636_;
	assign _1641_ = ~(_1640_ ^ _1635_);
	assign _1642_ = _1641_ ^ _1632_;
	assign \mchip.matrix_calculator.mul_logic.mult2.S [3] = ~(_1642_ ^ _1627_);
	assign _1643_ = _1627_ & ~_1642_;
	assign _1644_ = ~(_1640_ | _1635_);
	assign _1645_ = _1632_ & ~_1641_;
	assign _1646_ = _1645_ | _1644_;
	assign _1647_ = ~(_1631_ | _1001_);
	assign _1648_ = _1639_ | ~_1636_;
	assign _1649_ = _1637_ & ~_1638_;
	assign _1650_ = _1649_ | ~_1648_;
	assign _1651_ = _1615_ | _1037_;
	assign _1652_ = ~(_1623_ | _1021_);
	assign _1653_ = _1652_ ^ _1651_;
	assign _1654_ = _1653_ ^ _1650_;
	assign _1655_ = ~(_1654_ ^ _1647_);
	assign _1656_ = ~(_1655_ ^ _1646_);
	assign \mchip.matrix_calculator.mul_logic.mult2.S [4] = ~(_1656_ ^ _1643_);
	assign _1657_ = _1655_ & _1646_;
	assign _1658_ = _1643_ & ~_1656_;
	assign _1659_ = ~(_1658_ | _1657_);
	assign _1660_ = _1647_ & ~_1654_;
	assign _1661_ = _1650_ & ~_1653_;
	assign _1662_ = _1661_ | _1660_;
	assign _1663_ = ~(_1631_ | _1021_);
	assign _1664_ = _1651_ | ~_1652_;
	assign _1665_ = ~(_1623_ | _1037_);
	assign _1666_ = _1665_ ^ _1664_;
	assign _1667_ = ~(_1666_ ^ _1663_);
	assign _1668_ = ~(_1667_ ^ _1662_);
	assign \mchip.matrix_calculator.mul_logic.mult2.S [5] = _1668_ ^ _1659_;
	assign _1669_ = _1667_ & _1662_;
	assign _1670_ = _1657_ & ~_1668_;
	assign _1671_ = _1670_ | _1669_;
	assign _1672_ = _1668_ | _1656_;
	assign _1673_ = _1643_ & ~_1672_;
	assign _1674_ = _1673_ | _1671_;
	assign _1675_ = _1663_ & ~_1666_;
	assign _1676_ = _1665_ & ~_1664_;
	assign _1677_ = _1676_ | _1675_;
	assign _1678_ = ~(_1631_ | _1037_);
	assign _1679_ = _1678_ ^ _1677_;
	assign \mchip.matrix_calculator.mul_logic.mult2.S [6] = _1679_ ^ _1674_;
	assign _1680_ = _0992_ & _0991_;
	assign _1681_ = _0993_ & _0988_;
	assign \mchip.matrix_calculator.mul_logic.mult3.S [7] = _1681_ | _1680_;
	assign _1682_ = _0877_ & ~_0890_;
	assign _1683_ = _0880_ & ~_0889_;
	assign \mchip.matrix_calculator.mul_logic.add_out [9] = _1683_ | _1682_;
	assign _1684_ = _1185_ & _1184_;
	assign _1685_ = _1186_ & _1181_;
	assign \mchip.matrix_calculator.mul_logic.mult8.S [7] = _1685_ | _1684_;
	assign _1686_ = _1291_ & ~_1304_;
	assign _1687_ = _1294_ & ~_1303_;
	assign \mchip.matrix_calculator.mul_logic.add_out2 [9] = _1687_ | _1686_;
	assign _1688_ = _1396_ & _1395_;
	assign _1689_ = _1397_ & _1392_;
	assign \mchip.matrix_calculator.mul_logic.mult1.S [7] = _1689_ | _1688_;
	assign _1690_ = _1465_ & _1464_;
	assign _1691_ = _1466_ & _1461_;
	assign \mchip.matrix_calculator.mul_logic.mult5.S [7] = _1691_ | _1690_;
	assign _1692_ = _1534_ & _1533_;
	assign _1693_ = _1535_ & _1530_;
	assign \mchip.matrix_calculator.mul_logic.mult4.S [7] = _1693_ | _1692_;
	assign _1694_ = _1678_ & _1677_;
	assign _1695_ = _1679_ & _1674_;
	assign \mchip.matrix_calculator.mul_logic.mult2.S [7] = _1695_ | _1694_;
	assign _1696_ = \mchip.matrix_calculator.shift_register.Q [0] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1];
	assign _1697_ = \mchip.matrix_calculator.shift_register.Q [8] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _1698_ = ~(_1697_ | _1696_);
	assign _1699_ = \mchip.matrix_calculator.shift_register.Q [24] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _1700_ = \mchip.matrix_calculator.shift_register.Q [16] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _1701_ = _1700_ | _1699_;
	assign _1702_ = _1698_ & ~_1701_;
	assign _1703_ = \mchip.matrix_calculator.shift_register.Q [56] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _1704_ = \mchip.matrix_calculator.shift_register.Q [48] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _1705_ = _1704_ | _1703_;
	assign _1706_ = \mchip.matrix_calculator.shift_register.Q [40] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _1707_ = \mchip.matrix_calculator.shift_register.Q [32] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _1708_ = _1707_ | _1706_;
	assign _1709_ = _1708_ | _1705_;
	assign _1710_ = _1702_ & ~_1709_;
	assign _1711_ = ~(\mchip.matrix_calculator.add_logic.fsm.cur_state [9] | \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _1712_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [7] | \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _1713_ = _1711_ & ~_1712_;
	assign _1714_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [5] | \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _1715_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [8] | \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _1716_ = _1715_ | _1714_;
	assign _1717_ = _1713_ & ~_1716_;
	assign _1718_ = ~_1717_;
	assign _1719_ = _1718_ & ~_1710_;
	assign _1720_ = ~(\mchip.matrix_calculator.add_logic.fsm.cur_state [9] & \mchip.matrix_calculator.shift_register.Q [72]);
	assign _1721_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [1] & \mchip.matrix_calculator.shift_register.Q [64];
	assign _1722_ = _1720_ & ~_1721_;
	assign _1723_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [7] & \mchip.matrix_calculator.shift_register.Q [88];
	assign _1724_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [4] & \mchip.matrix_calculator.shift_register.Q [80];
	assign _1725_ = _1724_ | _1723_;
	assign _1726_ = _1722_ & ~_1725_;
	assign _1727_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [5] & \mchip.matrix_calculator.shift_register.Q [120];
	assign _1728_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [3] & \mchip.matrix_calculator.shift_register.Q [112];
	assign _1729_ = _1728_ | _1727_;
	assign _1730_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [8] & \mchip.matrix_calculator.shift_register.Q [104];
	assign _1731_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [2] & \mchip.matrix_calculator.shift_register.Q [96];
	assign _1732_ = _1731_ | _1730_;
	assign _1733_ = _1732_ | _1729_;
	assign _1734_ = _1726_ & ~_1733_;
	assign _1735_ = _1718_ & ~_1734_;
	assign \mchip.matrix_calculator.add_logic.add2.S [0] = _1735_ ^ _1719_;
	assign _1736_ = ~(\mchip.matrix_calculator.shift_register.Q [4] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _1737_ = \mchip.matrix_calculator.shift_register.Q [12] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _1738_ = _1736_ & ~_1737_;
	assign _1739_ = \mchip.matrix_calculator.shift_register.Q [28] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _1740_ = \mchip.matrix_calculator.shift_register.Q [20] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _1741_ = _1740_ | _1739_;
	assign _1742_ = _1738_ & ~_1741_;
	assign _1743_ = \mchip.matrix_calculator.shift_register.Q [60] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _1744_ = \mchip.matrix_calculator.shift_register.Q [52] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _1745_ = _1744_ | _1743_;
	assign _1746_ = \mchip.matrix_calculator.shift_register.Q [44] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _1747_ = \mchip.matrix_calculator.shift_register.Q [36] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _1748_ = _1747_ | _1746_;
	assign _1749_ = _1748_ | _1745_;
	assign _1750_ = _1742_ & ~_1749_;
	assign _1751_ = _1718_ & ~_1750_;
	assign _1752_ = ~(\mchip.matrix_calculator.shift_register.Q [68] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _1753_ = \mchip.matrix_calculator.shift_register.Q [76] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _1754_ = _1752_ & ~_1753_;
	assign _1755_ = \mchip.matrix_calculator.shift_register.Q [92] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _1756_ = \mchip.matrix_calculator.shift_register.Q [84] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _1757_ = _1756_ | _1755_;
	assign _1758_ = _1754_ & ~_1757_;
	assign _1759_ = \mchip.matrix_calculator.shift_register.Q [124] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _1760_ = \mchip.matrix_calculator.shift_register.Q [116] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _1761_ = _1760_ | _1759_;
	assign _1762_ = \mchip.matrix_calculator.shift_register.Q [108] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _1763_ = \mchip.matrix_calculator.shift_register.Q [100] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _1764_ = _1763_ | _1762_;
	assign _1765_ = _1764_ | _1761_;
	assign _1766_ = _1758_ & ~_1765_;
	assign _1767_ = _1718_ & ~_1766_;
	assign \mchip.matrix_calculator.add_logic.add1.S [0] = _1767_ ^ _1751_;
	assign _1768_ = \mchip.matrix_calculator.op_reg.Q [1] | \mchip.matrix_calculator.op_reg.Q [0];
	assign _1769_ = \mchip.matrix_calculator.fsm.cur_state [1] & ~_1768_;
	assign _1770_ = _1769_ | \mchip.sync13.sync ;
	assign _1771_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [0] & ~_1770_;
	assign _0041_ = _1771_ | \mchip.sync13.sync ;
	assign _1772_ = \mchip.sync9.sync  & ~\mchip.matrix_calculator.ed_de.tmp1 ;
	assign _1773_ = _1772_ | \mchip.sync13.sync ;
	assign _1774_ = \mchip.matrix_calculator.fsm.cur_state [20] & ~_1773_;
	assign _1775_ = ~\mchip.sync13.sync ;
	assign _1776_ = ~(_1772_ & _1775_);
	assign _1777_ = \mchip.matrix_calculator.fsm.cur_state [10] & ~_1776_;
	assign _0032_ = _1777_ | _1774_;
	assign _1778_ = \mchip.matrix_calculator.fsm.cur_state [19] & ~_1773_;
	assign _1779_ = \mchip.matrix_calculator.fsm.cur_state [9] & ~_1776_;
	assign _0031_ = _1779_ | _1778_;
	assign _1780_ = \mchip.matrix_calculator.fsm.cur_state [18] & ~_1773_;
	assign _1781_ = \mchip.matrix_calculator.fsm.cur_state [8] & ~_1776_;
	assign _0030_ = _1781_ | _1780_;
	assign _1782_ = \mchip.sync13.sync  | ~\mchip.matrix_calculator.add_logic.fsm.cur_state [6];
	assign _1783_ = \mchip.matrix_calculator.fsm.cur_state [7] & ~_1782_;
	assign _1784_ = \mchip.sync13.sync  | ~\mchip.matrix_calculator.mul_logic.fsm.cur_state [4];
	assign _1785_ = \mchip.matrix_calculator.fsm.cur_state [12] & ~_1784_;
	assign _1786_ = \mchip.matrix_calculator.fsm.cur_state [17] & ~\mchip.sync13.sync ;
	assign _1787_ = _1786_ | _1785_;
	assign _0029_ = _1787_ | _1783_;
	assign _1788_ = \mchip.matrix_calculator.fsm.cur_state [16] & ~_1773_;
	assign _1789_ = \mchip.matrix_calculator.fsm.cur_state [6] & ~_1776_;
	assign _0028_ = _1789_ | _1788_;
	assign _1790_ = \mchip.matrix_calculator.fsm.cur_state [15] & ~_1773_;
	assign _1791_ = \mchip.matrix_calculator.fsm.cur_state [5] & ~_1776_;
	assign _0027_ = _1791_ | _1790_;
	assign _1792_ = \mchip.matrix_calculator.fsm.cur_state [0] & ~_1773_;
	assign _0021_ = _1792_ | \mchip.sync13.sync ;
	assign _1793_ = \mchip.matrix_calculator.fsm.cur_state [11] & ~_1773_;
	assign _1794_ = \mchip.matrix_calculator.fsm.cur_state [0] & ~_1776_;
	assign _0023_ = _1794_ | _1793_;
	assign _1795_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [4] | \mchip.sync13.sync ;
	assign _1796_ = \mchip.matrix_calculator.fsm.cur_state [12] & ~_1795_;
	assign _1797_ = _1768_ | \mchip.sync13.sync ;
	assign _1798_ = \mchip.matrix_calculator.fsm.cur_state [1] & ~_1797_;
	assign _0024_ = _1798_ | _1796_;
	assign _1799_ = \mchip.matrix_calculator.fsm.cur_state [2] & ~_1776_;
	assign _1800_ = \mchip.matrix_calculator.fsm.cur_state [13] & ~_1773_;
	assign _0025_ = _1800_ | _1799_;
	assign _1801_ = \mchip.matrix_calculator.fsm.cur_state [3] & ~_1776_;
	assign _1802_ = \mchip.matrix_calculator.fsm.cur_state [14] & ~_1773_;
	assign _0026_ = _1802_ | _1801_;
	assign _1803_ = \mchip.matrix_calculator.fsm.cur_state [1] & \mchip.matrix_calculator.op_reg.Q [1];
	assign _1804_ = _1803_ | \mchip.sync13.sync ;
	assign _1805_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [0] & ~_1804_;
	assign _0020_ = _1805_ | \mchip.sync13.sync ;
	assign _2025_[0] = ~\mchip.matrix_calculator.index_counter.Q [0];
	assign _1806_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [9] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [10];
	assign _1807_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [7] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [8];
	assign _1808_ = _1807_ | _1806_;
	assign _1809_ = ~(\mchip.matrix_calculator.mul_logic.fsm.cur_state [2] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [1]);
	assign _1810_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [3] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [5];
	assign _1811_ = _1809_ & ~_1810_;
	assign \mchip.matrix_calculator.mul_logic.fsm.layer_2_en  = _1808_ | ~_1811_;
	assign _1812_ = \mchip.matrix_calculator.fsm.cur_state [10] & ~_1773_;
	assign _1813_ = \mchip.matrix_calculator.fsm.cur_state [15] & ~_1776_;
	assign _0022_ = _1813_ | _1812_;
	assign _1814_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [6] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [8];
	assign _1815_ = ~(_1814_ | _1806_);
	assign _0042_ = _1815_ & _1811_;
	assign _1816_ = \mchip.matrix_calculator.fsm.cur_state [9] & ~_1773_;
	assign _1817_ = \mchip.matrix_calculator.fsm.cur_state [14] & ~_1776_;
	assign _0040_ = _1817_ | _1816_;
	assign _1818_ = \mchip.matrix_calculator.fsm.cur_state [8] & ~_1773_;
	assign _1819_ = \mchip.matrix_calculator.fsm.cur_state [13] & ~_1776_;
	assign _0039_ = _1819_ | _1818_;
	assign _1820_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [6] | \mchip.sync13.sync ;
	assign _1821_ = \mchip.matrix_calculator.fsm.cur_state [7] & ~_1820_;
	assign _1822_ = \mchip.sync13.sync  | ~\mchip.matrix_calculator.op_reg.Q [1];
	assign _1823_ = \mchip.matrix_calculator.fsm.cur_state [1] & ~_1822_;
	assign _0038_ = _1823_ | _1821_;
	assign _1824_ = \mchip.matrix_calculator.fsm.cur_state [19] & ~_1776_;
	assign _1825_ = \mchip.matrix_calculator.fsm.cur_state [2] & ~_1773_;
	assign _0033_ = _1825_ | _1824_;
	assign _1826_ = \mchip.matrix_calculator.fsm.cur_state [6] & ~_1773_;
	assign _1827_ = \mchip.matrix_calculator.fsm.cur_state [11] & ~_1776_;
	assign _0037_ = _1827_ | _1826_;
	assign _1828_ = \mchip.matrix_calculator.fsm.cur_state [5] & ~_1773_;
	assign _1829_ = \mchip.matrix_calculator.fsm.cur_state [18] & ~_1776_;
	assign _0036_ = _1829_ | _1828_;
	assign _1830_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.op_reg.Q [0];
	assign _1831_ = _1830_ | \mchip.sync13.sync ;
	assign _1832_ = \mchip.matrix_calculator.fsm.cur_state [1] & ~_1831_;
	assign _1833_ = \mchip.matrix_calculator.fsm.cur_state [4] & ~\mchip.sync13.sync ;
	assign _0035_ = _1833_ | _1832_;
	assign _1834_ = \mchip.matrix_calculator.fsm.cur_state [3] & ~_1773_;
	assign _1835_ = \mchip.matrix_calculator.fsm.cur_state [16] & ~_1776_;
	assign _0034_ = _1835_ | _1834_;
	assign _1836_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [8] | \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _1837_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [5] | \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _1838_ = _1837_ | _1836_;
	assign _1839_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [3] | \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _1840_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [2] | \mchip.matrix_calculator.add_logic.fsm.cur_state [1];
	assign _1841_ = _1840_ | _1839_;
	assign \mchip.matrix_calculator.add_logic.fsm.shift_en  = _1841_ | _1838_;
	assign _1842_ = ~(\mchip.matrix_calculator.fsm.cur_state [2] | \mchip.matrix_calculator.fsm.cur_state [0]);
	assign _1843_ = \mchip.matrix_calculator.fsm.cur_state [3] | \mchip.matrix_calculator.fsm.cur_state [5];
	assign _1844_ = _1842_ & ~_1843_;
	assign _1845_ = \mchip.matrix_calculator.fsm.cur_state [9] | \mchip.matrix_calculator.fsm.cur_state [10];
	assign _1846_ = \mchip.matrix_calculator.fsm.cur_state [6] | \mchip.matrix_calculator.fsm.cur_state [8];
	assign _1847_ = _1846_ | _1845_;
	assign _1848_ = _1844_ & ~_1847_;
	assign _1849_ = \mchip.matrix_calculator.fsm.cur_state [19] | \mchip.matrix_calculator.fsm.cur_state [20];
	assign _1850_ = \mchip.matrix_calculator.fsm.cur_state [16] | \mchip.matrix_calculator.fsm.cur_state [18];
	assign _1851_ = _1850_ | _1849_;
	assign _1852_ = \mchip.matrix_calculator.fsm.cur_state [14] | \mchip.matrix_calculator.fsm.cur_state [15];
	assign _1853_ = \mchip.matrix_calculator.fsm.cur_state [13] | \mchip.matrix_calculator.fsm.cur_state [11];
	assign _1854_ = _1853_ | _1852_;
	assign _1855_ = _1854_ | _1851_;
	assign _1856_ = _1848_ & ~_1855_;
	assign \mchip.matrix_calculator.op_reg.en  = _1772_ & ~_1856_;
	assign _1857_ = \mchip.matrix_calculator.fsm.cur_state [12] & \mchip.matrix_calculator.mul_logic.fsm.cur_state [4];
	assign _1858_ = \mchip.matrix_calculator.fsm.cur_state [7] & \mchip.matrix_calculator.add_logic.fsm.cur_state [6];
	assign _1859_ = _1858_ | \mchip.matrix_calculator.fsm.cur_state [17];
	assign _1860_ = _1859_ | _1857_;
	assign _1861_ = ~(\mchip.matrix_calculator.fsm.cur_state [7] | \mchip.matrix_calculator.fsm.cur_state [17]);
	assign _1862_ = _1861_ & ~\mchip.matrix_calculator.fsm.cur_state [12];
	assign \mchip.finish  = _1860_ & ~_1862_;
	assign _1863_ = \mchip.matrix_calculator.sw_de.tmp1  | ~\mchip.sync10.sync ;
	assign \mchip.matrix_calculator.index_counter.en  = \mchip.finish  & ~_1863_;
	assign _1864_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [150] : \mchip.matrix_calculator.mul_logic.shift_register.Q [150]);
	assign _1865_ = ~\mchip.matrix_calculator.index_counter.Q [4];
	assign _1866_ = \mchip.matrix_calculator.index_counter.Q [2] | \mchip.matrix_calculator.index_counter.Q [3];
	assign _1867_ = \mchip.matrix_calculator.index_counter.Q [1] | ~\mchip.matrix_calculator.index_counter.Q [0];
	assign _1868_ = _1867_ | _1866_;
	assign _1869_ = _1865_ & ~_1868_;
	assign _1870_ = _1869_ & _1864_;
	assign _1871_ = \mchip.matrix_calculator.index_counter.Q [0] | ~\mchip.matrix_calculator.index_counter.Q [1];
	assign _1872_ = _1871_ | _1866_;
	assign _1873_ = _1865_ & ~_1872_;
	assign _1874_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [145];
	assign _1875_ = _1873_ & ~_1874_;
	assign _1876_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [140] : \mchip.matrix_calculator.mul_logic.shift_register.Q [140]);
	assign _1877_ = \mchip.matrix_calculator.index_counter.Q [1] & \mchip.matrix_calculator.index_counter.Q [0];
	assign _1878_ = _1866_ | ~_1877_;
	assign _1879_ = _1865_ & ~_1878_;
	assign _1880_ = _1879_ & _1876_;
	assign _1881_ = _1880_ | _1875_;
	assign _1882_ = _1881_ | _1870_;
	assign _1883_ = \mchip.matrix_calculator.index_counter.Q [3] | ~\mchip.matrix_calculator.index_counter.Q [2];
	assign _1884_ = \mchip.matrix_calculator.index_counter.Q [1] | \mchip.matrix_calculator.index_counter.Q [0];
	assign _1885_ = _1884_ | _1883_;
	assign _1886_ = _1865_ & ~_1885_;
	assign _1887_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [135];
	assign _1888_ = _1886_ & ~_1887_;
	assign _1889_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [130] : \mchip.matrix_calculator.mul_logic.shift_register.Q [130]);
	assign _1890_ = _1883_ | _1867_;
	assign _1891_ = _1865_ & ~_1890_;
	assign _1892_ = _1891_ & _1889_;
	assign _1893_ = _1892_ | _1888_;
	assign _1894_ = _1883_ | _1871_;
	assign _1895_ = _1865_ & ~_1894_;
	assign _1896_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [125];
	assign _1897_ = _1895_ & ~_1896_;
	assign _1898_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [120] : \mchip.matrix_calculator.mul_logic.shift_register.Q [120]);
	assign _1899_ = _1883_ | ~_1877_;
	assign _1900_ = _1865_ & ~_1899_;
	assign _1901_ = _1900_ & _1898_;
	assign _1902_ = _1901_ | _1897_;
	assign _1903_ = _1902_ | _1893_;
	assign _1904_ = _1903_ | _1882_;
	assign _1905_ = \mchip.matrix_calculator.index_counter.Q [2] | ~\mchip.matrix_calculator.index_counter.Q [3];
	assign _1906_ = _1905_ | _1884_;
	assign _1907_ = _1865_ & ~_1906_;
	assign _1908_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [115];
	assign _1909_ = _1907_ & ~_1908_;
	assign _1910_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [110] : \mchip.matrix_calculator.mul_logic.shift_register.Q [110]);
	assign _1911_ = _1905_ | _1867_;
	assign _1912_ = _1865_ & ~_1911_;
	assign _1913_ = _1912_ & _1910_;
	assign _1914_ = _1913_ | _1909_;
	assign _1915_ = _1905_ | _1871_;
	assign _1916_ = _1865_ & ~_1915_;
	assign _1917_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [105];
	assign _1918_ = _1916_ & ~_1917_;
	assign _1919_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [100] : \mchip.matrix_calculator.mul_logic.shift_register.Q [100]);
	assign _1920_ = _1905_ | ~_1877_;
	assign _1921_ = _1865_ & ~_1920_;
	assign _1922_ = _1921_ & _1919_;
	assign _1923_ = _1922_ | _1918_;
	assign _1924_ = _1923_ | _1914_;
	assign _1925_ = ~(\mchip.matrix_calculator.index_counter.Q [2] & \mchip.matrix_calculator.index_counter.Q [3]);
	assign _1926_ = _1925_ | _1884_;
	assign _1927_ = _1865_ & ~_1926_;
	assign _1928_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [95];
	assign _1929_ = _1927_ & ~_1928_;
	assign _1930_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [90] : \mchip.matrix_calculator.mul_logic.shift_register.Q [90]);
	assign _1931_ = _1925_ | _1867_;
	assign _1932_ = _1865_ & ~_1931_;
	assign _1933_ = _1932_ & _1930_;
	assign _1934_ = _1933_ | _1929_;
	assign _1935_ = _1925_ | _1871_;
	assign _1936_ = _1865_ & ~_1935_;
	assign _1937_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [85];
	assign _1938_ = _1936_ & ~_1937_;
	assign _1939_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [80] : \mchip.matrix_calculator.mul_logic.shift_register.Q [80]);
	assign _1940_ = _1925_ | ~_1877_;
	assign _1941_ = _1865_ & ~_1940_;
	assign _1942_ = _1941_ & _1939_;
	assign _1943_ = _1942_ | _1938_;
	assign _1944_ = _1943_ | _1934_;
	assign _1945_ = _1944_ | _1924_;
	assign _1946_ = _1945_ | _1904_;
	assign _1947_ = _1884_ | _1866_;
	assign _1948_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1947_;
	assign _1949_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [75];
	assign _1950_ = _1948_ & ~_1949_;
	assign _1951_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [70] : \mchip.matrix_calculator.mul_logic.shift_register.Q [70]);
	assign _1952_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1868_;
	assign _1953_ = _1952_ & _1951_;
	assign _1954_ = _1953_ | _1950_;
	assign _1955_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1872_;
	assign _1956_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [65];
	assign _1957_ = _1955_ & ~_1956_;
	assign _1958_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [60] : \mchip.matrix_calculator.mul_logic.shift_register.Q [60]);
	assign _1959_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1878_;
	assign _1960_ = _1959_ & _1958_;
	assign _1961_ = _1960_ | _1957_;
	assign _1962_ = _1961_ | _1954_;
	assign _1963_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1885_;
	assign _1964_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [55];
	assign _1965_ = _1963_ & ~_1964_;
	assign _1966_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [50] : \mchip.matrix_calculator.mul_logic.shift_register.Q [50]);
	assign _1967_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1890_;
	assign _1968_ = _1967_ & _1966_;
	assign _1969_ = _1968_ | _1965_;
	assign _1970_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1894_;
	assign _1971_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [45];
	assign _1972_ = _1970_ & ~_1971_;
	assign _1973_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [40] : \mchip.matrix_calculator.mul_logic.shift_register.Q [40]);
	assign _1974_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1899_;
	assign _1975_ = _1974_ & _1973_;
	assign _1976_ = _1975_ | _1972_;
	assign _1977_ = _1976_ | _1969_;
	assign _1978_ = _1977_ | _1962_;
	assign _1979_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1906_;
	assign _1980_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [35];
	assign _1981_ = _1979_ & ~_1980_;
	assign _1982_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [30] : \mchip.matrix_calculator.mul_logic.shift_register.Q [30]);
	assign _1983_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1911_;
	assign _1984_ = _1983_ & _1982_;
	assign _1985_ = _1984_ | _1981_;
	assign _1986_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1915_;
	assign _1987_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [25];
	assign _1988_ = _1986_ & ~_1987_;
	assign _1989_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [20] : \mchip.matrix_calculator.mul_logic.shift_register.Q [20]);
	assign _1990_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1920_;
	assign _1991_ = _1990_ & _1989_;
	assign _1992_ = _1991_ | _1988_;
	assign _1993_ = _1992_ | _1985_;
	assign _1994_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1926_;
	assign _1995_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [15];
	assign _1996_ = _1994_ & ~_1995_;
	assign _1997_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [10] : \mchip.matrix_calculator.mul_logic.shift_register.Q [10]);
	assign _1998_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1931_;
	assign _1999_ = _1998_ & _1997_;
	assign _2000_ = _1999_ | _1996_;
	assign _2001_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1935_;
	assign _2002_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [5];
	assign _2003_ = _2001_ & ~_2002_;
	assign _2004_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [0] : \mchip.matrix_calculator.mul_logic.shift_register.Q [0]);
	assign _2005_ = \mchip.matrix_calculator.index_counter.Q [4] & ~_1940_;
	assign _2006_ = _2005_ & _2004_;
	assign _2007_ = _2006_ | _2003_;
	assign _2008_ = _2007_ | _2000_;
	assign _2009_ = _2008_ | _1993_;
	assign _2010_ = _2009_ | _1978_;
	assign _2011_ = _2010_ | _1946_;
	assign _2012_ = _2005_ | _2001_;
	assign _2013_ = _1998_ | _1994_;
	assign _2014_ = _2013_ | _2012_;
	assign _2015_ = _1983_ | _1979_;
	assign _2016_ = _1990_ | _1986_;
	assign _2017_ = _2016_ | _2015_;
	assign _2018_ = _2017_ | _2014_;
	assign _2019_ = _1952_ | _1948_;
	assign _2020_ = _1959_ | _1955_;
	assign _2021_ = _2020_ | _2019_;
	assign _2022_ = _1967_ | _1963_;
	assign _2023_ = _1974_ | _1970_;
	assign _2024_ = _2023_ | _2022_;
	assign _0043_ = _2024_ | _2021_;
	assign _0044_ = _0043_ | _2018_;
	assign _0045_ = _1879_ | _1873_;
	assign _0046_ = _0045_ | _1869_;
	assign _0047_ = _1891_ | _1886_;
	assign _0048_ = _1900_ | _1895_;
	assign _0049_ = _0048_ | _0047_;
	assign _0050_ = _0049_ | _0046_;
	assign _0051_ = _1912_ | _1907_;
	assign _0052_ = _1921_ | _1916_;
	assign _0053_ = _0052_ | _0051_;
	assign _0054_ = _1932_ | _1927_;
	assign _0055_ = _1941_ | _1936_;
	assign _0056_ = _0055_ | _0054_;
	assign _0057_ = _0056_ | _0053_;
	assign _0058_ = _0057_ | _0050_;
	assign _0059_ = _0058_ | _0044_;
	assign _0060_ = \mchip.matrix_calculator.mul_logic.shift_register.Q [155] & ~\mchip.matrix_calculator.op_reg.Q [1];
	assign io_out[0] = (_0059_ ? _2011_ : _0060_);
	assign _0061_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [151] : \mchip.matrix_calculator.mul_logic.shift_register.Q [151]);
	assign _0062_ = _0061_ & _1869_;
	assign _0063_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [146];
	assign _0064_ = _1873_ & ~_0063_;
	assign _0065_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [141] : \mchip.matrix_calculator.mul_logic.shift_register.Q [141]);
	assign _0066_ = _0065_ & _1879_;
	assign _0067_ = _0066_ | _0064_;
	assign _0068_ = _0067_ | _0062_;
	assign _0069_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [136];
	assign _0070_ = _1886_ & ~_0069_;
	assign _0071_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [131] : \mchip.matrix_calculator.mul_logic.shift_register.Q [131]);
	assign _0072_ = _0071_ & _1891_;
	assign _0073_ = _0072_ | _0070_;
	assign _0074_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [126];
	assign _0075_ = _1895_ & ~_0074_;
	assign _0076_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [121] : \mchip.matrix_calculator.mul_logic.shift_register.Q [121]);
	assign _0077_ = _0076_ & _1900_;
	assign _0078_ = _0077_ | _0075_;
	assign _0079_ = _0078_ | _0073_;
	assign _0080_ = _0079_ | _0068_;
	assign _0081_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [116];
	assign _0082_ = _1907_ & ~_0081_;
	assign _0083_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [111] : \mchip.matrix_calculator.mul_logic.shift_register.Q [111]);
	assign _0084_ = _0083_ & _1912_;
	assign _0085_ = _0084_ | _0082_;
	assign _0086_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [106];
	assign _0087_ = _1916_ & ~_0086_;
	assign _0088_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [101] : \mchip.matrix_calculator.mul_logic.shift_register.Q [101]);
	assign _0089_ = _0088_ & _1921_;
	assign _0090_ = _0089_ | _0087_;
	assign _0091_ = _0090_ | _0085_;
	assign _0092_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [96];
	assign _0093_ = _1927_ & ~_0092_;
	assign _0094_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [91] : \mchip.matrix_calculator.mul_logic.shift_register.Q [91]);
	assign _0095_ = _0094_ & _1932_;
	assign _0096_ = _0095_ | _0093_;
	assign _0097_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [86];
	assign _0098_ = _1936_ & ~_0097_;
	assign _0099_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [81] : \mchip.matrix_calculator.mul_logic.shift_register.Q [81]);
	assign _0100_ = _0099_ & _1941_;
	assign _0101_ = _0100_ | _0098_;
	assign _0102_ = _0101_ | _0096_;
	assign _0103_ = _0102_ | _0091_;
	assign _0104_ = _0103_ | _0080_;
	assign _0105_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [76];
	assign _0106_ = _1948_ & ~_0105_;
	assign _0107_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [71] : \mchip.matrix_calculator.mul_logic.shift_register.Q [71]);
	assign _0108_ = _0107_ & _1952_;
	assign _0109_ = _0108_ | _0106_;
	assign _0110_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [66];
	assign _0111_ = _1955_ & ~_0110_;
	assign _0112_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [61] : \mchip.matrix_calculator.mul_logic.shift_register.Q [61]);
	assign _0113_ = _0112_ & _1959_;
	assign _0114_ = _0113_ | _0111_;
	assign _0115_ = _0114_ | _0109_;
	assign _0116_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [56];
	assign _0117_ = _1963_ & ~_0116_;
	assign _0118_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [51] : \mchip.matrix_calculator.mul_logic.shift_register.Q [51]);
	assign _0119_ = _0118_ & _1967_;
	assign _0120_ = _0119_ | _0117_;
	assign _0121_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [46];
	assign _0122_ = _1970_ & ~_0121_;
	assign _0123_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [41] : \mchip.matrix_calculator.mul_logic.shift_register.Q [41]);
	assign _0124_ = _0123_ & _1974_;
	assign _0125_ = _0124_ | _0122_;
	assign _0126_ = _0125_ | _0120_;
	assign _0127_ = _0126_ | _0115_;
	assign _0128_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [36];
	assign _0129_ = _1979_ & ~_0128_;
	assign _0130_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [31] : \mchip.matrix_calculator.mul_logic.shift_register.Q [31]);
	assign _0131_ = _0130_ & _1983_;
	assign _0132_ = _0131_ | _0129_;
	assign _0133_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [26];
	assign _0134_ = _1986_ & ~_0133_;
	assign _0135_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [21] : \mchip.matrix_calculator.mul_logic.shift_register.Q [21]);
	assign _0136_ = _0135_ & _1990_;
	assign _0137_ = _0136_ | _0134_;
	assign _0138_ = _0137_ | _0132_;
	assign _0139_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [16];
	assign _0140_ = _1994_ & ~_0139_;
	assign _0141_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [11] : \mchip.matrix_calculator.mul_logic.shift_register.Q [11]);
	assign _0142_ = _0141_ & _1998_;
	assign _0143_ = _0142_ | _0140_;
	assign _0144_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [6];
	assign _0145_ = _2001_ & ~_0144_;
	assign _0146_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [1] : \mchip.matrix_calculator.mul_logic.shift_register.Q [1]);
	assign _0147_ = _0146_ & _2005_;
	assign _0148_ = _0147_ | _0145_;
	assign _0149_ = _0148_ | _0143_;
	assign _0150_ = _0149_ | _0138_;
	assign _0151_ = _0150_ | _0127_;
	assign _0152_ = _0151_ | _0104_;
	assign _0153_ = \mchip.matrix_calculator.mul_logic.shift_register.Q [156] & ~\mchip.matrix_calculator.op_reg.Q [1];
	assign io_out[1] = (_0059_ ? _0152_ : _0153_);
	assign _0154_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [152] : \mchip.matrix_calculator.mul_logic.shift_register.Q [152]);
	assign _0155_ = _0154_ & _1869_;
	assign _0156_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [147];
	assign _0157_ = _1873_ & ~_0156_;
	assign _0158_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [142] : \mchip.matrix_calculator.mul_logic.shift_register.Q [142]);
	assign _0159_ = _0158_ & _1879_;
	assign _0160_ = _0159_ | _0157_;
	assign _0161_ = _0160_ | _0155_;
	assign _0162_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [137];
	assign _0163_ = _1886_ & ~_0162_;
	assign _0164_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [132] : \mchip.matrix_calculator.mul_logic.shift_register.Q [132]);
	assign _0165_ = _0164_ & _1891_;
	assign _0166_ = _0165_ | _0163_;
	assign _0167_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [127];
	assign _0168_ = _1895_ & ~_0167_;
	assign _0169_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [122] : \mchip.matrix_calculator.mul_logic.shift_register.Q [122]);
	assign _0170_ = _0169_ & _1900_;
	assign _0171_ = _0170_ | _0168_;
	assign _0172_ = _0171_ | _0166_;
	assign _0173_ = _0172_ | _0161_;
	assign _0174_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [117];
	assign _0175_ = _1907_ & ~_0174_;
	assign _0176_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [112] : \mchip.matrix_calculator.mul_logic.shift_register.Q [112]);
	assign _0177_ = _0176_ & _1912_;
	assign _0178_ = _0177_ | _0175_;
	assign _0179_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [107];
	assign _0180_ = _1916_ & ~_0179_;
	assign _0181_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [102] : \mchip.matrix_calculator.mul_logic.shift_register.Q [102]);
	assign _0182_ = _0181_ & _1921_;
	assign _0183_ = _0182_ | _0180_;
	assign _0184_ = _0183_ | _0178_;
	assign _0185_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [97];
	assign _0186_ = _1927_ & ~_0185_;
	assign _0187_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [92] : \mchip.matrix_calculator.mul_logic.shift_register.Q [92]);
	assign _0188_ = _0187_ & _1932_;
	assign _0189_ = _0188_ | _0186_;
	assign _0190_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [87];
	assign _0191_ = _1936_ & ~_0190_;
	assign _0192_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [82] : \mchip.matrix_calculator.mul_logic.shift_register.Q [82]);
	assign _0193_ = _0192_ & _1941_;
	assign _0194_ = _0193_ | _0191_;
	assign _0195_ = _0194_ | _0189_;
	assign _0196_ = _0195_ | _0184_;
	assign _0197_ = _0196_ | _0173_;
	assign _0198_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [77];
	assign _0199_ = _1948_ & ~_0198_;
	assign _0200_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [72] : \mchip.matrix_calculator.mul_logic.shift_register.Q [72]);
	assign _0201_ = _0200_ & _1952_;
	assign _0202_ = _0201_ | _0199_;
	assign _0203_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [67];
	assign _0204_ = _1955_ & ~_0203_;
	assign _0205_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [62] : \mchip.matrix_calculator.mul_logic.shift_register.Q [62]);
	assign _0206_ = _0205_ & _1959_;
	assign _0207_ = _0206_ | _0204_;
	assign _0208_ = _0207_ | _0202_;
	assign _0209_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [57];
	assign _0210_ = _1963_ & ~_0209_;
	assign _0211_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [52] : \mchip.matrix_calculator.mul_logic.shift_register.Q [52]);
	assign _0212_ = _0211_ & _1967_;
	assign _0213_ = _0212_ | _0210_;
	assign _0214_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [47];
	assign _0215_ = _1970_ & ~_0214_;
	assign _0216_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [42] : \mchip.matrix_calculator.mul_logic.shift_register.Q [42]);
	assign _0217_ = _0216_ & _1974_;
	assign _0218_ = _0217_ | _0215_;
	assign _0219_ = _0218_ | _0213_;
	assign _0220_ = _0219_ | _0208_;
	assign _0221_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [37];
	assign _0222_ = _1979_ & ~_0221_;
	assign _0223_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [32] : \mchip.matrix_calculator.mul_logic.shift_register.Q [32]);
	assign _0224_ = _0223_ & _1983_;
	assign _0225_ = _0224_ | _0222_;
	assign _0226_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [27];
	assign _0227_ = _1986_ & ~_0226_;
	assign _0228_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [22] : \mchip.matrix_calculator.mul_logic.shift_register.Q [22]);
	assign _0229_ = _0228_ & _1990_;
	assign _0230_ = _0229_ | _0227_;
	assign _0231_ = _0230_ | _0225_;
	assign _0232_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [17];
	assign _0233_ = _1994_ & ~_0232_;
	assign _0234_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [12] : \mchip.matrix_calculator.mul_logic.shift_register.Q [12]);
	assign _0235_ = _0234_ & _1998_;
	assign _0236_ = _0235_ | _0233_;
	assign _0237_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [7];
	assign _0238_ = _2001_ & ~_0237_;
	assign _0239_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [2] : \mchip.matrix_calculator.mul_logic.shift_register.Q [2]);
	assign _0240_ = _0239_ & _2005_;
	assign _0241_ = _0240_ | _0238_;
	assign _0242_ = _0241_ | _0236_;
	assign _0243_ = _0242_ | _0231_;
	assign _0244_ = _0243_ | _0220_;
	assign _0245_ = _0244_ | _0197_;
	assign _0246_ = \mchip.matrix_calculator.mul_logic.shift_register.Q [157] & ~\mchip.matrix_calculator.op_reg.Q [1];
	assign io_out[2] = (_0059_ ? _0245_ : _0246_);
	assign _0247_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [153] : \mchip.matrix_calculator.mul_logic.shift_register.Q [153]);
	assign _0248_ = _0247_ & _1869_;
	assign _0249_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [148];
	assign _0250_ = _1873_ & ~_0249_;
	assign _0251_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [143] : \mchip.matrix_calculator.mul_logic.shift_register.Q [143]);
	assign _0252_ = _0251_ & _1879_;
	assign _0253_ = _0252_ | _0250_;
	assign _0254_ = _0253_ | _0248_;
	assign _0255_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [138];
	assign _0256_ = _1886_ & ~_0255_;
	assign _0257_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [133] : \mchip.matrix_calculator.mul_logic.shift_register.Q [133]);
	assign _0258_ = _0257_ & _1891_;
	assign _0259_ = _0258_ | _0256_;
	assign _0260_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [128];
	assign _0261_ = _1895_ & ~_0260_;
	assign _0262_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [123] : \mchip.matrix_calculator.mul_logic.shift_register.Q [123]);
	assign _0263_ = _0262_ & _1900_;
	assign _0264_ = _0263_ | _0261_;
	assign _0265_ = _0264_ | _0259_;
	assign _0266_ = _0265_ | _0254_;
	assign _0267_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [118];
	assign _0268_ = _1907_ & ~_0267_;
	assign _0269_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [113] : \mchip.matrix_calculator.mul_logic.shift_register.Q [113]);
	assign _0270_ = _0269_ & _1912_;
	assign _0271_ = _0270_ | _0268_;
	assign _0272_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [108];
	assign _0273_ = _1916_ & ~_0272_;
	assign _0274_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [103] : \mchip.matrix_calculator.mul_logic.shift_register.Q [103]);
	assign _0275_ = _0274_ & _1921_;
	assign _0276_ = _0275_ | _0273_;
	assign _0277_ = _0276_ | _0271_;
	assign _0278_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [98];
	assign _0279_ = _1927_ & ~_0278_;
	assign _0280_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [93] : \mchip.matrix_calculator.mul_logic.shift_register.Q [93]);
	assign _0281_ = _0280_ & _1932_;
	assign _0282_ = _0281_ | _0279_;
	assign _0283_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [88];
	assign _0284_ = _1936_ & ~_0283_;
	assign _0285_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [83] : \mchip.matrix_calculator.mul_logic.shift_register.Q [83]);
	assign _0286_ = _0285_ & _1941_;
	assign _0287_ = _0286_ | _0284_;
	assign _0288_ = _0287_ | _0282_;
	assign _0289_ = _0288_ | _0277_;
	assign _0290_ = _0289_ | _0266_;
	assign _0291_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [78];
	assign _0292_ = _1948_ & ~_0291_;
	assign _0293_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [73] : \mchip.matrix_calculator.mul_logic.shift_register.Q [73]);
	assign _0294_ = _0293_ & _1952_;
	assign _0295_ = _0294_ | _0292_;
	assign _0296_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [68];
	assign _0297_ = _1955_ & ~_0296_;
	assign _0298_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [63] : \mchip.matrix_calculator.mul_logic.shift_register.Q [63]);
	assign _0299_ = _0298_ & _1959_;
	assign _0300_ = _0299_ | _0297_;
	assign _0301_ = _0300_ | _0295_;
	assign _0302_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [58];
	assign _0303_ = _1963_ & ~_0302_;
	assign _0304_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [53] : \mchip.matrix_calculator.mul_logic.shift_register.Q [53]);
	assign _0305_ = _0304_ & _1967_;
	assign _0306_ = _0305_ | _0303_;
	assign _0307_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [48];
	assign _0308_ = _1970_ & ~_0307_;
	assign _0309_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [43] : \mchip.matrix_calculator.mul_logic.shift_register.Q [43]);
	assign _0310_ = _0309_ & _1974_;
	assign _0311_ = _0310_ | _0308_;
	assign _0312_ = _0311_ | _0306_;
	assign _0313_ = _0312_ | _0301_;
	assign _0314_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [38];
	assign _0315_ = _1979_ & ~_0314_;
	assign _0316_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [33] : \mchip.matrix_calculator.mul_logic.shift_register.Q [33]);
	assign _0317_ = _0316_ & _1983_;
	assign _0318_ = _0317_ | _0315_;
	assign _0319_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [28];
	assign _0320_ = _1986_ & ~_0319_;
	assign _0321_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [23] : \mchip.matrix_calculator.mul_logic.shift_register.Q [23]);
	assign _0322_ = _0321_ & _1990_;
	assign _0323_ = _0322_ | _0320_;
	assign _0324_ = _0323_ | _0318_;
	assign _0325_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [18];
	assign _0326_ = _1994_ & ~_0325_;
	assign _0327_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [13] : \mchip.matrix_calculator.mul_logic.shift_register.Q [13]);
	assign _0328_ = _0327_ & _1998_;
	assign _0329_ = _0328_ | _0326_;
	assign _0330_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [8];
	assign _0331_ = _2001_ & ~_0330_;
	assign _0332_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [3] : \mchip.matrix_calculator.mul_logic.shift_register.Q [3]);
	assign _0333_ = _0332_ & _2005_;
	assign _0334_ = _0333_ | _0331_;
	assign _0335_ = _0334_ | _0329_;
	assign _0336_ = _0335_ | _0324_;
	assign _0337_ = _0336_ | _0313_;
	assign _0338_ = _0337_ | _0290_;
	assign _0339_ = \mchip.matrix_calculator.mul_logic.shift_register.Q [158] & ~\mchip.matrix_calculator.op_reg.Q [1];
	assign io_out[3] = (_0059_ ? _0338_ : _0339_);
	assign _0340_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [154] : \mchip.matrix_calculator.mul_logic.shift_register.Q [154]);
	assign _0341_ = _0340_ & _1869_;
	assign _0342_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [149];
	assign _0343_ = _1873_ & ~_0342_;
	assign _0344_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [144] : \mchip.matrix_calculator.mul_logic.shift_register.Q [144]);
	assign _0345_ = _0344_ & _1879_;
	assign _0346_ = _0345_ | _0343_;
	assign _0347_ = _0346_ | _0341_;
	assign _0348_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [139];
	assign _0349_ = _1886_ & ~_0348_;
	assign _0350_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [134] : \mchip.matrix_calculator.mul_logic.shift_register.Q [134]);
	assign _0351_ = _0350_ & _1891_;
	assign _0352_ = _0351_ | _0349_;
	assign _0353_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [129];
	assign _0354_ = _1895_ & ~_0353_;
	assign _0355_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [124] : \mchip.matrix_calculator.mul_logic.shift_register.Q [124]);
	assign _0356_ = _0355_ & _1900_;
	assign _0357_ = _0356_ | _0354_;
	assign _0358_ = _0357_ | _0352_;
	assign _0359_ = _0358_ | _0347_;
	assign _0360_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [119];
	assign _0361_ = _1907_ & ~_0360_;
	assign _0362_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [114] : \mchip.matrix_calculator.mul_logic.shift_register.Q [114]);
	assign _0363_ = _0362_ & _1912_;
	assign _0364_ = _0363_ | _0361_;
	assign _0365_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [109];
	assign _0366_ = _1916_ & ~_0365_;
	assign _0367_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [104] : \mchip.matrix_calculator.mul_logic.shift_register.Q [104]);
	assign _0368_ = _0367_ & _1921_;
	assign _0369_ = _0368_ | _0366_;
	assign _0370_ = _0369_ | _0364_;
	assign _0371_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [99];
	assign _0372_ = _1927_ & ~_0371_;
	assign _0373_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [94] : \mchip.matrix_calculator.mul_logic.shift_register.Q [94]);
	assign _0374_ = _0373_ & _1932_;
	assign _0375_ = _0374_ | _0372_;
	assign _0376_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [89];
	assign _0377_ = _1936_ & ~_0376_;
	assign _0378_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [84] : \mchip.matrix_calculator.mul_logic.shift_register.Q [84]);
	assign _0379_ = _0378_ & _1941_;
	assign _0380_ = _0379_ | _0377_;
	assign _0381_ = _0380_ | _0375_;
	assign _0382_ = _0381_ | _0370_;
	assign _0383_ = _0382_ | _0359_;
	assign _0384_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [79];
	assign _0385_ = _1948_ & ~_0384_;
	assign _0386_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [74] : \mchip.matrix_calculator.mul_logic.shift_register.Q [74]);
	assign _0387_ = _0386_ & _1952_;
	assign _0388_ = _0387_ | _0385_;
	assign _0389_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [69];
	assign _0390_ = _1955_ & ~_0389_;
	assign _0391_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [64] : \mchip.matrix_calculator.mul_logic.shift_register.Q [64]);
	assign _0392_ = _0391_ & _1959_;
	assign _0393_ = _0392_ | _0390_;
	assign _0394_ = _0393_ | _0388_;
	assign _0395_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [59];
	assign _0396_ = _1963_ & ~_0395_;
	assign _0397_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [54] : \mchip.matrix_calculator.mul_logic.shift_register.Q [54]);
	assign _0398_ = _0397_ & _1967_;
	assign _0399_ = _0398_ | _0396_;
	assign _0400_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [49];
	assign _0401_ = _1970_ & ~_0400_;
	assign _0402_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [44] : \mchip.matrix_calculator.mul_logic.shift_register.Q [44]);
	assign _0403_ = _0402_ & _1974_;
	assign _0404_ = _0403_ | _0401_;
	assign _0405_ = _0404_ | _0399_;
	assign _0406_ = _0405_ | _0394_;
	assign _0407_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [39];
	assign _0408_ = _1979_ & ~_0407_;
	assign _0409_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [34] : \mchip.matrix_calculator.mul_logic.shift_register.Q [34]);
	assign _0410_ = _0409_ & _1983_;
	assign _0411_ = _0410_ | _0408_;
	assign _0412_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [29];
	assign _0413_ = _1986_ & ~_0412_;
	assign _0414_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [24] : \mchip.matrix_calculator.mul_logic.shift_register.Q [24]);
	assign _0415_ = _0414_ & _1990_;
	assign _0416_ = _0415_ | _0413_;
	assign _0417_ = _0416_ | _0411_;
	assign _0418_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [19];
	assign _0419_ = _1994_ & ~_0418_;
	assign _0420_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [14] : \mchip.matrix_calculator.mul_logic.shift_register.Q [14]);
	assign _0421_ = _0420_ & _1998_;
	assign _0422_ = _0421_ | _0419_;
	assign _0423_ = \mchip.matrix_calculator.op_reg.Q [1] | ~\mchip.matrix_calculator.mul_logic.shift_register.Q [9];
	assign _0424_ = _2001_ & ~_0423_;
	assign _0425_ = (\mchip.matrix_calculator.op_reg.Q [1] ? \mchip.matrix_calculator.add_logic.shift1.Q [4] : \mchip.matrix_calculator.mul_logic.shift_register.Q [4]);
	assign _0426_ = _0425_ & _2005_;
	assign _0427_ = _0426_ | _0424_;
	assign _0428_ = _0427_ | _0422_;
	assign _0429_ = _0428_ | _0417_;
	assign _0430_ = _0429_ | _0406_;
	assign _0431_ = _0430_ | _0383_;
	assign _0432_ = \mchip.matrix_calculator.mul_logic.shift_register.Q [159] & ~\mchip.matrix_calculator.op_reg.Q [1];
	assign io_out[4] = (_0059_ ? _0431_ : _0432_);
	assign _0433_ = \mchip.matrix_calculator.fsm.cur_state [1] & ~_1830_;
	assign _0434_ = _0433_ | \mchip.matrix_calculator.fsm.cur_state [4];
	assign _0435_ = ~(\mchip.matrix_calculator.fsm.cur_state [4] | \mchip.matrix_calculator.fsm.cur_state [1]);
	assign \mchip.error  = _0434_ & ~_0435_;
	assign _0012_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [6] & ~\mchip.sync13.sync ;
	assign _0011_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [9] & ~\mchip.sync13.sync ;
	assign _0010_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [10] & ~\mchip.sync13.sync ;
	assign _0008_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [4] & ~\mchip.sync13.sync ;
	assign _0009_ = \mchip.matrix_calculator.fsm.cur_state [20] & ~_1776_;
	assign _0436_ = ~(\mchip.matrix_calculator.mul_logic.fsm.cur_state [7] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [4]);
	assign _0013_ = _1775_ & ~_0436_;
	assign _0014_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [8] & ~\mchip.sync13.sync ;
	assign _0437_ = ~(_1769_ & _1775_);
	assign _0015_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [0] & ~_0437_;
	assign _0016_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [1] & ~\mchip.sync13.sync ;
	assign _0017_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [2] & ~\mchip.sync13.sync ;
	assign _0018_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [3] & ~\mchip.sync13.sync ;
	assign _0019_ = \mchip.matrix_calculator.mul_logic.fsm.cur_state [5] & ~\mchip.sync13.sync ;
	assign _0000_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [9] & ~\mchip.sync13.sync ;
	assign _0007_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [3] & ~\mchip.sync13.sync ;
	assign _0006_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [2] & ~\mchip.sync13.sync ;
	assign _0438_ = ~(\mchip.matrix_calculator.add_logic.fsm.cur_state [6] | \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0005_ = _1775_ & ~_0438_;
	assign _0439_ = ~(_1803_ & _1775_);
	assign _0004_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [0] & ~_0439_;
	assign _0003_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [7] & ~\mchip.sync13.sync ;
	assign _0002_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [5] & ~\mchip.sync13.sync ;
	assign _0001_ = \mchip.matrix_calculator.add_logic.fsm.cur_state [8] & ~\mchip.sync13.sync ;
	assign _0440_ = ~(\mchip.matrix_calculator.mul_logic.fsm.cur_state [6] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [3]);
	assign _0441_ = \mchip.matrix_calculator.shift_register.Q [124] & ~_0440_;
	assign _0442_ = ~(\mchip.matrix_calculator.mul_logic.fsm.cur_state [9] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [2]);
	assign _0443_ = \mchip.matrix_calculator.shift_register.Q [108] & ~_0442_;
	assign _0444_ = _0443_ | _0441_;
	assign _0445_ = ~(\mchip.matrix_calculator.mul_logic.fsm.cur_state [8] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [5]);
	assign _0446_ = \mchip.matrix_calculator.shift_register.Q [92] & ~_0445_;
	assign _0447_ = ~(\mchip.matrix_calculator.mul_logic.fsm.cur_state [10] | \mchip.matrix_calculator.mul_logic.fsm.cur_state [1]);
	assign _0448_ = \mchip.matrix_calculator.shift_register.Q [76] & ~_0447_;
	assign _0449_ = _0448_ | _0446_;
	assign _0450_ = _0449_ | _0444_;
	assign _0451_ = _0447_ & _0445_;
	assign _0452_ = ~(_0442_ & _0440_);
	assign _0453_ = _0451_ & ~_0452_;
	assign _0454_ = _0450_ & ~_0453_;
	assign _0455_ = _1811_ | ~\mchip.matrix_calculator.shift_register.Q [52];
	assign _0456_ = \mchip.matrix_calculator.shift_register.Q [60] & ~_1815_;
	assign _0457_ = _0455_ & ~_0456_;
	assign _0458_ = _0457_ | _0042_;
	assign \mchip.matrix_calculator.mul_logic.mult1.S [0] = _0454_ & ~_0458_;
	assign _2026_[1] = ~(_1871_ & _1867_);
	assign _2026_[2] = _1877_ ^ \mchip.matrix_calculator.index_counter.Q [2];
	assign _0459_ = _1877_ & \mchip.matrix_calculator.index_counter.Q [2];
	assign _2026_[3] = _0459_ ^ \mchip.matrix_calculator.index_counter.Q [3];
	assign _2026_[4] = _1940_ ^ _1865_;
	assign _0460_ = _1735_ | ~_1719_;
	assign _0461_ = ~(\mchip.matrix_calculator.shift_register.Q [1] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0462_ = \mchip.matrix_calculator.shift_register.Q [9] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0463_ = _0461_ & ~_0462_;
	assign _0464_ = \mchip.matrix_calculator.shift_register.Q [25] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0465_ = \mchip.matrix_calculator.shift_register.Q [17] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0466_ = _0465_ | _0464_;
	assign _0467_ = _0463_ & ~_0466_;
	assign _0468_ = \mchip.matrix_calculator.shift_register.Q [57] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0469_ = \mchip.matrix_calculator.shift_register.Q [49] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0470_ = _0469_ | _0468_;
	assign _0471_ = \mchip.matrix_calculator.shift_register.Q [41] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0472_ = \mchip.matrix_calculator.shift_register.Q [33] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0473_ = _0472_ | _0471_;
	assign _0474_ = _0473_ | _0470_;
	assign _0475_ = _0467_ & ~_0474_;
	assign _0476_ = _1718_ & ~_0475_;
	assign _0477_ = ~_0476_;
	assign _0478_ = ~(_0476_ ^ _1719_);
	assign _0479_ = (\mchip.matrix_calculator.op_reg.Q [0] ? _0477_ : _0478_);
	assign _0480_ = ~(\mchip.matrix_calculator.shift_register.Q [65] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0481_ = \mchip.matrix_calculator.shift_register.Q [73] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0482_ = _0480_ & ~_0481_;
	assign _0483_ = \mchip.matrix_calculator.shift_register.Q [89] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0484_ = \mchip.matrix_calculator.shift_register.Q [81] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0485_ = _0484_ | _0483_;
	assign _0486_ = _0482_ & ~_0485_;
	assign _0487_ = \mchip.matrix_calculator.shift_register.Q [121] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0488_ = \mchip.matrix_calculator.shift_register.Q [113] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0489_ = _0488_ | _0487_;
	assign _0490_ = \mchip.matrix_calculator.shift_register.Q [105] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0491_ = \mchip.matrix_calculator.shift_register.Q [97] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0492_ = _0491_ | _0490_;
	assign _0493_ = _0492_ | _0489_;
	assign _0494_ = _0486_ & ~_0493_;
	assign _0495_ = _1718_ & ~_0494_;
	assign _0496_ = _0495_ ^ _0479_;
	assign \mchip.matrix_calculator.add_logic.add2.S [1] = _0496_ ^ _0460_;
	assign _0497_ = _0495_ & _0479_;
	assign _0498_ = _0496_ & _0460_;
	assign _0499_ = _0498_ | _0497_;
	assign _0500_ = ~(\mchip.matrix_calculator.shift_register.Q [2] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0501_ = \mchip.matrix_calculator.shift_register.Q [10] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0502_ = _0500_ & ~_0501_;
	assign _0503_ = \mchip.matrix_calculator.shift_register.Q [26] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0504_ = \mchip.matrix_calculator.shift_register.Q [18] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0505_ = _0504_ | _0503_;
	assign _0506_ = _0502_ & ~_0505_;
	assign _0507_ = \mchip.matrix_calculator.shift_register.Q [58] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0508_ = \mchip.matrix_calculator.shift_register.Q [50] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0509_ = _0508_ | _0507_;
	assign _0510_ = \mchip.matrix_calculator.shift_register.Q [42] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0511_ = \mchip.matrix_calculator.shift_register.Q [34] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0512_ = _0511_ | _0510_;
	assign _0513_ = _0512_ | _0509_;
	assign _0514_ = _0506_ & ~_0513_;
	assign _0515_ = _1718_ & ~_0514_;
	assign _0516_ = ~_0515_;
	assign _0517_ = ~(_0476_ | _1719_);
	assign _0518_ = _0515_ ^ _0517_;
	assign _0519_ = (\mchip.matrix_calculator.op_reg.Q [0] ? _0516_ : _0518_);
	assign _0520_ = ~(\mchip.matrix_calculator.shift_register.Q [66] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0521_ = \mchip.matrix_calculator.shift_register.Q [74] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0522_ = _0520_ & ~_0521_;
	assign _0523_ = \mchip.matrix_calculator.shift_register.Q [90] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0524_ = \mchip.matrix_calculator.shift_register.Q [82] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0525_ = _0524_ | _0523_;
	assign _0526_ = _0522_ & ~_0525_;
	assign _0527_ = \mchip.matrix_calculator.shift_register.Q [122] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0528_ = \mchip.matrix_calculator.shift_register.Q [114] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0529_ = _0528_ | _0527_;
	assign _0530_ = \mchip.matrix_calculator.shift_register.Q [106] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0531_ = \mchip.matrix_calculator.shift_register.Q [98] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0532_ = _0531_ | _0530_;
	assign _0533_ = _0532_ | _0529_;
	assign _0534_ = _0526_ & ~_0533_;
	assign _0535_ = _1718_ & ~_0534_;
	assign _0536_ = _0535_ ^ _0519_;
	assign \mchip.matrix_calculator.add_logic.add2.S [2] = _0536_ ^ _0499_;
	assign _0537_ = _0535_ & _0519_;
	assign _0538_ = _0536_ & _0499_;
	assign _0539_ = _0538_ | _0537_;
	assign _0540_ = ~(\mchip.matrix_calculator.shift_register.Q [3] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0541_ = \mchip.matrix_calculator.shift_register.Q [11] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0542_ = _0540_ & ~_0541_;
	assign _0543_ = \mchip.matrix_calculator.shift_register.Q [27] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0544_ = \mchip.matrix_calculator.shift_register.Q [19] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0545_ = _0544_ | _0543_;
	assign _0546_ = _0542_ & ~_0545_;
	assign _0547_ = \mchip.matrix_calculator.shift_register.Q [59] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0548_ = \mchip.matrix_calculator.shift_register.Q [51] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0549_ = _0548_ | _0547_;
	assign _0550_ = \mchip.matrix_calculator.shift_register.Q [43] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0551_ = \mchip.matrix_calculator.shift_register.Q [35] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0552_ = _0551_ | _0550_;
	assign _0553_ = _0552_ | _0549_;
	assign _0554_ = _0546_ & ~_0553_;
	assign _0555_ = _1718_ & ~_0554_;
	assign _0556_ = _0515_ | ~_0517_;
	assign _0557_ = _0555_ ^ _0556_;
	assign _0558_ = (\mchip.matrix_calculator.op_reg.Q [0] ? _0555_ : _0557_);
	assign _0559_ = ~(\mchip.matrix_calculator.shift_register.Q [67] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0560_ = \mchip.matrix_calculator.shift_register.Q [75] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0561_ = _0559_ & ~_0560_;
	assign _0562_ = \mchip.matrix_calculator.shift_register.Q [91] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0563_ = \mchip.matrix_calculator.shift_register.Q [83] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0564_ = _0563_ | _0562_;
	assign _0565_ = _0561_ & ~_0564_;
	assign _0566_ = \mchip.matrix_calculator.shift_register.Q [123] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0567_ = \mchip.matrix_calculator.shift_register.Q [115] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0568_ = _0567_ | _0566_;
	assign _0569_ = \mchip.matrix_calculator.shift_register.Q [107] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0570_ = \mchip.matrix_calculator.shift_register.Q [99] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0571_ = _0570_ | _0569_;
	assign _0572_ = _0571_ | _0568_;
	assign _0573_ = _0565_ & ~_0572_;
	assign _0574_ = _1718_ & ~_0573_;
	assign _0575_ = ~(_0574_ ^ _0558_);
	assign \mchip.matrix_calculator.add_logic.add2.S [3] = _0575_ ^ _0539_;
	assign _0576_ = _0558_ | ~_0574_;
	assign _0577_ = _0575_ & _0537_;
	assign _0578_ = _0576_ & ~_0577_;
	assign _0579_ = ~(_0575_ & _0536_);
	assign _0580_ = _0499_ & ~_0579_;
	assign _0581_ = _0578_ & ~_0580_;
	assign _0582_ = ~\mchip.matrix_calculator.op_reg.Q [0];
	assign _0583_ = _0555_ | _0515_;
	assign _0584_ = _0517_ & ~_0583_;
	assign _0585_ = _0582_ & ~_0584_;
	assign \mchip.matrix_calculator.add_logic.add2.S [4] = _0585_ ^ _0581_;
	assign _0586_ = _1767_ | ~_1751_;
	assign _0587_ = ~(\mchip.matrix_calculator.shift_register.Q [5] & \mchip.matrix_calculator.add_logic.fsm.cur_state [1]);
	assign _0588_ = \mchip.matrix_calculator.shift_register.Q [13] & \mchip.matrix_calculator.add_logic.fsm.cur_state [9];
	assign _0589_ = _0587_ & ~_0588_;
	assign _0590_ = \mchip.matrix_calculator.shift_register.Q [29] & \mchip.matrix_calculator.add_logic.fsm.cur_state [7];
	assign _0591_ = \mchip.matrix_calculator.shift_register.Q [21] & \mchip.matrix_calculator.add_logic.fsm.cur_state [4];
	assign _0592_ = _0591_ | _0590_;
	assign _0593_ = _0589_ & ~_0592_;
	assign _0594_ = \mchip.matrix_calculator.shift_register.Q [61] & \mchip.matrix_calculator.add_logic.fsm.cur_state [5];
	assign _0595_ = \mchip.matrix_calculator.shift_register.Q [53] & \mchip.matrix_calculator.add_logic.fsm.cur_state [3];
	assign _0596_ = _0595_ | _0594_;
	assign _0597_ = \mchip.matrix_calculator.shift_register.Q [45] & \mchip.matrix_calculator.add_logic.fsm.cur_state [8];
	assign _0598_ = \mchip.matrix_calculator.shift_register.Q [37] & \mchip.matrix_calculator.add_logic.fsm.cur_state [2];
	assign _0599_ = _0598_ | _0597_;
	assign _0600_ = _0599_ | _0596_;
	assign _0601_ = _0593_ & ~_0600_;
	assign _0602_ = _1718_ & ~_0601_;
	assign _0603_ = ~_0602_;
	assign _0604_ = ~(_0602_ ^ _1751_);
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [0] <= _0041_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [1] <= _0010_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [2] <= _0011_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [3] <= _0012_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [4] <= _0013_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [5] <= _0014_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [6] <= _0015_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [7] <= _0016_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [8] <= _0017_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [9] <= _0018_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.mul_logic.fsm.cur_state [10] <= _0019_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [0] <= _0021_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [1] <= _0009_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [2] <= _0033_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [3] <= _0034_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [4] <= _0035_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [5] <= _0036_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [6] <= _0037_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [7] <= _0038_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [8] <= _0039_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [9] <= _0040_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [10] <= _0022_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [11] <= _0023_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [12] <= _0024_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [13] <= _0025_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [14] <= _0026_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [15] <= _0027_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [16] <= _0028_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [17] <= _0029_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [18] <= _0030_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [19] <= _0031_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.fsm.cur_state [20] <= _0032_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [0] <= _0020_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [1] <= _0000_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [2] <= _0001_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [3] <= _0002_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [4] <= _0003_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [5] <= _0004_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [6] <= _0005_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [7] <= _0006_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [8] <= _0007_;
	always @(posedge io_in[12]) \mchip.matrix_calculator.add_logic.fsm.cur_state [9] <= _0008_;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[0] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[0]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[0]  <= \mchip.matrix_calculator.add_logic.add2.S [0];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [0] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[0] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[1] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[1]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[1]  <= \mchip.matrix_calculator.add_logic.add2.S [1];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [1] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[1] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[2] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[2]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[2]  <= \mchip.matrix_calculator.add_logic.add2.S [2];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [2] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[2] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[3] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[3]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[3]  <= \mchip.matrix_calculator.add_logic.add2.S [3];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [3] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[3] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[4] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[4]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[4]  <= \mchip.matrix_calculator.add_logic.add2.S [4];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [4] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[4] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[10] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[10]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[10]  <= \mchip.matrix_calculator.add_logic.add1.S [0];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [10] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[10] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[11] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[11]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[11]  <= \mchip.matrix_calculator.add_logic.add1.S [1];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [11] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[11] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[12] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[12]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[12]  <= \mchip.matrix_calculator.add_logic.add1.S [2];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [12] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[12] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[13] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[13]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[13]  <= \mchip.matrix_calculator.add_logic.add1.S [3];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [13] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[13] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[14] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[14]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[14]  <= \mchip.matrix_calculator.add_logic.add1.S [4];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [14] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[14] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[20] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[20]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[20]  <= \mchip.matrix_calculator.add_logic.shift1.Q [0];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [20] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[20] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[21] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[21]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[21]  <= \mchip.matrix_calculator.add_logic.shift1.Q [1];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [21] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[21] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[22] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[22]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[22]  <= \mchip.matrix_calculator.add_logic.shift1.Q [2];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [22] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[22] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[23] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[23]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[23]  <= \mchip.matrix_calculator.add_logic.shift1.Q [3];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [23] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[23] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[24] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[24]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[24]  <= \mchip.matrix_calculator.add_logic.shift1.Q [4];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [24] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[24] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[30] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[30]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[30]  <= \mchip.matrix_calculator.add_logic.shift1.Q [10];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [30] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[30] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[31] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[31]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[31]  <= \mchip.matrix_calculator.add_logic.shift1.Q [11];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [31] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[31] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[32] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[32]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[32]  <= \mchip.matrix_calculator.add_logic.shift1.Q [12];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [32] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[32] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[33] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[33]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[33]  <= \mchip.matrix_calculator.add_logic.shift1.Q [13];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [33] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[33] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[34] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[34]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[34]  <= \mchip.matrix_calculator.add_logic.shift1.Q [14];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [34] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[34] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[40] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[40]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[40]  <= \mchip.matrix_calculator.add_logic.shift1.Q [20];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [40] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[40] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[41] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[41]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[41]  <= \mchip.matrix_calculator.add_logic.shift1.Q [21];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [41] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[41] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[42] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[42]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[42]  <= \mchip.matrix_calculator.add_logic.shift1.Q [22];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [42] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[42] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[43] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[43]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[43]  <= \mchip.matrix_calculator.add_logic.shift1.Q [23];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [43] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[43] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[44] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[44]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[44]  <= \mchip.matrix_calculator.add_logic.shift1.Q [24];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [44] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[44] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[50] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[50]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[50]  <= \mchip.matrix_calculator.add_logic.shift1.Q [30];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [50] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[50] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[51] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[51]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[51]  <= \mchip.matrix_calculator.add_logic.shift1.Q [31];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [51] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[51] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[52] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[52]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[52]  <= \mchip.matrix_calculator.add_logic.shift1.Q [32];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [52] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[52] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[53] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[53]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[53]  <= \mchip.matrix_calculator.add_logic.shift1.Q [33];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [53] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[53] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[54] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[54]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[54]  <= \mchip.matrix_calculator.add_logic.shift1.Q [34];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [54] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[54] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[60] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[60]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[60]  <= \mchip.matrix_calculator.add_logic.shift1.Q [40];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [60] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[60] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[61] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[61]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[61]  <= \mchip.matrix_calculator.add_logic.shift1.Q [41];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [61] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[61] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[62] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[62]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[62]  <= \mchip.matrix_calculator.add_logic.shift1.Q [42];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [62] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[62] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[63] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[63]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[63]  <= \mchip.matrix_calculator.add_logic.shift1.Q [43];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [63] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[63] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[64] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[64]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[64]  <= \mchip.matrix_calculator.add_logic.shift1.Q [44];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [64] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[64] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[70] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[70]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[70]  <= \mchip.matrix_calculator.add_logic.shift1.Q [50];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [70] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[70] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[71] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[71]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[71]  <= \mchip.matrix_calculator.add_logic.shift1.Q [51];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [71] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[71] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[72] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[72]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[72]  <= \mchip.matrix_calculator.add_logic.shift1.Q [52];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [72] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[72] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[73] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[73]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[73]  <= \mchip.matrix_calculator.add_logic.shift1.Q [53];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [73] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[73] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[74] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[74]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[74]  <= \mchip.matrix_calculator.add_logic.shift1.Q [54];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [74] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[74] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[80] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[80]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[80]  <= \mchip.matrix_calculator.add_logic.shift1.Q [60];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [80] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[80] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[81] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[81]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[81]  <= \mchip.matrix_calculator.add_logic.shift1.Q [61];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [81] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[81] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[82] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[82]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[82]  <= \mchip.matrix_calculator.add_logic.shift1.Q [62];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [82] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[82] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[83] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[83]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[83]  <= \mchip.matrix_calculator.add_logic.shift1.Q [63];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [83] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[83] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[84] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[84]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[84]  <= \mchip.matrix_calculator.add_logic.shift1.Q [64];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [84] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[84] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[90] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[90]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[90]  <= \mchip.matrix_calculator.add_logic.shift1.Q [70];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [90] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[90] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[91] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[91]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[91]  <= \mchip.matrix_calculator.add_logic.shift1.Q [71];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [91] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[91] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[92] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[92]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[92]  <= \mchip.matrix_calculator.add_logic.shift1.Q [72];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [92] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[92] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[93] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[93]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[93]  <= \mchip.matrix_calculator.add_logic.shift1.Q [73];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [93] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[93] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[94] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[94]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[94]  <= \mchip.matrix_calculator.add_logic.shift1.Q [74];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [94] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[94] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[100] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[100]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[100]  <= \mchip.matrix_calculator.add_logic.shift1.Q [80];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [100] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[100] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[101] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[101]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[101]  <= \mchip.matrix_calculator.add_logic.shift1.Q [81];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [101] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[101] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[102] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[102]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[102]  <= \mchip.matrix_calculator.add_logic.shift1.Q [82];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [102] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[102] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[103] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[103]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[103]  <= \mchip.matrix_calculator.add_logic.shift1.Q [83];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [103] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[103] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[104] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[104]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[104]  <= \mchip.matrix_calculator.add_logic.shift1.Q [84];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [104] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[104] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[110] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[110]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[110]  <= \mchip.matrix_calculator.add_logic.shift1.Q [90];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [110] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[110] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[111] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[111]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[111]  <= \mchip.matrix_calculator.add_logic.shift1.Q [91];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [111] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[111] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[112] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[112]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[112]  <= \mchip.matrix_calculator.add_logic.shift1.Q [92];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [112] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[112] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[113] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[113]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[113]  <= \mchip.matrix_calculator.add_logic.shift1.Q [93];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [113] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[113] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[114] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[114]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[114]  <= \mchip.matrix_calculator.add_logic.shift1.Q [94];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [114] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[114] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[120] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[120]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[120]  <= \mchip.matrix_calculator.add_logic.shift1.Q [100];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [120] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[120] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[121] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[121]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[121]  <= \mchip.matrix_calculator.add_logic.shift1.Q [101];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [121] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[121] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[122] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[122]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[122]  <= \mchip.matrix_calculator.add_logic.shift1.Q [102];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [122] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[122] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[123] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[123]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[123]  <= \mchip.matrix_calculator.add_logic.shift1.Q [103];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [123] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[123] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[124] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[124]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[124]  <= \mchip.matrix_calculator.add_logic.shift1.Q [104];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [124] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[124] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[130] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[130]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[130]  <= \mchip.matrix_calculator.add_logic.shift1.Q [110];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [130] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[130] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[131] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[131]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[131]  <= \mchip.matrix_calculator.add_logic.shift1.Q [111];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [131] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[131] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[132] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[132]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[132]  <= \mchip.matrix_calculator.add_logic.shift1.Q [112];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [132] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[132] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[133] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[133]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[133]  <= \mchip.matrix_calculator.add_logic.shift1.Q [113];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [133] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[133] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[134] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[134]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[134]  <= \mchip.matrix_calculator.add_logic.shift1.Q [114];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [134] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[134] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[140] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[140]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[140]  <= \mchip.matrix_calculator.add_logic.shift1.Q [120];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [140] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[140] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[141] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[141]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[141]  <= \mchip.matrix_calculator.add_logic.shift1.Q [121];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [141] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[141] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[142] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[142]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[142]  <= \mchip.matrix_calculator.add_logic.shift1.Q [122];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [142] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[142] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[143] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[143]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[143]  <= \mchip.matrix_calculator.add_logic.shift1.Q [123];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [143] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[143] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[144] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[144]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[144]  <= \mchip.matrix_calculator.add_logic.shift1.Q [124];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [144] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[144] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[150] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[150]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[150]  <= \mchip.matrix_calculator.add_logic.shift1.Q [130];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [150] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[150] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[151] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[151]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[151]  <= \mchip.matrix_calculator.add_logic.shift1.Q [131];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [151] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[151] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[152] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[152]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[152]  <= \mchip.matrix_calculator.add_logic.shift1.Q [132];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [152] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[152] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[153] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[153]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[153]  <= \mchip.matrix_calculator.add_logic.shift1.Q [133];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [153] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[153] ;
	reg \mchip.matrix_calculator.add_logic.shift1.Q_reg[154] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[154]  <= 1'h0;
		else if (\mchip.matrix_calculator.add_logic.fsm.shift_en )
			\mchip.matrix_calculator.add_logic.shift1.Q_reg[154]  <= \mchip.matrix_calculator.add_logic.shift1.Q [134];
	assign \mchip.matrix_calculator.add_logic.shift1.Q [154] = \mchip.matrix_calculator.add_logic.shift1.Q_reg[154] ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [0] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [0] <= \mchip.sync1.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [1] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [1] <= \mchip.sync2.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [2] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [2] <= \mchip.sync3.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [3] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [3] <= \mchip.sync4.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [4] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [4] <= \mchip.sync5.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [5] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [5] <= \mchip.sync6.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [6] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [6] <= \mchip.sync7.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [7] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [7] <= \mchip.sync8.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [8] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [8] <= \mchip.matrix_calculator.shift_register.Q [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [9] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [9] <= \mchip.matrix_calculator.shift_register.Q [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [10] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [10] <= \mchip.matrix_calculator.shift_register.Q [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [11] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [11] <= \mchip.matrix_calculator.shift_register.Q [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [12] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [12] <= \mchip.matrix_calculator.shift_register.Q [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [13] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [13] <= \mchip.matrix_calculator.shift_register.Q [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [14] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [14] <= \mchip.matrix_calculator.shift_register.Q [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [15] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [15] <= \mchip.matrix_calculator.shift_register.Q [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [16] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [16] <= \mchip.matrix_calculator.shift_register.Q [8];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [17] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [17] <= \mchip.matrix_calculator.shift_register.Q [9];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [18] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [18] <= \mchip.matrix_calculator.shift_register.Q [10];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [19] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [19] <= \mchip.matrix_calculator.shift_register.Q [11];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [20] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [20] <= \mchip.matrix_calculator.shift_register.Q [12];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [21] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [21] <= \mchip.matrix_calculator.shift_register.Q [13];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [22] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [22] <= \mchip.matrix_calculator.shift_register.Q [14];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [23] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [23] <= \mchip.matrix_calculator.shift_register.Q [15];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [24] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [24] <= \mchip.matrix_calculator.shift_register.Q [16];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [25] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [25] <= \mchip.matrix_calculator.shift_register.Q [17];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [26] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [26] <= \mchip.matrix_calculator.shift_register.Q [18];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [27] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [27] <= \mchip.matrix_calculator.shift_register.Q [19];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [28] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [28] <= \mchip.matrix_calculator.shift_register.Q [20];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [29] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [29] <= \mchip.matrix_calculator.shift_register.Q [21];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [30] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [30] <= \mchip.matrix_calculator.shift_register.Q [22];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [31] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [31] <= \mchip.matrix_calculator.shift_register.Q [23];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [32] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [32] <= \mchip.matrix_calculator.shift_register.Q [24];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [33] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [33] <= \mchip.matrix_calculator.shift_register.Q [25];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [34] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [34] <= \mchip.matrix_calculator.shift_register.Q [26];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [35] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [35] <= \mchip.matrix_calculator.shift_register.Q [27];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [36] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [36] <= \mchip.matrix_calculator.shift_register.Q [28];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [37] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [37] <= \mchip.matrix_calculator.shift_register.Q [29];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [38] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [38] <= \mchip.matrix_calculator.shift_register.Q [30];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [39] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [39] <= \mchip.matrix_calculator.shift_register.Q [31];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [40] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [40] <= \mchip.matrix_calculator.shift_register.Q [32];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [41] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [41] <= \mchip.matrix_calculator.shift_register.Q [33];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [42] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [42] <= \mchip.matrix_calculator.shift_register.Q [34];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [43] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [43] <= \mchip.matrix_calculator.shift_register.Q [35];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [44] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [44] <= \mchip.matrix_calculator.shift_register.Q [36];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [45] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [45] <= \mchip.matrix_calculator.shift_register.Q [37];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [46] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [46] <= \mchip.matrix_calculator.shift_register.Q [38];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [47] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [47] <= \mchip.matrix_calculator.shift_register.Q [39];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [48] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [48] <= \mchip.matrix_calculator.shift_register.Q [40];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [49] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [49] <= \mchip.matrix_calculator.shift_register.Q [41];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [50] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [50] <= \mchip.matrix_calculator.shift_register.Q [42];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [51] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [51] <= \mchip.matrix_calculator.shift_register.Q [43];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [52] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [52] <= \mchip.matrix_calculator.shift_register.Q [44];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [53] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [53] <= \mchip.matrix_calculator.shift_register.Q [45];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [54] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [54] <= \mchip.matrix_calculator.shift_register.Q [46];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [55] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [55] <= \mchip.matrix_calculator.shift_register.Q [47];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [56] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [56] <= \mchip.matrix_calculator.shift_register.Q [48];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [57] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [57] <= \mchip.matrix_calculator.shift_register.Q [49];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [58] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [58] <= \mchip.matrix_calculator.shift_register.Q [50];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [59] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [59] <= \mchip.matrix_calculator.shift_register.Q [51];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [60] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [60] <= \mchip.matrix_calculator.shift_register.Q [52];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [61] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [61] <= \mchip.matrix_calculator.shift_register.Q [53];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [62] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [62] <= \mchip.matrix_calculator.shift_register.Q [54];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [63] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [63] <= \mchip.matrix_calculator.shift_register.Q [55];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [64] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [64] <= \mchip.matrix_calculator.shift_register.Q [56];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [65] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [65] <= \mchip.matrix_calculator.shift_register.Q [57];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [66] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [66] <= \mchip.matrix_calculator.shift_register.Q [58];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [67] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [67] <= \mchip.matrix_calculator.shift_register.Q [59];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [68] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [68] <= \mchip.matrix_calculator.shift_register.Q [60];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [69] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [69] <= \mchip.matrix_calculator.shift_register.Q [61];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [70] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [70] <= \mchip.matrix_calculator.shift_register.Q [62];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [71] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [71] <= \mchip.matrix_calculator.shift_register.Q [63];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [72] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [72] <= \mchip.matrix_calculator.shift_register.Q [64];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [73] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [73] <= \mchip.matrix_calculator.shift_register.Q [65];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [74] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [74] <= \mchip.matrix_calculator.shift_register.Q [66];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [75] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [75] <= \mchip.matrix_calculator.shift_register.Q [67];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [76] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [76] <= \mchip.matrix_calculator.shift_register.Q [68];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [77] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [77] <= \mchip.matrix_calculator.shift_register.Q [69];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [78] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [78] <= \mchip.matrix_calculator.shift_register.Q [70];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [79] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [79] <= \mchip.matrix_calculator.shift_register.Q [71];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [80] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [80] <= \mchip.matrix_calculator.shift_register.Q [72];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [81] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [81] <= \mchip.matrix_calculator.shift_register.Q [73];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [82] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [82] <= \mchip.matrix_calculator.shift_register.Q [74];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [83] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [83] <= \mchip.matrix_calculator.shift_register.Q [75];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [84] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [84] <= \mchip.matrix_calculator.shift_register.Q [76];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [85] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [85] <= \mchip.matrix_calculator.shift_register.Q [77];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [86] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [86] <= \mchip.matrix_calculator.shift_register.Q [78];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [87] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [87] <= \mchip.matrix_calculator.shift_register.Q [79];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [88] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [88] <= \mchip.matrix_calculator.shift_register.Q [80];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [89] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [89] <= \mchip.matrix_calculator.shift_register.Q [81];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [90] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [90] <= \mchip.matrix_calculator.shift_register.Q [82];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [91] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [91] <= \mchip.matrix_calculator.shift_register.Q [83];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [92] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [92] <= \mchip.matrix_calculator.shift_register.Q [84];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [93] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [93] <= \mchip.matrix_calculator.shift_register.Q [85];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [94] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [94] <= \mchip.matrix_calculator.shift_register.Q [86];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [95] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [95] <= \mchip.matrix_calculator.shift_register.Q [87];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [96] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [96] <= \mchip.matrix_calculator.shift_register.Q [88];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [97] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [97] <= \mchip.matrix_calculator.shift_register.Q [89];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [98] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [98] <= \mchip.matrix_calculator.shift_register.Q [90];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [99] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [99] <= \mchip.matrix_calculator.shift_register.Q [91];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [100] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [100] <= \mchip.matrix_calculator.shift_register.Q [92];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [101] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [101] <= \mchip.matrix_calculator.shift_register.Q [93];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [102] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [102] <= \mchip.matrix_calculator.shift_register.Q [94];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [103] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [103] <= \mchip.matrix_calculator.shift_register.Q [95];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [104] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [104] <= \mchip.matrix_calculator.shift_register.Q [96];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [105] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [105] <= \mchip.matrix_calculator.shift_register.Q [97];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [106] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [106] <= \mchip.matrix_calculator.shift_register.Q [98];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [107] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [107] <= \mchip.matrix_calculator.shift_register.Q [99];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [108] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [108] <= \mchip.matrix_calculator.shift_register.Q [100];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [109] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [109] <= \mchip.matrix_calculator.shift_register.Q [101];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [110] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [110] <= \mchip.matrix_calculator.shift_register.Q [102];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [111] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [111] <= \mchip.matrix_calculator.shift_register.Q [103];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [112] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [112] <= \mchip.matrix_calculator.shift_register.Q [104];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [113] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [113] <= \mchip.matrix_calculator.shift_register.Q [105];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [114] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [114] <= \mchip.matrix_calculator.shift_register.Q [106];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [115] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [115] <= \mchip.matrix_calculator.shift_register.Q [107];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [116] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [116] <= \mchip.matrix_calculator.shift_register.Q [108];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [117] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [117] <= \mchip.matrix_calculator.shift_register.Q [109];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [118] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [118] <= \mchip.matrix_calculator.shift_register.Q [110];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [119] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [119] <= \mchip.matrix_calculator.shift_register.Q [111];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [120] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [120] <= \mchip.matrix_calculator.shift_register.Q [112];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [121] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [121] <= \mchip.matrix_calculator.shift_register.Q [113];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [122] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [122] <= \mchip.matrix_calculator.shift_register.Q [114];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [123] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [123] <= \mchip.matrix_calculator.shift_register.Q [115];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [124] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [124] <= \mchip.matrix_calculator.shift_register.Q [116];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [125] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [125] <= \mchip.matrix_calculator.shift_register.Q [117];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [126] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [126] <= \mchip.matrix_calculator.shift_register.Q [118];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.shift_register.Q [127] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.shift_register.Q [127] <= \mchip.matrix_calculator.shift_register.Q [119];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.op_reg.Q [0] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.op_reg.Q [0] <= \mchip.sync11.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.op_reg.Q [1] <= 1'h0;
		else if (\mchip.matrix_calculator.op_reg.en )
			\mchip.matrix_calculator.op_reg.Q [1] <= \mchip.sync12.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [0] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [0] <= \mchip.matrix_calculator.mul_logic.add_out2 [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [1] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [1] <= \mchip.matrix_calculator.mul_logic.add_out2 [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [2] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [2] <= \mchip.matrix_calculator.mul_logic.add_out2 [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [3] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [3] <= \mchip.matrix_calculator.mul_logic.add_out2 [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [4] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [4] <= \mchip.matrix_calculator.mul_logic.add_out2 [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [5] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [5] <= \mchip.matrix_calculator.mul_logic.add_out2 [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [6] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [6] <= \mchip.matrix_calculator.mul_logic.add_out2 [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [7] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [7] <= \mchip.matrix_calculator.mul_logic.add_out2 [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [8] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [8] <= \mchip.matrix_calculator.mul_logic.add_out2 [8];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [9] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [9] <= \mchip.matrix_calculator.mul_logic.add_out2 [9];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [10] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [10] <= \mchip.matrix_calculator.mul_logic.add_out [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [11] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [11] <= \mchip.matrix_calculator.mul_logic.add_out [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [12] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [12] <= \mchip.matrix_calculator.mul_logic.add_out [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [13] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [13] <= \mchip.matrix_calculator.mul_logic.add_out [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [14] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [14] <= \mchip.matrix_calculator.mul_logic.add_out [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [15] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [15] <= \mchip.matrix_calculator.mul_logic.add_out [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [16] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [16] <= \mchip.matrix_calculator.mul_logic.add_out [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [17] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [17] <= \mchip.matrix_calculator.mul_logic.add_out [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [18] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [18] <= \mchip.matrix_calculator.mul_logic.add_out [8];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [19] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [19] <= \mchip.matrix_calculator.mul_logic.add_out [9];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [20] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [20] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [21] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [21] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [22] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [22] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [23] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [23] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [24] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [24] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [25] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [25] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [26] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [26] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [27] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [27] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [28] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [28] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [8];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [29] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [29] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [9];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [30] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [30] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [10];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [31] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [31] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [11];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [32] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [32] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [12];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [33] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [33] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [13];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [34] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [34] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [14];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [35] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [35] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [15];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [36] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [36] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [16];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [37] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [37] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [17];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [38] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [38] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [18];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [39] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [39] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [19];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [40] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [40] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [20];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [41] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [41] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [21];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [42] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [42] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [22];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [43] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [43] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [23];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [44] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [44] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [24];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [45] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [45] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [25];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [46] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [46] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [26];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [47] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [47] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [27];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [48] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [48] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [28];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [49] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [49] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [29];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [50] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [50] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [30];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [51] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [51] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [31];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [52] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [52] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [32];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [53] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [53] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [33];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [54] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [54] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [34];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [55] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [55] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [35];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [56] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [56] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [36];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [57] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [57] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [37];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [58] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [58] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [38];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [59] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [59] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [39];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [60] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [60] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [40];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [61] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [61] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [41];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [62] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [62] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [42];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [63] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [63] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [43];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [64] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [64] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [44];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [65] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [65] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [45];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [66] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [66] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [46];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [67] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [67] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [47];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [68] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [68] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [48];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [69] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [69] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [49];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [70] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [70] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [50];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [71] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [71] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [51];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [72] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [72] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [52];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [73] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [73] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [53];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [74] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [74] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [54];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [75] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [75] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [55];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [76] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [76] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [56];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [77] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [77] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [57];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [78] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [78] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [58];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [79] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [79] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [59];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [80] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [80] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [60];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [81] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [81] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [61];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [82] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [82] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [62];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [83] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [83] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [63];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [84] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [84] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [64];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [85] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [85] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [65];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [86] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [86] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [66];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [87] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [87] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [67];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [88] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [88] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [68];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [89] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [89] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [69];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [90] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [90] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [70];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [91] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [91] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [71];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [92] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [92] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [72];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [93] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [93] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [73];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [94] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [94] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [74];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [95] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [95] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [75];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [96] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [96] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [76];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [97] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [97] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [77];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [98] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [98] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [78];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [99] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [99] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [79];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [100] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [100] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [80];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [101] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [101] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [81];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [102] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [102] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [82];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [103] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [103] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [83];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [104] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [104] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [84];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [105] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [105] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [85];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [106] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [106] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [86];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [107] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [107] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [87];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [108] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [108] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [88];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [109] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [109] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [89];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [110] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [110] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [90];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [111] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [111] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [91];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [112] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [112] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [92];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [113] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [113] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [93];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [114] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [114] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [94];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [115] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [115] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [95];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [116] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [116] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [96];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [117] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [117] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [97];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [118] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [118] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [98];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [119] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [119] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [99];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [120] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [120] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [100];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [121] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [121] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [101];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [122] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [122] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [102];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [123] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [123] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [103];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [124] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [124] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [104];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [125] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [125] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [105];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [126] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [126] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [106];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [127] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [127] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [107];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [128] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [128] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [108];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [129] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [129] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [109];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [130] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [130] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [110];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [131] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [131] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [111];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [132] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [132] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [112];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [133] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [133] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [113];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [134] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [134] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [114];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [135] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [135] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [115];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [136] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [136] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [116];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [137] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [137] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [117];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [138] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [138] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [118];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [139] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [139] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [119];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [140] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [140] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [120];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [141] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [141] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [121];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [142] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [142] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [122];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [143] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [143] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [123];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [144] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [144] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [124];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [145] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [145] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [125];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [146] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [146] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [126];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [147] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [147] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [127];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [148] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [148] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [128];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [149] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [149] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [129];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [150] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [150] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [130];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [151] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [151] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [131];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [152] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [152] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [132];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [153] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [153] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [133];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [154] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [154] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [134];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [155] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [155] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [135];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [156] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [156] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [136];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [157] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [157] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [137];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [158] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [158] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [138];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [159] <= 1'h0;
		else if (\mchip.matrix_calculator.mul_logic.fsm.layer_2_en )
			\mchip.matrix_calculator.mul_logic.shift_register.Q [159] <= \mchip.matrix_calculator.mul_logic.shift_register.Q [139];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [0] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [0] <= \mchip.matrix_calculator.mul_logic.mult8.S [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [1] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [1] <= \mchip.matrix_calculator.mul_logic.mult8.S [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [2] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [2] <= \mchip.matrix_calculator.mul_logic.mult8.S [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [3] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [3] <= \mchip.matrix_calculator.mul_logic.mult8.S [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [4] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [4] <= \mchip.matrix_calculator.mul_logic.mult8.S [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [5] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [5] <= \mchip.matrix_calculator.mul_logic.mult8.S [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [6] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [6] <= \mchip.matrix_calculator.mul_logic.mult8.S [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [7] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [7] <= \mchip.matrix_calculator.mul_logic.mult8.S [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [8] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [8] <= \mchip.matrix_calculator.mul_logic.mult7.S [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [9] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [9] <= \mchip.matrix_calculator.mul_logic.mult7.S [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [10] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [10] <= \mchip.matrix_calculator.mul_logic.mult7.S [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [11] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [11] <= \mchip.matrix_calculator.mul_logic.mult7.S [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [12] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [12] <= \mchip.matrix_calculator.mul_logic.mult7.S [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [13] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [13] <= \mchip.matrix_calculator.mul_logic.mult7.S [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [14] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [14] <= \mchip.matrix_calculator.mul_logic.mult7.S [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [15] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [15] <= \mchip.matrix_calculator.mul_logic.mult7.S [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [16] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [16] <= \mchip.matrix_calculator.mul_logic.mult6.S [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [17] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [17] <= \mchip.matrix_calculator.mul_logic.mult6.S [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [18] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [18] <= \mchip.matrix_calculator.mul_logic.mult6.S [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [19] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [19] <= \mchip.matrix_calculator.mul_logic.mult6.S [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [20] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [20] <= \mchip.matrix_calculator.mul_logic.mult6.S [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [21] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [21] <= \mchip.matrix_calculator.mul_logic.mult6.S [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [22] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [22] <= \mchip.matrix_calculator.mul_logic.mult6.S [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [23] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [23] <= \mchip.matrix_calculator.mul_logic.mult6.S [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [24] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [24] <= \mchip.matrix_calculator.mul_logic.mult5.S [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [25] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [25] <= \mchip.matrix_calculator.mul_logic.mult5.S [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [26] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [26] <= \mchip.matrix_calculator.mul_logic.mult5.S [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [27] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [27] <= \mchip.matrix_calculator.mul_logic.mult5.S [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [28] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [28] <= \mchip.matrix_calculator.mul_logic.mult5.S [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [29] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [29] <= \mchip.matrix_calculator.mul_logic.mult5.S [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [30] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [30] <= \mchip.matrix_calculator.mul_logic.mult5.S [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [31] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [31] <= \mchip.matrix_calculator.mul_logic.mult5.S [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [0] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [0] <= \mchip.matrix_calculator.mul_logic.mult4.S [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [1] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [1] <= \mchip.matrix_calculator.mul_logic.mult4.S [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [2] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [2] <= \mchip.matrix_calculator.mul_logic.mult4.S [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [3] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [3] <= \mchip.matrix_calculator.mul_logic.mult4.S [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [4] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [4] <= \mchip.matrix_calculator.mul_logic.mult4.S [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [5] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [5] <= \mchip.matrix_calculator.mul_logic.mult4.S [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [6] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [6] <= \mchip.matrix_calculator.mul_logic.mult4.S [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [7] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [7] <= \mchip.matrix_calculator.mul_logic.mult4.S [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [8] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [8] <= \mchip.matrix_calculator.mul_logic.mult3.S [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [9] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [9] <= \mchip.matrix_calculator.mul_logic.mult3.S [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [10] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [10] <= \mchip.matrix_calculator.mul_logic.mult3.S [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [11] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [11] <= \mchip.matrix_calculator.mul_logic.mult3.S [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [12] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [12] <= \mchip.matrix_calculator.mul_logic.mult3.S [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [13] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [13] <= \mchip.matrix_calculator.mul_logic.mult3.S [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [14] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [14] <= \mchip.matrix_calculator.mul_logic.mult3.S [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [15] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [15] <= \mchip.matrix_calculator.mul_logic.mult3.S [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [16] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [16] <= \mchip.matrix_calculator.mul_logic.mult2.S [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [17] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [17] <= \mchip.matrix_calculator.mul_logic.mult2.S [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [18] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [18] <= \mchip.matrix_calculator.mul_logic.mult2.S [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [19] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [19] <= \mchip.matrix_calculator.mul_logic.mult2.S [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [20] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [20] <= \mchip.matrix_calculator.mul_logic.mult2.S [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [21] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [21] <= \mchip.matrix_calculator.mul_logic.mult2.S [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [22] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [22] <= \mchip.matrix_calculator.mul_logic.mult2.S [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [23] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [23] <= \mchip.matrix_calculator.mul_logic.mult2.S [7];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [24] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [24] <= \mchip.matrix_calculator.mul_logic.mult1.S [0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [25] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [25] <= \mchip.matrix_calculator.mul_logic.mult1.S [1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [26] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [26] <= \mchip.matrix_calculator.mul_logic.mult1.S [2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [27] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [27] <= \mchip.matrix_calculator.mul_logic.mult1.S [3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [28] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [28] <= \mchip.matrix_calculator.mul_logic.mult1.S [4];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [29] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [29] <= \mchip.matrix_calculator.mul_logic.mult1.S [5];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [30] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [30] <= \mchip.matrix_calculator.mul_logic.mult1.S [6];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [31] <= 1'h0;
		else if (!_0042_)
			\mchip.matrix_calculator.mul_logic.layer_1_reg.Q [31] <= \mchip.matrix_calculator.mul_logic.mult1.S [7];
	always @(posedge io_in[12]) \mchip.matrix_calculator.sw_de.tmp1  <= \mchip.sync10.sync ;
	always @(posedge io_in[12]) \mchip.matrix_calculator.ed_de.tmp1  <= \mchip.sync9.sync ;
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.index_counter.Q [0] <= 1'h0;
		else if (\mchip.matrix_calculator.index_counter.en )
			\mchip.matrix_calculator.index_counter.Q [0] <= _2025_[0];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.index_counter.Q [1] <= 1'h0;
		else if (\mchip.matrix_calculator.index_counter.en )
			\mchip.matrix_calculator.index_counter.Q [1] <= _2026_[1];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.index_counter.Q [2] <= 1'h0;
		else if (\mchip.matrix_calculator.index_counter.en )
			\mchip.matrix_calculator.index_counter.Q [2] <= _2026_[2];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.index_counter.Q [3] <= 1'h0;
		else if (\mchip.matrix_calculator.index_counter.en )
			\mchip.matrix_calculator.index_counter.Q [3] <= _2026_[3];
	always @(posedge io_in[12])
		if (\mchip.sync13.sync )
			\mchip.matrix_calculator.index_counter.Q [4] <= 1'h0;
		else if (\mchip.matrix_calculator.index_counter.en )
			\mchip.matrix_calculator.index_counter.Q [4] <= _2026_[4];
	always @(posedge io_in[12]) \mchip.sync13.tmp1  <= io_in[13];
	always @(posedge io_in[12]) \mchip.sync12.tmp1  <= io_in[11];
	always @(posedge io_in[12]) \mchip.sync11.tmp1  <= io_in[10];
	always @(posedge io_in[12]) \mchip.sync10.tmp1  <= io_in[9];
	always @(posedge io_in[12]) \mchip.sync9.tmp1  <= io_in[8];
	always @(posedge io_in[12]) \mchip.sync8.tmp1  <= io_in[7];
	always @(posedge io_in[12]) \mchip.sync7.tmp1  <= io_in[6];
	always @(posedge io_in[12]) \mchip.sync6.tmp1  <= io_in[5];
	always @(posedge io_in[12]) \mchip.sync5.tmp1  <= io_in[4];
	always @(posedge io_in[12]) \mchip.sync4.tmp1  <= io_in[3];
	always @(posedge io_in[12]) \mchip.sync3.tmp1  <= io_in[2];
	always @(posedge io_in[12]) \mchip.sync2.tmp1  <= io_in[1];
	always @(posedge io_in[12]) \mchip.sync1.tmp1  <= io_in[0];
	always @(posedge io_in[12]) \mchip.sync13.sync  <= \mchip.sync13.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync12.sync  <= \mchip.sync12.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync11.sync  <= \mchip.sync11.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync10.sync  <= \mchip.sync10.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync9.sync  <= \mchip.sync9.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync8.sync  <= \mchip.sync8.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync7.sync  <= \mchip.sync7.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync6.sync  <= \mchip.sync6.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync5.sync  <= \mchip.sync5.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync4.sync  <= \mchip.sync4.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync3.sync  <= \mchip.sync3.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync2.sync  <= \mchip.sync2.tmp1 ;
	always @(posedge io_in[12]) \mchip.sync1.sync  <= \mchip.sync1.tmp1 ;
	assign _2025_[4:1] = \mchip.matrix_calculator.index_counter.Q [4:1];
	assign _2026_[0] = _2025_[0];
	assign io_out[13:5] = {3'h0, \mchip.matrix_calculator.index_counter.Q [4:1], \mchip.error , \mchip.finish };
	assign \mchip.clock  = io_in[12];
	assign \mchip.data_in  = {\mchip.sync8.sync , \mchip.sync7.sync , \mchip.sync6.sync , \mchip.sync5.sync , \mchip.sync4.sync , \mchip.sync3.sync , \mchip.sync2.sync , \mchip.sync1.sync };
	assign \mchip.data_out  = io_out[4:0];
	assign \mchip.enter  = \mchip.sync9.sync ;
	assign \mchip.index  = \mchip.matrix_calculator.index_counter.Q [4:1];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {1'h0, \mchip.matrix_calculator.index_counter.Q [4:1], \mchip.error , \mchip.finish , io_out[4:0]};
	assign \mchip.matrix_calculator.add_finish  = \mchip.matrix_calculator.add_logic.fsm.cur_state [6];
	assign \mchip.matrix_calculator.add_logic.add1_out  = \mchip.matrix_calculator.add_logic.add1.S ;
	assign \mchip.matrix_calculator.add_logic.add2_out  = \mchip.matrix_calculator.add_logic.add2.S ;
	assign \mchip.matrix_calculator.add_logic.clk  = io_in[12];
	assign \mchip.matrix_calculator.add_logic.finish  = \mchip.matrix_calculator.add_logic.fsm.cur_state [6];
	assign \mchip.matrix_calculator.add_logic.fsm.clk  = io_in[12];
	assign \mchip.matrix_calculator.add_logic.fsm.finish  = \mchip.matrix_calculator.add_logic.fsm.cur_state [6];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A  = \mchip.matrix_calculator.shift_register.Q [127:64];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_1  = \mchip.matrix_calculator.shift_register.Q [127:124];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_10  = \mchip.matrix_calculator.shift_register.Q [91:88];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_11  = \mchip.matrix_calculator.shift_register.Q [87:84];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_12  = \mchip.matrix_calculator.shift_register.Q [83:80];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_13  = \mchip.matrix_calculator.shift_register.Q [79:76];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_14  = \mchip.matrix_calculator.shift_register.Q [75:72];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_15  = \mchip.matrix_calculator.shift_register.Q [71:68];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_16  = \mchip.matrix_calculator.shift_register.Q [67:64];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_2  = \mchip.matrix_calculator.shift_register.Q [123:120];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_3  = \mchip.matrix_calculator.shift_register.Q [119:116];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_4  = \mchip.matrix_calculator.shift_register.Q [115:112];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_5  = \mchip.matrix_calculator.shift_register.Q [111:108];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_6  = \mchip.matrix_calculator.shift_register.Q [107:104];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_7  = \mchip.matrix_calculator.shift_register.Q [103:100];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_8  = \mchip.matrix_calculator.shift_register.Q [99:96];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_A_9  = \mchip.matrix_calculator.shift_register.Q [95:92];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B  = \mchip.matrix_calculator.shift_register.Q [63:0];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_1  = \mchip.matrix_calculator.shift_register.Q [63:60];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_10  = \mchip.matrix_calculator.shift_register.Q [27:24];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_11  = \mchip.matrix_calculator.shift_register.Q [23:20];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_12  = \mchip.matrix_calculator.shift_register.Q [19:16];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_13  = \mchip.matrix_calculator.shift_register.Q [15:12];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_14  = \mchip.matrix_calculator.shift_register.Q [11:8];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_15  = \mchip.matrix_calculator.shift_register.Q [7:4];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_16  = \mchip.matrix_calculator.shift_register.Q [3:0];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_2  = \mchip.matrix_calculator.shift_register.Q [59:56];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_3  = \mchip.matrix_calculator.shift_register.Q [55:52];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_4  = \mchip.matrix_calculator.shift_register.Q [51:48];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_5  = \mchip.matrix_calculator.shift_register.Q [47:44];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_6  = \mchip.matrix_calculator.shift_register.Q [43:40];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_7  = \mchip.matrix_calculator.shift_register.Q [39:36];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_8  = \mchip.matrix_calculator.shift_register.Q [35:32];
	assign \mchip.matrix_calculator.add_logic.fsm.mat_B_9  = \mchip.matrix_calculator.shift_register.Q [31:28];
	assign \mchip.matrix_calculator.add_logic.fsm.rst  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.add_logic.mat_A  = \mchip.matrix_calculator.shift_register.Q [127:64];
	assign \mchip.matrix_calculator.add_logic.mat_B  = \mchip.matrix_calculator.shift_register.Q [63:0];
	assign \mchip.matrix_calculator.add_logic.mat_out  = {5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [154:150], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [144:140], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [134:130], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [124:120], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [114:110], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [104:100], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [94:90], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [84:80], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [74:70], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [64:60], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [54:50], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [44:40], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [34:30], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [24:20], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [14:10], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [4:0]};
	assign \mchip.matrix_calculator.add_logic.rst  = \mchip.sync13.sync ;
	assign {\mchip.matrix_calculator.add_logic.shift1.Q [159:155], \mchip.matrix_calculator.add_logic.shift1.Q [149:145], \mchip.matrix_calculator.add_logic.shift1.Q [139:135], \mchip.matrix_calculator.add_logic.shift1.Q [129:125], \mchip.matrix_calculator.add_logic.shift1.Q [119:115], \mchip.matrix_calculator.add_logic.shift1.Q [109:105], \mchip.matrix_calculator.add_logic.shift1.Q [99:95], \mchip.matrix_calculator.add_logic.shift1.Q [89:85], \mchip.matrix_calculator.add_logic.shift1.Q [79:75], \mchip.matrix_calculator.add_logic.shift1.Q [69:65], \mchip.matrix_calculator.add_logic.shift1.Q [59:55], \mchip.matrix_calculator.add_logic.shift1.Q [49:45], \mchip.matrix_calculator.add_logic.shift1.Q [39:35], \mchip.matrix_calculator.add_logic.shift1.Q [29:25], \mchip.matrix_calculator.add_logic.shift1.Q [19:15], \mchip.matrix_calculator.add_logic.shift1.Q [9:5]} = 80'h00000000000000000000;
	assign \mchip.matrix_calculator.add_logic.shift1.clock  = io_in[12];
	assign \mchip.matrix_calculator.add_logic.shift1.data_in  = {5'h00, \mchip.matrix_calculator.add_logic.add1.S , 5'h00, \mchip.matrix_calculator.add_logic.add2.S };
	assign \mchip.matrix_calculator.add_logic.shift1.en  = \mchip.matrix_calculator.add_logic.fsm.shift_en ;
	assign \mchip.matrix_calculator.add_logic.shift1.rst  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.add_logic.shift_en  = \mchip.matrix_calculator.add_logic.fsm.shift_en ;
	assign \mchip.matrix_calculator.add_logic.shift_in  = {5'h00, \mchip.matrix_calculator.add_logic.add1.S , 5'h00, \mchip.matrix_calculator.add_logic.add2.S };
	assign \mchip.matrix_calculator.add_logic.sign  = \mchip.matrix_calculator.op_reg.Q [0];
	assign \mchip.matrix_calculator.add_output  = {5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [154:150], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [144:140], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [134:130], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [124:120], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [114:110], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [104:100], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [94:90], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [84:80], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [74:70], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [64:60], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [54:50], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [44:40], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [34:30], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [24:20], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [14:10], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [4:0]};
	assign \mchip.matrix_calculator.clk  = io_in[12];
	assign \mchip.matrix_calculator.data_in  = {\mchip.sync8.sync , \mchip.sync7.sync , \mchip.sync6.sync , \mchip.sync5.sync , \mchip.sync4.sync , \mchip.sync3.sync , \mchip.sync2.sync , \mchip.sync1.sync };
	assign \mchip.matrix_calculator.data_out  = io_out[4:0];
	assign \mchip.matrix_calculator.ed_de.clk  = io_in[12];
	assign \mchip.matrix_calculator.ed_de.signal  = \mchip.sync9.sync ;
	assign \mchip.matrix_calculator.enter  = \mchip.sync9.sync ;
	assign \mchip.matrix_calculator.error  = \mchip.error ;
	assign \mchip.matrix_calculator.finish  = \mchip.finish ;
	assign \mchip.matrix_calculator.fsm.add_finish  = \mchip.matrix_calculator.add_logic.fsm.cur_state [6];
	assign \mchip.matrix_calculator.fsm.clk  = io_in[12];
	assign \mchip.matrix_calculator.fsm.error  = \mchip.error ;
	assign \mchip.matrix_calculator.fsm.finish  = \mchip.finish ;
	assign \mchip.matrix_calculator.fsm.input_op  = \mchip.matrix_calculator.op_reg.Q ;
	assign \mchip.matrix_calculator.fsm.mul_finish  = \mchip.matrix_calculator.mul_logic.fsm.cur_state [4];
	assign \mchip.matrix_calculator.fsm.rst  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.index  = \mchip.matrix_calculator.index_counter.Q [4:1];
	assign \mchip.matrix_calculator.index_count  = \mchip.matrix_calculator.index_counter.Q ;
	assign \mchip.matrix_calculator.index_counter.clear  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.index_counter.clock  = io_in[12];
	assign \mchip.matrix_calculator.input_matrix  = \mchip.matrix_calculator.shift_register.Q ;
	assign \mchip.matrix_calculator.input_matrix_A  = \mchip.matrix_calculator.shift_register.Q [127:64];
	assign \mchip.matrix_calculator.input_matrix_B  = \mchip.matrix_calculator.shift_register.Q [63:0];
	assign \mchip.matrix_calculator.input_op  = \mchip.matrix_calculator.op_reg.Q ;
	assign \mchip.matrix_calculator.mul_finish  = \mchip.matrix_calculator.mul_logic.fsm.cur_state [4];
	assign \mchip.matrix_calculator.mul_logic.add_in1  = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [31:24];
	assign \mchip.matrix_calculator.mul_logic.add_in2  = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [23:16];
	assign \mchip.matrix_calculator.mul_logic.add_in3  = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [15:8];
	assign \mchip.matrix_calculator.mul_logic.add_in4  = \mchip.matrix_calculator.mul_logic.layer_1_reg.Q [7:0];
	assign \mchip.matrix_calculator.mul_logic.add_in5  = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [31:24];
	assign \mchip.matrix_calculator.mul_logic.add_in6  = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [23:16];
	assign \mchip.matrix_calculator.mul_logic.add_in7  = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [15:8];
	assign \mchip.matrix_calculator.mul_logic.add_in8  = \mchip.matrix_calculator.mul_logic.layer_1_2_reg.Q [7:0];
	assign \mchip.matrix_calculator.mul_logic.clk  = io_in[12];
	assign \mchip.matrix_calculator.mul_logic.finish  = \mchip.matrix_calculator.mul_logic.fsm.cur_state [4];
	assign \mchip.matrix_calculator.mul_logic.fsm.clk  = io_in[12];
	assign \mchip.matrix_calculator.mul_logic.fsm.finish  = \mchip.matrix_calculator.mul_logic.fsm.cur_state [4];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A  = \mchip.matrix_calculator.shift_register.Q [127:64];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_1  = \mchip.matrix_calculator.shift_register.Q [127:124];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_10  = \mchip.matrix_calculator.shift_register.Q [91:88];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_11  = \mchip.matrix_calculator.shift_register.Q [87:84];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_12  = \mchip.matrix_calculator.shift_register.Q [83:80];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_13  = \mchip.matrix_calculator.shift_register.Q [79:76];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_14  = \mchip.matrix_calculator.shift_register.Q [75:72];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_15  = \mchip.matrix_calculator.shift_register.Q [71:68];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_16  = \mchip.matrix_calculator.shift_register.Q [67:64];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_2  = \mchip.matrix_calculator.shift_register.Q [123:120];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_3  = \mchip.matrix_calculator.shift_register.Q [119:116];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_4  = \mchip.matrix_calculator.shift_register.Q [115:112];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_5  = \mchip.matrix_calculator.shift_register.Q [111:108];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_6  = \mchip.matrix_calculator.shift_register.Q [107:104];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_7  = \mchip.matrix_calculator.shift_register.Q [103:100];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_8  = \mchip.matrix_calculator.shift_register.Q [99:96];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_A_9  = \mchip.matrix_calculator.shift_register.Q [95:92];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B  = \mchip.matrix_calculator.shift_register.Q [63:0];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_1  = \mchip.matrix_calculator.shift_register.Q [63:60];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_10  = \mchip.matrix_calculator.shift_register.Q [27:24];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_11  = \mchip.matrix_calculator.shift_register.Q [23:20];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_12  = \mchip.matrix_calculator.shift_register.Q [19:16];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_13  = \mchip.matrix_calculator.shift_register.Q [15:12];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_14  = \mchip.matrix_calculator.shift_register.Q [11:8];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_15  = \mchip.matrix_calculator.shift_register.Q [7:4];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_16  = \mchip.matrix_calculator.shift_register.Q [3:0];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_2  = \mchip.matrix_calculator.shift_register.Q [59:56];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_3  = \mchip.matrix_calculator.shift_register.Q [55:52];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_4  = \mchip.matrix_calculator.shift_register.Q [51:48];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_5  = \mchip.matrix_calculator.shift_register.Q [47:44];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_6  = \mchip.matrix_calculator.shift_register.Q [43:40];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_7  = \mchip.matrix_calculator.shift_register.Q [39:36];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_8  = \mchip.matrix_calculator.shift_register.Q [35:32];
	assign \mchip.matrix_calculator.mul_logic.fsm.mat_B_9  = \mchip.matrix_calculator.shift_register.Q [31:28];
	assign \mchip.matrix_calculator.mul_logic.fsm.rst  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.mul_logic.layer_1_2_reg.D  = {\mchip.matrix_calculator.mul_logic.mult5.S , \mchip.matrix_calculator.mul_logic.mult6.S , \mchip.matrix_calculator.mul_logic.mult7.S , \mchip.matrix_calculator.mul_logic.mult8.S };
	assign \mchip.matrix_calculator.mul_logic.layer_1_2_reg.clear  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.mul_logic.layer_1_2_reg.clock  = io_in[12];
	assign \mchip.matrix_calculator.mul_logic.layer_1_reg.D  = {\mchip.matrix_calculator.mul_logic.mult1.S , \mchip.matrix_calculator.mul_logic.mult2.S , \mchip.matrix_calculator.mul_logic.mult3.S , \mchip.matrix_calculator.mul_logic.mult4.S };
	assign \mchip.matrix_calculator.mul_logic.layer_1_reg.clear  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.mul_logic.layer_1_reg.clock  = io_in[12];
	assign \mchip.matrix_calculator.mul_logic.layer_2_en  = \mchip.matrix_calculator.mul_logic.fsm.layer_2_en ;
	assign \mchip.matrix_calculator.mul_logic.mat_A  = \mchip.matrix_calculator.shift_register.Q [127:64];
	assign \mchip.matrix_calculator.mul_logic.mat_B  = \mchip.matrix_calculator.shift_register.Q [63:0];
	assign \mchip.matrix_calculator.mul_logic.mat_out  = \mchip.matrix_calculator.mul_logic.shift_register.Q ;
	assign \mchip.matrix_calculator.mul_logic.mult1_out  = \mchip.matrix_calculator.mul_logic.mult1.S ;
	assign \mchip.matrix_calculator.mul_logic.mult2_out  = \mchip.matrix_calculator.mul_logic.mult2.S ;
	assign \mchip.matrix_calculator.mul_logic.mult3_out  = \mchip.matrix_calculator.mul_logic.mult3.S ;
	assign \mchip.matrix_calculator.mul_logic.mult4_out  = \mchip.matrix_calculator.mul_logic.mult4.S ;
	assign \mchip.matrix_calculator.mul_logic.mult5_out  = \mchip.matrix_calculator.mul_logic.mult5.S ;
	assign \mchip.matrix_calculator.mul_logic.mult6_out  = \mchip.matrix_calculator.mul_logic.mult6.S ;
	assign \mchip.matrix_calculator.mul_logic.mult7_out  = \mchip.matrix_calculator.mul_logic.mult7.S ;
	assign \mchip.matrix_calculator.mul_logic.mult8_out  = \mchip.matrix_calculator.mul_logic.mult8.S ;
	assign \mchip.matrix_calculator.mul_logic.rst  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.mul_logic.shift_register.clock  = io_in[12];
	assign \mchip.matrix_calculator.mul_logic.shift_register.data_in  = {\mchip.matrix_calculator.mul_logic.add_out , \mchip.matrix_calculator.mul_logic.add_out2 };
	assign \mchip.matrix_calculator.mul_logic.shift_register.en  = \mchip.matrix_calculator.mul_logic.fsm.layer_2_en ;
	assign \mchip.matrix_calculator.mul_logic.shift_register.rst  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.mul_output  = \mchip.matrix_calculator.mul_logic.shift_register.Q ;
	assign \mchip.matrix_calculator.op_reg.D  = {\mchip.sync12.sync , \mchip.sync11.sync };
	assign \mchip.matrix_calculator.op_reg.clear  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.op_reg.clock  = io_in[12];
	assign \mchip.matrix_calculator.operation  = {\mchip.sync12.sync , \mchip.sync11.sync };
	assign \mchip.matrix_calculator.output_mux.I0  = \mchip.matrix_calculator.mul_logic.shift_register.Q ;
	assign \mchip.matrix_calculator.output_mux.I1  = {5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [154:150], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [144:140], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [134:130], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [124:120], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [114:110], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [104:100], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [94:90], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [84:80], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [74:70], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [64:60], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [54:50], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [44:40], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [34:30], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [24:20], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [14:10], 5'h00, \mchip.matrix_calculator.add_logic.shift1.Q [4:0]};
	assign \mchip.matrix_calculator.output_mux.S  = \mchip.matrix_calculator.op_reg.Q [1];
	assign \mchip.matrix_calculator.rst  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.shift_register.clock  = io_in[12];
	assign \mchip.matrix_calculator.shift_register.data_in  = {\mchip.sync8.sync , \mchip.sync7.sync , \mchip.sync6.sync , \mchip.sync5.sync , \mchip.sync4.sync , \mchip.sync3.sync , \mchip.sync2.sync , \mchip.sync1.sync };
	assign \mchip.matrix_calculator.shift_register.en  = \mchip.matrix_calculator.op_reg.en ;
	assign \mchip.matrix_calculator.shift_register.rst  = \mchip.sync13.sync ;
	assign \mchip.matrix_calculator.sw  = \mchip.sync10.sync ;
	assign \mchip.matrix_calculator.sw_de.clk  = io_in[12];
	assign \mchip.matrix_calculator.sw_de.signal  = \mchip.sync10.sync ;
	assign \mchip.operation  = {\mchip.sync12.sync , \mchip.sync11.sync };
	assign \mchip.reset  = io_in[13];
	assign \mchip.rst  = \mchip.sync13.sync ;
	assign \mchip.sw  = \mchip.sync10.sync ;
	assign \mchip.sync1.async  = io_in[0];
	assign \mchip.sync1.clock  = io_in[12];
	assign \mchip.sync1.tmp2  = \mchip.sync1.tmp1 ;
	assign \mchip.sync10.async  = io_in[9];
	assign \mchip.sync10.clock  = io_in[12];
	assign \mchip.sync10.tmp2  = \mchip.sync10.tmp1 ;
	assign \mchip.sync11.async  = io_in[10];
	assign \mchip.sync11.clock  = io_in[12];
	assign \mchip.sync11.tmp2  = \mchip.sync11.tmp1 ;
	assign \mchip.sync12.async  = io_in[11];
	assign \mchip.sync12.clock  = io_in[12];
	assign \mchip.sync12.tmp2  = \mchip.sync12.tmp1 ;
	assign \mchip.sync13.async  = io_in[13];
	assign \mchip.sync13.clock  = io_in[12];
	assign \mchip.sync13.tmp2  = \mchip.sync13.tmp1 ;
	assign \mchip.sync2.async  = io_in[1];
	assign \mchip.sync2.clock  = io_in[12];
	assign \mchip.sync2.tmp2  = \mchip.sync2.tmp1 ;
	assign \mchip.sync3.async  = io_in[2];
	assign \mchip.sync3.clock  = io_in[12];
	assign \mchip.sync3.tmp2  = \mchip.sync3.tmp1 ;
	assign \mchip.sync4.async  = io_in[3];
	assign \mchip.sync4.clock  = io_in[12];
	assign \mchip.sync4.tmp2  = \mchip.sync4.tmp1 ;
	assign \mchip.sync5.async  = io_in[4];
	assign \mchip.sync5.clock  = io_in[12];
	assign \mchip.sync5.tmp2  = \mchip.sync5.tmp1 ;
	assign \mchip.sync6.async  = io_in[5];
	assign \mchip.sync6.clock  = io_in[12];
	assign \mchip.sync6.tmp2  = \mchip.sync6.tmp1 ;
	assign \mchip.sync7.async  = io_in[6];
	assign \mchip.sync7.clock  = io_in[12];
	assign \mchip.sync7.tmp2  = \mchip.sync7.tmp1 ;
	assign \mchip.sync8.async  = io_in[7];
	assign \mchip.sync8.clock  = io_in[12];
	assign \mchip.sync8.tmp2  = \mchip.sync8.tmp1 ;
	assign \mchip.sync9.async  = io_in[8];
	assign \mchip.sync9.clock  = io_in[12];
	assign \mchip.sync9.tmp2  = \mchip.sync9.tmp1 ;
endmodule
module d15_spencer2_pianotiles (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	reg _0044_;
	reg _0045_;
	reg _0046_;
	reg _0047_;
	reg _0048_;
	reg _0049_;
	reg _0050_;
	reg _0051_;
	reg _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire [11:0] _0509_;
	wire [11:0] _0510_;
	wire [4:0] _0511_;
	wire [4:0] _0512_;
	wire [2:0] _0513_;
	wire [6:0] _0514_;
	wire [6:0] _0515_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.my_chip.async2sync0.async ;
	wire \mchip.my_chip.async2sync0.clk ;
	reg \mchip.my_chip.async2sync0.metastable ;
	reg \mchip.my_chip.async2sync0.sync ;
	wire \mchip.my_chip.async2sync1.async ;
	wire \mchip.my_chip.async2sync1.clk ;
	reg \mchip.my_chip.async2sync1.metastable ;
	reg \mchip.my_chip.async2sync1.sync ;
	wire \mchip.my_chip.async2sync2.async ;
	wire \mchip.my_chip.async2sync2.clk ;
	reg \mchip.my_chip.async2sync2.metastable ;
	reg \mchip.my_chip.async2sync2.sync ;
	wire \mchip.my_chip.async2sync3.async ;
	wire \mchip.my_chip.async2sync3.clk ;
	reg \mchip.my_chip.async2sync3.metastable ;
	reg \mchip.my_chip.async2sync3.sync ;
	wire \mchip.my_chip.async2sync4.async ;
	wire \mchip.my_chip.async2sync4.clk ;
	reg \mchip.my_chip.async2sync4.metastable ;
	reg \mchip.my_chip.async2sync4.sync ;
	wire \mchip.my_chip.async2sync5.async ;
	wire \mchip.my_chip.async2sync5.clk ;
	reg \mchip.my_chip.async2sync5.metastable ;
	reg \mchip.my_chip.async2sync5.sync ;
	wire \mchip.my_chip.async2sync6.async ;
	wire \mchip.my_chip.async2sync6.clk ;
	reg \mchip.my_chip.async2sync6.metastable ;
	reg \mchip.my_chip.async2sync6.sync ;
	wire [6:0] \mchip.my_chip.btn ;
	wire \mchip.my_chip.clk ;
	wire [6:0] \mchip.my_chip.col ;
	wire [5:0] \mchip.my_chip.game.btn ;
	wire [3:0] \mchip.my_chip.game.buttondetector.btn ;
	wire \mchip.my_chip.game.buttondetector.clk ;
	wire [6:0] \mchip.my_chip.game.buttondetector.col ;
	reg \mchip.my_chip.game.buttondetector.game_over ;
	wire [7:0] \mchip.my_chip.game.buttondetector.mask ;
	reg [3:0] \mchip.my_chip.game.buttondetector.press_reg ;
	wire [2:0] \mchip.my_chip.game.buttondetector.row ;
	wire \mchip.my_chip.game.buttondetector.rst_n ;
	wire [3:0] \mchip.my_chip.game.buttondetector.tiles ;
	wire \mchip.my_chip.game.clk ;
	wire [6:0] \mchip.my_chip.game.col ;
	reg [11:0] \mchip.my_chip.game.count ;
	wire [11:0] \mchip.my_chip.game.count_end ;
	wire \mchip.my_chip.game.dc ;
	wire [63:0] \mchip.my_chip.game.displaytext.a ;
	wire \mchip.my_chip.game.displaytext.clk ;
	wire [6:0] \mchip.my_chip.game.displaytext.col ;
	wire [7:0] \mchip.my_chip.game.displaytext.data ;
	wire [63:0] \mchip.my_chip.game.displaytext.e ;
	wire [63:0] \mchip.my_chip.game.displaytext.g ;
	wire \mchip.my_chip.game.displaytext.game_over ;
	wire [63:0] \mchip.my_chip.game.displaytext.l ;
	wire [63:0] \mchip.my_chip.game.displaytext.m ;
	wire [63:0] \mchip.my_chip.game.displaytext.o ;
	wire [63:0] \mchip.my_chip.game.displaytext.p ;
	wire [2:0] \mchip.my_chip.game.displaytext.place ;
	wire [63:0] \mchip.my_chip.game.displaytext.r ;
	wire [2:0] \mchip.my_chip.game.displaytext.row ;
	wire \mchip.my_chip.game.displaytext.rst_n ;
	wire [63:0] \mchip.my_chip.game.displaytext.v ;
	wire [63:0] \mchip.my_chip.game.displaytext.y ;
	wire \mchip.my_chip.game.displaytiles.clk ;
	wire [6:0] \mchip.my_chip.game.displaytiles.col ;
	wire [7:0] \mchip.my_chip.game.displaytiles.data ;
	wire [7:0] \mchip.my_chip.game.displaytiles.horz_mask ;
	wire [2:0] \mchip.my_chip.game.displaytiles.place ;
	wire [2:0] \mchip.my_chip.game.displaytiles.row ;
	wire \mchip.my_chip.game.displaytiles.rst_n ;
	wire [4:0] \mchip.my_chip.game.displaytiles.tile_loc ;
	wire [19:0] \mchip.my_chip.game.displaytiles.tiles ;
	wire [7:0] \mchip.my_chip.game.displaytiles.vert_mask ;
	wire \mchip.my_chip.game.frame ;
	wire \mchip.my_chip.game.game_over ;
	wire [7:0] \mchip.my_chip.game.mask ;
	wire [3:0] \mchip.my_chip.game.new_tiles ;
	reg \mchip.my_chip.game.pframe ;
	wire [2:0] \mchip.my_chip.game.place ;
	wire \mchip.my_chip.game.random.clk ;
	wire \mchip.my_chip.game.random.next_bit ;
	reg [23:0] \mchip.my_chip.game.random.random_reg ;
	wire \mchip.my_chip.game.random.rst_n ;
	wire [2:0] \mchip.my_chip.game.row ;
	wire \mchip.my_chip.game.rst_n ;
	reg [6:0] \mchip.my_chip.game.state ;
	wire [7:0] \mchip.my_chip.game.text_data ;
	wire [7:0] \mchip.my_chip.game.tile_data ;
	wire [19:0] \mchip.my_chip.game.tiles ;
	wire \mchip.my_chip.game.tilesreg.clk ;
	wire [3:0] \mchip.my_chip.game.tilesreg.new_tiles ;
	wire \mchip.my_chip.game.tilesreg.rst_n ;
	wire [19:0] \mchip.my_chip.game.tilesreg.tiles ;
	wire \mchip.my_chip.oled_clk ;
	wire \mchip.my_chip.oled_cs_n ;
	wire \mchip.my_chip.oled_dc ;
	wire \mchip.my_chip.oled_mosi ;
	wire \mchip.my_chip.oled_res_n ;
	wire [2:0] \mchip.my_chip.place ;
	wire [2:0] \mchip.my_chip.row ;
	wire \mchip.my_chip.rst_n ;
	wire [5:0] \mchip.my_chip.sbtn ;
	wire \mchip.my_chip.spi.clk ;
	reg [6:0] \mchip.my_chip.spi.col ;
	reg [4:0] \mchip.my_chip.spi.count ;
	wire [4:0] \mchip.my_chip.spi.count_end ;
	wire \mchip.my_chip.spi.dc ;
	wire \mchip.my_chip.spi.mosi ;
	wire [31:0] \mchip.my_chip.spi.out_byte ;
	wire [2:0] \mchip.my_chip.spi.place ;
	reg [2:0] \mchip.my_chip.spi.row ;
	wire \mchip.my_chip.spi.rst_n ;
	wire \mchip.my_chip.spi.spi_clk ;
	reg [12:0] \mchip.my_chip.spi.state ;
	wire \mchip.reset ;
	assign _0511_[0] = ~\mchip.my_chip.spi.count [0];
	assign _0053_ = \mchip.my_chip.game.state [1] | \mchip.my_chip.game.state [5];
	assign _0054_ = ~(_0053_ | \mchip.my_chip.game.state [6]);
	assign _0055_ = ~(_0054_ ^ \mchip.my_chip.game.count [10]);
	assign _0056_ = _0055_ | \mchip.my_chip.game.count [11];
	assign _0057_ = ~(\mchip.my_chip.game.count [8] & \mchip.my_chip.game.count [9]);
	assign _0058_ = _0057_ | _0056_;
	assign _0059_ = \mchip.my_chip.game.state [6] | \mchip.my_chip.game.state [1];
	assign _0060_ = ~(_0059_ | _0054_);
	assign _0061_ = _0060_ ^ \mchip.my_chip.game.count [7];
	assign _0062_ = ~(_0061_ & \mchip.my_chip.game.count [6]);
	assign _0063_ = ~(\mchip.my_chip.game.state [6] | \mchip.my_chip.game.state [5]);
	assign _0064_ = _0063_ & ~_0054_;
	assign _0065_ = _0064_ ^ \mchip.my_chip.game.count [5];
	assign _0066_ = ~(_0065_ & \mchip.my_chip.game.count [4]);
	assign _0067_ = ~(_0066_ | _0062_);
	assign _0068_ = \mchip.my_chip.game.count [0] & \mchip.my_chip.game.count [1];
	assign _0069_ = ~(\mchip.my_chip.game.count [2] & \mchip.my_chip.game.count [3]);
	assign _0070_ = _0068_ & ~_0069_;
	assign _0071_ = ~(_0070_ & _0067_);
	assign _0025_ = _0071_ | _0058_;
	assign _0024_ = \mchip.my_chip.async2sync0.sync  & ~_0025_;
	assign _0072_ = ~(\mchip.my_chip.spi.state [5] | \mchip.my_chip.spi.state [8]);
	assign _0073_ = ~(_0072_ ^ \mchip.my_chip.spi.count [4]);
	assign _0074_ = ~\mchip.my_chip.spi.count [2];
	assign _0075_ = ~(\mchip.my_chip.spi.state [7] | \mchip.my_chip.spi.state [11]);
	assign _0076_ = \mchip.my_chip.spi.state [1] | \mchip.my_chip.spi.state [4];
	assign _0077_ = _0075_ & ~_0076_;
	assign _0078_ = _0077_ ^ \mchip.my_chip.spi.count [3];
	assign _0079_ = _0078_ & ~_0074_;
	assign _0080_ = \mchip.my_chip.spi.count [1] & \mchip.my_chip.spi.count [0];
	assign _0081_ = ~(_0080_ & _0079_);
	assign _0082_ = _0081_ | _0073_;
	assign _0020_ = ~(_0082_ & \mchip.my_chip.async2sync0.sync );
	assign _0083_ = \mchip.my_chip.spi.state [9] & ~_0020_;
	assign _0084_ = ~\mchip.my_chip.async2sync0.sync ;
	assign _0085_ = _0082_ | _0084_;
	assign _0086_ = \mchip.my_chip.spi.state [2] & ~_0085_;
	assign _0019_ = _0086_ | _0083_;
	assign _0087_ = \mchip.my_chip.spi.state [5] & ~_0085_;
	assign _0088_ = \mchip.my_chip.spi.col [2] & \mchip.my_chip.spi.col [3];
	assign _0089_ = ~(\mchip.my_chip.spi.col [0] & \mchip.my_chip.spi.col [1]);
	assign _0090_ = _0088_ & ~_0089_;
	assign _0091_ = ~\mchip.my_chip.spi.col [6];
	assign _0092_ = ~(\mchip.my_chip.spi.col [4] & \mchip.my_chip.spi.col [5]);
	assign _0093_ = _0092_ | _0091_;
	assign _0094_ = _0093_ | ~_0090_;
	assign _0095_ = _0094_ | _0082_;
	assign _0096_ = ~(\mchip.my_chip.spi.row [0] & \mchip.my_chip.spi.row [1]);
	assign _0097_ = \mchip.my_chip.spi.row [2] & ~_0096_;
	assign _0098_ = _0095_ | ~_0097_;
	assign _0099_ = _0098_ | _0082_;
	assign _0100_ = ~(_0099_ & \mchip.my_chip.async2sync0.sync );
	assign _0101_ = \mchip.my_chip.spi.state [3] & ~_0100_;
	assign _0013_ = _0101_ | _0087_;
	assign _0042_ = \mchip.my_chip.spi.state [3] & ~_0095_;
	assign _0102_ = \mchip.my_chip.spi.state [3] & ~_0099_;
	assign _0103_ = _0042_ | _0084_;
	assign _0021_ = _0103_ | _0102_;
	assign _0104_ = \mchip.my_chip.spi.state [1] & ~_0085_;
	assign _0105_ = \mchip.my_chip.spi.state [4] & ~_0020_;
	assign _0014_ = _0105_ | _0104_;
	assign _0106_ = \mchip.my_chip.spi.state [8] & ~_0085_;
	assign _0107_ = \mchip.my_chip.spi.state [5] & ~_0020_;
	assign _0015_ = _0107_ | _0106_;
	assign _0022_ = _0102_ | _0084_;
	assign _0108_ = \mchip.my_chip.spi.state [9] & ~_0085_;
	assign _0109_ = \mchip.my_chip.spi.state [6] & ~_0020_;
	assign _0016_ = _0109_ | _0108_;
	assign _0110_ = \mchip.my_chip.spi.state [0] & ~_0085_;
	assign _0111_ = \mchip.my_chip.spi.state [7] & ~_0020_;
	assign _0017_ = _0111_ | _0110_;
	assign _0112_ = \mchip.my_chip.spi.state [12] & ~_0085_;
	assign _0113_ = \mchip.my_chip.spi.state [8] & ~_0020_;
	assign _0114_ = _0099_ | _0084_;
	assign _0115_ = \mchip.my_chip.spi.state [3] & ~_0114_;
	assign _0116_ = _0115_ | _0113_;
	assign _0018_ = _0116_ | _0112_;
	assign _0117_ = \mchip.my_chip.spi.state [2] & ~_0020_;
	assign _0118_ = \mchip.my_chip.spi.state [11] & ~_0085_;
	assign _0012_ = _0118_ | _0117_;
	assign _0119_ = \mchip.my_chip.async2sync6.sync  | \mchip.my_chip.async2sync5.sync ;
	assign _0120_ = _0119_ | \mchip.my_chip.async2sync4.sync ;
	assign _0121_ = _0120_ | \mchip.my_chip.async2sync3.sync ;
	assign _0122_ = _0121_ | \mchip.my_chip.async2sync2.sync ;
	assign _0123_ = _0122_ | _0084_;
	assign _0124_ = \mchip.my_chip.game.state [0] & ~_0123_;
	assign _0125_ = _0051_ & \mchip.my_chip.async2sync0.sync ;
	assign _0126_ = _0050_ & \mchip.my_chip.async2sync0.sync ;
	assign _0127_ = _0126_ & _0125_;
	assign _0128_ = _0052_ & \mchip.my_chip.async2sync0.sync ;
	assign _0129_ = _0128_ & _0127_;
	assign _0130_ = ~(_0129_ & \mchip.my_chip.async2sync0.sync );
	assign _0131_ = \mchip.my_chip.game.state [3] & ~_0130_;
	assign _0132_ = _0131_ | _0084_;
	assign _0001_ = _0132_ | _0124_;
	assign _0023_ = ~(_0025_ & \mchip.my_chip.async2sync0.sync );
	assign _0133_ = \mchip.my_chip.game.buttondetector.game_over  | ~\mchip.my_chip.async2sync0.sync ;
	assign _0134_ = _0049_ & \mchip.my_chip.async2sync0.sync ;
	assign _0135_ = _0048_ & \mchip.my_chip.async2sync0.sync ;
	assign _0136_ = _0047_ & \mchip.my_chip.async2sync0.sync ;
	assign _0137_ = _0046_ & \mchip.my_chip.async2sync0.sync ;
	assign _0138_ = _0045_ & \mchip.my_chip.async2sync0.sync ;
	assign _0139_ = ~(_0135_ | _0134_);
	assign _0140_ = _0133_ | ~_0139_;
	assign _0141_ = \mchip.my_chip.game.state [1] & ~_0140_;
	assign _0142_ = ~_0134_;
	assign _0143_ = _0135_ & ~_0136_;
	assign _0144_ = _0138_ & _0137_;
	assign _0145_ = _0143_ & ~_0144_;
	assign _0146_ = _0135_ & ~_0145_;
	assign _0147_ = _0142_ & ~_0146_;
	assign _0148_ = _0137_ & ~_0138_;
	assign _0149_ = ~(_0148_ & _0143_);
	assign _0150_ = _0142_ & ~_0149_;
	assign _0151_ = _0147_ & ~_0150_;
	assign _0152_ = _0151_ | _0133_;
	assign _0153_ = \mchip.my_chip.game.state [6] & ~_0152_;
	assign _0002_ = _0153_ | _0141_;
	assign _0154_ = \mchip.my_chip.game.buttondetector.game_over  & \mchip.my_chip.async2sync0.sync ;
	assign _0155_ = _0154_ & ~_0054_;
	assign _0156_ = _0129_ | _0084_;
	assign _0157_ = \mchip.my_chip.game.state [3] & ~_0156_;
	assign _0004_ = _0157_ | _0155_;
	assign _0158_ = \mchip.my_chip.spi.state [12] & ~_0020_;
	assign _0159_ = \mchip.my_chip.spi.state [6] & ~_0085_;
	assign _0010_ = _0159_ | _0158_;
	assign _0160_ = \mchip.my_chip.spi.state [4] & ~_0085_;
	assign _0161_ = \mchip.my_chip.spi.state [11] & ~_0020_;
	assign _0009_ = _0161_ | _0160_;
	assign _0162_ = ~(_0122_ | _0025_);
	assign _0163_ = ~(_0162_ & \mchip.my_chip.async2sync0.sync );
	assign _0164_ = \mchip.my_chip.game.state [4] & ~_0163_;
	assign _0165_ = \mchip.my_chip.game.state [2] & ~_0023_;
	assign _0003_ = _0165_ | _0164_;
	assign _0166_ = \mchip.my_chip.game.tilesreg.tiles [15] ^ \mchip.my_chip.game.buttondetector.press_reg [3];
	assign _0167_ = \mchip.my_chip.game.tilesreg.tiles [14] ^ \mchip.my_chip.game.buttondetector.press_reg [2];
	assign _0168_ = _0167_ | _0166_;
	assign _0169_ = \mchip.my_chip.game.tilesreg.tiles [13] ^ \mchip.my_chip.game.buttondetector.press_reg [1];
	assign _0170_ = \mchip.my_chip.game.tilesreg.tiles [12] ^ \mchip.my_chip.game.buttondetector.press_reg [0];
	assign _0171_ = _0170_ | _0169_;
	assign _0026_ = _0171_ | _0168_;
	assign \mchip.my_chip.game.displaytiles.horz_mask [7] = ~\mchip.my_chip.spi.row [0];
	assign _0172_ = \mchip.my_chip.spi.state [1] & ~_0020_;
	assign _0173_ = \mchip.my_chip.spi.state [7] & ~_0085_;
	assign _0011_ = _0173_ | _0172_;
	assign _0174_ = \mchip.my_chip.spi.state [0] & ~_0020_;
	assign _0008_ = _0174_ | _0084_;
	assign _0509_[0] = ~\mchip.my_chip.game.count [0];
	assign _0514_[0] = ~\mchip.my_chip.spi.col [0];
	assign _0175_ = _0133_ | ~_0151_;
	assign _0176_ = \mchip.my_chip.game.state [6] & ~_0175_;
	assign _0177_ = _0024_ & \mchip.my_chip.game.state [2];
	assign _0007_ = _0177_ | _0176_;
	assign _0178_ = _0139_ | _0133_;
	assign _0179_ = \mchip.my_chip.game.state [1] & ~_0178_;
	assign _0180_ = \mchip.my_chip.game.state [5] & ~_0133_;
	assign _0006_ = _0180_ | _0179_;
	assign _0181_ = _0162_ | _0084_;
	assign _0182_ = \mchip.my_chip.game.state [4] & ~_0181_;
	assign _0183_ = ~(_0122_ & \mchip.my_chip.async2sync0.sync );
	assign _0184_ = \mchip.my_chip.game.state [0] & ~_0183_;
	assign _0005_ = _0184_ | _0182_;
	assign _0185_ = _0080_ & ~_0074_;
	assign _0186_ = _0094_ | ~_0097_;
	assign \mchip.my_chip.game.frame  = _0185_ & ~_0186_;
	assign _0043_ = \mchip.my_chip.spi.state [3] & ~_0082_;
	assign _0030_ = ~(_0138_ | _0054_);
	assign _0187_ = _0138_ ^ _0137_;
	assign _0031_ = _0187_ & ~_0054_;
	assign _0188_ = ~_0054_;
	assign _0189_ = ~_0136_;
	assign _0190_ = _0144_ ^ _0189_;
	assign _0032_ = _0188_ & ~_0190_;
	assign _0191_ = ~(_0144_ & _0136_);
	assign _0192_ = _0191_ ^ _0135_;
	assign _0033_ = _0188_ & ~_0192_;
	assign _0193_ = ~(_0136_ & _0135_);
	assign _0194_ = _0144_ & ~_0193_;
	assign _0195_ = _0194_ ^ _0142_;
	assign _0034_ = _0188_ & ~_0195_;
	assign _0027_ = \mchip.my_chip.game.state [3] & ~_0126_;
	assign _0196_ = ~(_0126_ ^ _0125_);
	assign _0028_ = \mchip.my_chip.game.state [3] & ~_0196_;
	assign _0197_ = ~(_0128_ ^ _0127_);
	assign _0029_ = \mchip.my_chip.game.state [3] & ~_0197_;
	assign _0198_ = \mchip.my_chip.game.random.random_reg [3] ^ \mchip.my_chip.game.random.random_reg [1];
	assign _0199_ = ~(\mchip.my_chip.game.random.random_reg [14] ^ \mchip.my_chip.game.random.random_reg [11]);
	assign _0200_ = _0198_ & ~_0199_;
	assign _0201_ = ~(_0059_ | \mchip.my_chip.game.state [5]);
	assign \mchip.my_chip.game.tilesreg.new_tiles [0] = _0200_ & ~_0201_;
	assign _0202_ = ~(\mchip.my_chip.game.random.random_reg [12] ^ \mchip.my_chip.game.random.random_reg [13]);
	assign _0203_ = ~(\mchip.my_chip.game.random.random_reg [7] ^ \mchip.my_chip.game.random.random_reg [2]);
	assign _0204_ = ~(_0203_ | _0202_);
	assign \mchip.my_chip.game.tilesreg.new_tiles [1] = _0204_ & ~_0201_;
	assign _0205_ = ~(\mchip.my_chip.game.random.random_reg [10] ^ \mchip.my_chip.game.random.random_reg [15]);
	assign _0206_ = ~(\mchip.my_chip.game.random.random_reg [4] ^ \mchip.my_chip.game.random.random_reg [5]);
	assign _0207_ = ~(_0206_ | _0205_);
	assign \mchip.my_chip.game.tilesreg.new_tiles [2] = _0207_ & ~_0201_;
	assign _0208_ = ~(\mchip.my_chip.game.random.random_reg [6] ^ \mchip.my_chip.game.random.random_reg [9]);
	assign _0209_ = ~(\mchip.my_chip.game.random.random_reg [0] ^ \mchip.my_chip.game.random.random_reg [8]);
	assign _0210_ = ~(_0209_ | _0208_);
	assign \mchip.my_chip.game.tilesreg.new_tiles [3] = _0210_ & ~_0201_;
	assign _0211_ = _0044_ & \mchip.my_chip.async2sync0.sync ;
	assign _0040_ = ~_0211_;
	assign \mchip.my_chip.async2sync6.async  = ~io_in[13];
	assign _0000_ = \mchip.my_chip.spi.state [10] & \mchip.my_chip.async2sync0.sync ;
	assign _0036_ = \mchip.my_chip.async2sync1.sync  | \mchip.my_chip.game.buttondetector.press_reg [0];
	assign _0037_ = \mchip.my_chip.game.buttondetector.press_reg [1] | \mchip.my_chip.async2sync2.sync ;
	assign _0038_ = \mchip.my_chip.game.buttondetector.press_reg [2] | \mchip.my_chip.async2sync4.sync ;
	assign _0039_ = \mchip.my_chip.game.buttondetector.press_reg [3] | \mchip.my_chip.async2sync6.sync ;
	assign _0212_ = \mchip.my_chip.game.random.random_reg [23] ^ \mchip.my_chip.game.random.random_reg [22];
	assign _0213_ = _0212_ ^ \mchip.my_chip.game.random.random_reg [21];
	assign _0214_ = _0213_ ^ \mchip.my_chip.game.random.random_reg [16];
	assign \mchip.my_chip.game.random.next_bit  = _0214_ ^ \mchip.my_chip.game.random.random_reg [0];
	assign _0215_ = \mchip.my_chip.async2sync1.sync  ^ \mchip.my_chip.async2sync2.sync ;
	assign _0216_ = _0215_ ^ \mchip.my_chip.async2sync4.sync ;
	assign _0217_ = ~(_0216_ ^ \mchip.my_chip.async2sync5.sync );
	assign _0218_ = _0217_ ^ \mchip.my_chip.async2sync6.sync ;
	assign _0219_ = ~(_0218_ | _0025_);
	assign _0041_ = _0219_ ^ \mchip.my_chip.game.random.random_reg [23];
	assign _0035_ = \mchip.my_chip.game.frame  & ~\mchip.my_chip.game.pframe ;
	assign _0220_ = ~\mchip.my_chip.spi.count [1];
	assign _0221_ = ~_0072_;
	assign _0222_ = \mchip.my_chip.spi.state [10] | \mchip.my_chip.spi.state [3];
	assign _0223_ = _0072_ & ~_0222_;
	assign _0224_ = \mchip.my_chip.spi.state [9] | \mchip.my_chip.spi.state [2];
	assign _0225_ = \mchip.my_chip.spi.state [12] | \mchip.my_chip.spi.state [6];
	assign _0226_ = _0225_ | _0224_;
	assign _0227_ = _0223_ & ~_0226_;
	assign _0228_ = \mchip.my_chip.spi.state [7] | \mchip.my_chip.spi.state [1];
	assign _0229_ = \mchip.my_chip.spi.state [11] | \mchip.my_chip.spi.state [4];
	assign _0230_ = _0229_ | _0228_;
	assign _0231_ = _0230_ | \mchip.my_chip.spi.state [0];
	assign _0232_ = _0227_ & ~_0231_;
	assign _0233_ = _0232_ | ~_0221_;
	assign _0234_ = _0233_ | \mchip.my_chip.spi.count [0];
	assign _0235_ = (\mchip.my_chip.spi.count [0] ? \mchip.my_chip.spi.state [5] : \mchip.my_chip.spi.state [8]);
	assign _0236_ = _0232_ | ~_0235_;
	assign _0237_ = (\mchip.my_chip.spi.count [2] ? _0236_ : _0234_);
	assign _0238_ = _0237_ | _0220_;
	assign _0239_ = _0078_ & ~_0238_;
	assign _0240_ = ~(_0077_ & \mchip.my_chip.spi.count [3]);
	assign _0241_ = _0072_ ^ \mchip.my_chip.spi.count [4];
	assign _0242_ = _0241_ ^ _0240_;
	assign _0243_ = ~\mchip.my_chip.spi.row [2];
	assign _0244_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.tilesreg.tiles [1] : \mchip.my_chip.game.tilesreg.tiles [0]);
	assign _0245_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.tilesreg.tiles [3] : \mchip.my_chip.game.tilesreg.tiles [2]);
	assign _0246_ = (\mchip.my_chip.spi.row [2] ? _0245_ : _0244_);
	assign _0247_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.tilesreg.tiles [5] : \mchip.my_chip.game.tilesreg.tiles [4]);
	assign _0248_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.tilesreg.tiles [7] : \mchip.my_chip.game.tilesreg.tiles [6]);
	assign _0249_ = (\mchip.my_chip.spi.row [2] ? _0248_ : _0247_);
	assign _0250_ = (\mchip.my_chip.spi.col [5] ? _0249_ : _0246_);
	assign _0251_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.tilesreg.tiles [9] : \mchip.my_chip.game.tilesreg.tiles [8]);
	assign _0252_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.tilesreg.tiles [11] : \mchip.my_chip.game.tilesreg.tiles [10]);
	assign _0253_ = (\mchip.my_chip.spi.row [2] ? _0252_ : _0251_);
	assign _0254_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.tilesreg.tiles [13] : \mchip.my_chip.game.tilesreg.tiles [12]);
	assign _0255_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.tilesreg.tiles [15] : \mchip.my_chip.game.tilesreg.tiles [14]);
	assign _0256_ = (\mchip.my_chip.spi.row [2] ? _0255_ : _0254_);
	assign _0257_ = (\mchip.my_chip.spi.col [5] ? _0256_ : _0253_);
	assign _0258_ = (\mchip.my_chip.spi.col [6] ? _0257_ : _0250_);
	assign _0259_ = ~_0258_;
	assign _0260_ = ~(\mchip.my_chip.spi.col [2] | \mchip.my_chip.spi.col [3]);
	assign _0261_ = \mchip.my_chip.spi.col [0] | \mchip.my_chip.spi.col [1];
	assign _0262_ = _0260_ & ~_0261_;
	assign _0263_ = \mchip.my_chip.spi.col [4] | ~\mchip.my_chip.spi.col [5];
	assign _0264_ = _0263_ | _0091_;
	assign _0265_ = _0262_ & ~_0264_;
	assign _0266_ = \mchip.my_chip.spi.col [5] | ~\mchip.my_chip.spi.col [4];
	assign _0267_ = _0266_ | _0091_;
	assign _0268_ = _0090_ & ~_0267_;
	assign _0269_ = \mchip.my_chip.spi.col [4] | \mchip.my_chip.spi.col [5];
	assign _0270_ = _0269_ | _0091_;
	assign _0271_ = _0262_ & ~_0270_;
	assign _0272_ = _0092_ | \mchip.my_chip.spi.col [6];
	assign _0273_ = _0090_ & ~_0272_;
	assign _0274_ = _0263_ | \mchip.my_chip.spi.col [6];
	assign _0275_ = _0262_ & ~_0274_;
	assign _0276_ = _0266_ | \mchip.my_chip.spi.col [6];
	assign _0277_ = _0090_ & ~_0276_;
	assign _0278_ = _0269_ | \mchip.my_chip.spi.col [6];
	assign _0279_ = _0262_ & ~_0278_;
	assign _0280_ = _0279_ | _0277_;
	assign _0281_ = _0280_ | _0275_;
	assign _0282_ = _0281_ | _0273_;
	assign _0283_ = _0282_ | _0271_;
	assign _0284_ = _0283_ | _0268_;
	assign _0285_ = _0284_ | _0265_;
	assign _0286_ = _0285_ | ~_0094_;
	assign _0287_ = _0286_ | \mchip.my_chip.spi.row [0];
	assign _0288_ = _0287_ | _0259_;
	assign _0289_ = _0288_ | ~_0188_;
	assign _0290_ = \mchip.my_chip.spi.state [3] & ~_0289_;
	assign _0291_ = _0290_ | \mchip.my_chip.spi.state [10];
	assign _0292_ = _0291_ | \mchip.my_chip.spi.state [8];
	assign _0293_ = _0292_ | _0226_;
	assign _0294_ = ~(_0293_ | _0229_);
	assign _0295_ = ~(_0294_ | _0232_);
	assign _0296_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.buttondetector.press_reg [1] : \mchip.my_chip.game.buttondetector.press_reg [0]);
	assign _0297_ = (\mchip.my_chip.spi.row [1] ? \mchip.my_chip.game.buttondetector.press_reg [3] : \mchip.my_chip.game.buttondetector.press_reg [2]);
	assign _0298_ = (\mchip.my_chip.spi.row [2] ? _0297_ : _0296_);
	assign _0299_ = \mchip.my_chip.spi.col [5] & \mchip.my_chip.spi.col [6];
	assign _0300_ = ~(_0299_ & _0298_);
	assign _0301_ = _0286_ | _0259_;
	assign _0302_ = ~(_0301_ ^ _0300_);
	assign _0303_ = _0302_ | _0054_;
	assign _0304_ = ~\mchip.my_chip.game.state [3];
	assign _0305_ = \mchip.my_chip.spi.row [0] | ~\mchip.my_chip.spi.row [1];
	assign _0306_ = \mchip.my_chip.spi.row [2] & ~_0305_;
	assign _0307_ = ~(_0211_ ^ \mchip.my_chip.spi.col [3]);
	assign _0308_ = \mchip.my_chip.spi.row [0] | \mchip.my_chip.spi.row [1];
	assign _0309_ = \mchip.my_chip.spi.row [2] & ~_0308_;
	assign _0310_ = _0096_ | \mchip.my_chip.spi.row [2];
	assign _0311_ = _0305_ | \mchip.my_chip.spi.row [2];
	assign _0312_ = _0307_ | \mchip.my_chip.spi.col [2];
	assign _0313_ = _0312_ | _0311_;
	assign _0314_ = _0313_ | ~_0310_;
	assign _0315_ = _0314_ | _0309_;
	assign _0316_ = \mchip.my_chip.spi.row [1] | ~\mchip.my_chip.spi.row [0];
	assign _0317_ = \mchip.my_chip.spi.row [2] & ~_0316_;
	assign _0318_ = (_0317_ ? _0307_ : _0315_);
	assign _0319_ = _0318_ | _0306_;
	assign _0320_ = _0319_ | _0097_;
	assign _0321_ = _0320_ | _0304_;
	assign _0322_ = \mchip.my_chip.game.state [2] | \mchip.my_chip.game.state [0];
	assign _0323_ = \mchip.my_chip.game.state [4] | \mchip.my_chip.game.state [3];
	assign _0324_ = _0323_ | _0322_;
	assign _0325_ = _0321_ | ~_0324_;
	assign _0326_ = _0325_ & _0303_;
	assign _0327_ = _0054_ & ~_0324_;
	assign _0328_ = _0327_ | _0326_;
	assign _0329_ = \mchip.my_chip.spi.state [3] & ~_0328_;
	assign _0330_ = _0329_ | \mchip.my_chip.spi.state [10];
	assign _0331_ = _0330_ | _0221_;
	assign _0332_ = _0331_ | \mchip.my_chip.spi.state [9];
	assign _0333_ = _0332_ | _0229_;
	assign _0334_ = _0333_ | _0232_;
	assign _0335_ = (\mchip.my_chip.spi.count [0] ? _0334_ : _0295_);
	assign _0336_ = _0225_ | \mchip.my_chip.spi.state [2];
	assign _0337_ = ~\mchip.my_chip.spi.col [2];
	assign _0338_ = _0337_ & ~_0261_;
	assign _0339_ = _0338_ | _0307_;
	assign _0340_ = (_0310_ ? _0313_ : _0339_);
	assign _0341_ = (_0309_ ? _0307_ : _0340_);
	assign _0342_ = (_0317_ ? _0307_ : _0341_);
	assign _0343_ = (\mchip.my_chip.spi.col [2] ? _0089_ : _0261_);
	assign _0344_ = _0307_ | ~_0343_;
	assign _0345_ = _0308_ | \mchip.my_chip.spi.row [2];
	assign _0346_ = _0345_ | _0307_;
	assign _0347_ = _0243_ & ~_0316_;
	assign _0348_ = (_0347_ ? _0307_ : _0346_);
	assign _0349_ = ~(_0089_ & \mchip.my_chip.spi.col [2]);
	assign _0350_ = _0349_ | _0307_;
	assign _0351_ = (_0311_ ? _0348_ : _0350_);
	assign _0352_ = (_0310_ ? _0351_ : _0344_);
	assign _0353_ = (_0309_ ? _0307_ : _0352_);
	assign _0354_ = ~(\mchip.my_chip.spi.col [0] | \mchip.my_chip.spi.col [1]);
	assign _0515_[1] = _0089_ & ~_0354_;
	assign _0355_ = ~(_0515_[1] & _0337_);
	assign _0356_ = _0355_ | _0307_;
	assign _0357_ = (_0317_ ? _0356_ : _0353_);
	assign _0358_ = (_0306_ ? _0339_ : _0357_);
	assign _0359_ = (_0097_ ? _0344_ : _0358_);
	assign _0360_ = (\mchip.my_chip.game.state [3] ? _0359_ : _0342_);
	assign _0361_ = _0360_ | ~_0324_;
	assign _0362_ = _0188_ & ~_0301_;
	assign _0363_ = _0361_ & ~_0362_;
	assign _0364_ = _0363_ | _0327_;
	assign _0365_ = \mchip.my_chip.spi.state [3] & ~_0364_;
	assign _0366_ = _0365_ | \mchip.my_chip.spi.state [10];
	assign _0367_ = _0366_ | _0221_;
	assign _0368_ = ~(_0367_ | _0336_);
	assign _0369_ = _0368_ & ~\mchip.my_chip.spi.state [11];
	assign _0370_ = ~(_0369_ | _0232_);
	assign _0371_ = _0307_ | _0261_;
	assign _0372_ = _0515_[1] | _0337_;
	assign _0373_ = _0372_ | _0307_;
	assign _0374_ = _0373_ | _0311_;
	assign _0375_ = (_0310_ ? _0374_ : _0371_);
	assign _0376_ = _0089_ | _0337_;
	assign _0377_ = _0376_ | _0307_;
	assign _0378_ = (_0309_ ? _0377_ : _0375_);
	assign _0379_ = (_0317_ ? _0371_ : _0378_);
	assign _0380_ = _0343_ | _0307_;
	assign _0381_ = (\mchip.my_chip.spi.col [2] ? _0515_[1] : _0261_);
	assign _0382_ = _0381_ | _0307_;
	assign _0383_ = _0371_ | _0345_;
	assign _0384_ = (_0347_ ? _0382_ : _0383_);
	assign _0385_ = (_0311_ ? _0384_ : _0377_);
	assign _0386_ = (_0310_ ? _0385_ : _0380_);
	assign _0387_ = (_0309_ ? _0382_ : _0386_);
	assign _0388_ = (\mchip.my_chip.spi.col [2] ? _0261_ : _0089_);
	assign _0389_ = _0388_ | _0307_;
	assign _0390_ = (_0317_ ? _0389_ : _0387_);
	assign _0391_ = (_0306_ ? _0371_ : _0390_);
	assign _0392_ = (_0097_ ? _0380_ : _0391_);
	assign _0393_ = (\mchip.my_chip.game.state [3] ? _0392_ : _0379_);
	assign _0394_ = _0324_ & ~_0393_;
	assign _0395_ = _0303_ & ~_0394_;
	assign _0396_ = _0395_ | _0327_;
	assign _0397_ = \mchip.my_chip.spi.state [3] & ~_0396_;
	assign _0398_ = _0397_ | \mchip.my_chip.spi.state [10];
	assign _0399_ = ~(_0398_ | _0221_);
	assign _0400_ = ~(_0399_ & _0075_);
	assign _0401_ = _0400_ | _0232_;
	assign _0402_ = (\mchip.my_chip.spi.count [0] ? _0401_ : _0370_);
	assign _0403_ = (\mchip.my_chip.spi.count [1] ? _0402_ : _0335_);
	assign _0404_ = \mchip.my_chip.spi.state [12] | \mchip.my_chip.spi.state [9];
	assign _0405_ = _0307_ | _0337_;
	assign _0406_ = _0405_ | _0311_;
	assign _0407_ = (_0310_ ? _0406_ : _0371_);
	assign _0408_ = (_0309_ ? _0377_ : _0407_);
	assign _0409_ = (_0317_ ? _0371_ : _0408_);
	assign _0410_ = (_0097_ ? _0382_ : _0391_);
	assign _0411_ = (\mchip.my_chip.game.state [3] ? _0410_ : _0409_);
	assign _0412_ = _0324_ & ~_0411_;
	assign _0413_ = ~(_0412_ | _0362_);
	assign _0414_ = _0413_ | _0327_;
	assign _0415_ = \mchip.my_chip.spi.state [3] & ~_0414_;
	assign _0416_ = _0415_ | \mchip.my_chip.spi.state [10];
	assign _0417_ = _0416_ | _0221_;
	assign _0418_ = ~(_0417_ | _0404_);
	assign _0419_ = _0418_ & ~\mchip.my_chip.spi.state [4];
	assign _0420_ = (_0309_ ? _0377_ : _0340_);
	assign _0421_ = _0354_ | \mchip.my_chip.spi.col [2];
	assign _0422_ = _0421_ | _0307_;
	assign _0423_ = (_0317_ ? _0422_ : _0420_);
	assign _0424_ = _0307_ | _0354_;
	assign _0425_ = _0424_ | _0345_;
	assign _0426_ = (_0347_ ? _0380_ : _0425_);
	assign _0427_ = (_0311_ ? _0426_ : _0350_);
	assign _0428_ = (_0310_ ? _0427_ : _0344_);
	assign _0429_ = (_0309_ ? _0380_ : _0428_);
	assign _0430_ = (_0317_ ? _0356_ : _0429_);
	assign _0431_ = (_0306_ ? _0339_ : _0430_);
	assign _0432_ = (\mchip.my_chip.spi.col [2] ? _0089_ : _0515_[1]);
	assign _0433_ = _0307_ | ~_0432_;
	assign _0434_ = (_0097_ ? _0433_ : _0431_);
	assign _0435_ = (\mchip.my_chip.game.state [3] ? _0434_ : _0423_);
	assign _0436_ = _0324_ & ~_0435_;
	assign _0437_ = _0303_ & ~_0436_;
	assign _0438_ = _0437_ | _0327_;
	assign _0439_ = \mchip.my_chip.spi.state [3] & ~_0438_;
	assign _0440_ = _0439_ | \mchip.my_chip.spi.state [10];
	assign _0441_ = _0440_ | _0221_;
	assign _0442_ = ~(_0441_ | _0225_);
	assign _0443_ = \mchip.my_chip.spi.state [7] | \mchip.my_chip.spi.state [4];
	assign _0444_ = _0442_ & ~_0443_;
	assign _0445_ = (\mchip.my_chip.spi.count [0] ? _0444_ : _0419_);
	assign _0446_ = ~(_0445_ | _0232_);
	assign _0447_ = _0325_ & ~_0362_;
	assign _0448_ = _0447_ | _0327_;
	assign _0449_ = \mchip.my_chip.spi.state [3] & ~_0448_;
	assign _0450_ = _0449_ | \mchip.my_chip.spi.state [10];
	assign _0451_ = _0450_ | _0221_;
	assign _0452_ = _0451_ | \mchip.my_chip.spi.state [12];
	assign _0453_ = _0452_ | \mchip.my_chip.spi.state [4];
	assign _0454_ = \mchip.my_chip.spi.state [12] | \mchip.my_chip.spi.state [2];
	assign _0455_ = _0286_ | \mchip.my_chip.game.displaytiles.horz_mask [7];
	assign _0456_ = _0258_ & ~_0455_;
	assign _0457_ = _0456_ ^ _0300_;
	assign _0458_ = _0457_ | _0054_;
	assign _0459_ = _0458_ | _0327_;
	assign _0460_ = \mchip.my_chip.spi.state [3] & ~_0459_;
	assign _0461_ = _0460_ | \mchip.my_chip.spi.state [10];
	assign _0462_ = _0461_ | _0221_;
	assign _0463_ = _0462_ | _0454_;
	assign _0464_ = _0463_ | _0229_;
	assign _0465_ = (\mchip.my_chip.spi.count [0] ? _0464_ : _0453_);
	assign _0466_ = _0465_ | _0232_;
	assign _0467_ = (\mchip.my_chip.spi.count [1] ? _0466_ : _0446_);
	assign _0468_ = (\mchip.my_chip.spi.count [2] ? _0467_ : _0403_);
	assign _0469_ = ~\mchip.my_chip.spi.state [7];
	assign _0470_ = _0469_ & ~_0229_;
	assign _0471_ = ~(_0470_ | _0232_);
	assign _0472_ = \mchip.my_chip.spi.state [11] & ~_0232_;
	assign _0473_ = (\mchip.my_chip.spi.count [0] ? _0472_ : _0471_);
	assign _0474_ = \mchip.my_chip.spi.state [1] & ~_0232_;
	assign _0475_ = (\mchip.my_chip.spi.count [0] ? _0472_ : _0474_);
	assign _0476_ = (\mchip.my_chip.spi.count [1] ? _0475_ : _0473_);
	assign _0477_ = (\mchip.my_chip.spi.count [0] ? _0469_ : _0075_);
	assign _0478_ = ~(_0477_ | _0232_);
	assign _0479_ = _0471_ & ~_0511_[0];
	assign _0480_ = (\mchip.my_chip.spi.count [1] ? _0479_ : _0478_);
	assign _0481_ = (\mchip.my_chip.spi.count [2] ? _0480_ : _0476_);
	assign _0482_ = (_0078_ ? _0468_ : _0481_);
	assign _0483_ = (_0242_ ? _0239_ : _0482_);
	assign _0484_ = ~(\mchip.my_chip.spi.state [2] | \mchip.my_chip.spi.state [1]);
	assign _0485_ = \mchip.my_chip.spi.state [3] | \mchip.my_chip.spi.state [4];
	assign _0486_ = _0484_ & ~_0485_;
	assign _0487_ = \mchip.my_chip.spi.state [8] | \mchip.my_chip.spi.state [7];
	assign _0488_ = \mchip.my_chip.spi.state [6] | \mchip.my_chip.spi.state [5];
	assign _0489_ = _0488_ | _0487_;
	assign _0490_ = _0486_ & ~_0489_;
	assign _0491_ = \mchip.my_chip.spi.state [9] | \mchip.my_chip.spi.state [11];
	assign _0492_ = _0491_ | \mchip.my_chip.spi.state [12];
	assign _0493_ = _0490_ & ~_0492_;
	assign \mchip.my_chip.oled_mosi  = _0483_ & ~_0493_;
	assign \mchip.my_chip.oled_clk  = ~(_0493_ | io_in[12]);
	assign _0515_[2] = _0089_ ^ _0337_;
	assign _0515_[3] = ~(_0376_ ^ \mchip.my_chip.spi.col [3]);
	assign _0515_[4] = _0090_ ^ \mchip.my_chip.spi.col [4];
	assign _0494_ = _0090_ & \mchip.my_chip.spi.col [4];
	assign _0515_[5] = _0494_ ^ \mchip.my_chip.spi.col [5];
	assign _0495_ = _0090_ & ~_0092_;
	assign _0515_[6] = _0495_ ^ \mchip.my_chip.spi.col [6];
	assign _0513_[1] = ~(_0316_ & _0305_);
	assign _0513_[2] = _0096_ ^ _0243_;
	assign _0510_[1] = \mchip.my_chip.game.count [0] ^ \mchip.my_chip.game.count [1];
	assign _0510_[2] = _0068_ ^ \mchip.my_chip.game.count [2];
	assign _0496_ = _0068_ & \mchip.my_chip.game.count [2];
	assign _0510_[3] = _0496_ ^ \mchip.my_chip.game.count [3];
	assign _0510_[4] = _0070_ ^ \mchip.my_chip.game.count [4];
	assign _0497_ = _0070_ & \mchip.my_chip.game.count [4];
	assign _0510_[5] = _0497_ ^ \mchip.my_chip.game.count [5];
	assign _0498_ = ~(\mchip.my_chip.game.count [4] & \mchip.my_chip.game.count [5]);
	assign _0499_ = _0070_ & ~_0498_;
	assign _0510_[6] = _0499_ ^ \mchip.my_chip.game.count [6];
	assign _0500_ = _0499_ & \mchip.my_chip.game.count [6];
	assign _0510_[7] = _0500_ ^ \mchip.my_chip.game.count [7];
	assign _0501_ = ~(\mchip.my_chip.game.count [6] & \mchip.my_chip.game.count [7]);
	assign _0502_ = ~(_0501_ | _0498_);
	assign _0503_ = ~(_0502_ & _0070_);
	assign _0510_[8] = ~(_0503_ ^ \mchip.my_chip.game.count [8]);
	assign _0504_ = \mchip.my_chip.game.count [8] & ~_0503_;
	assign _0510_[9] = _0504_ ^ \mchip.my_chip.game.count [9];
	assign _0505_ = ~(_0503_ | _0057_);
	assign _0510_[10] = _0505_ ^ \mchip.my_chip.game.count [10];
	assign _0506_ = _0505_ & \mchip.my_chip.game.count [10];
	assign _0510_[11] = _0506_ ^ \mchip.my_chip.game.count [11];
	assign _0512_[1] = \mchip.my_chip.spi.count [1] ^ \mchip.my_chip.spi.count [0];
	assign _0512_[2] = _0080_ ^ \mchip.my_chip.spi.count [2];
	assign _0512_[3] = _0185_ ^ \mchip.my_chip.spi.count [3];
	assign _0507_ = ~(\mchip.my_chip.spi.count [2] & \mchip.my_chip.spi.count [3]);
	assign _0508_ = _0080_ & ~_0507_;
	assign _0512_[4] = _0508_ ^ \mchip.my_chip.spi.count [4];
	always @(posedge io_in[12]) \mchip.my_chip.game.state [0] <= _0001_;
	always @(posedge io_in[12]) \mchip.my_chip.game.state [1] <= _0002_;
	always @(posedge io_in[12]) \mchip.my_chip.game.state [2] <= _0003_;
	always @(posedge io_in[12]) \mchip.my_chip.game.state [3] <= _0004_;
	always @(posedge io_in[12]) \mchip.my_chip.game.state [4] <= _0005_;
	always @(posedge io_in[12]) \mchip.my_chip.game.state [5] <= _0006_;
	always @(posedge io_in[12]) \mchip.my_chip.game.state [6] <= _0007_;
	always @(posedge io_in[12]) \mchip.my_chip.async2sync1.sync  <= \mchip.my_chip.async2sync1.metastable ;
	always @(posedge io_in[12]) \mchip.my_chip.async2sync2.sync  <= \mchip.my_chip.async2sync2.metastable ;
	always @(posedge io_in[12]) \mchip.my_chip.async2sync3.sync  <= \mchip.my_chip.async2sync3.metastable ;
	always @(posedge io_in[12]) \mchip.my_chip.async2sync4.sync  <= \mchip.my_chip.async2sync4.metastable ;
	always @(posedge io_in[12]) \mchip.my_chip.async2sync5.sync  <= \mchip.my_chip.async2sync5.metastable ;
	always @(posedge io_in[12]) \mchip.my_chip.async2sync6.sync  <= \mchip.my_chip.async2sync6.metastable ;
	always @(posedge io_in[12]) \mchip.my_chip.async2sync0.metastable  <= io_in[0];
	always @(posedge io_in[12]) \mchip.my_chip.async2sync1.metastable  <= io_in[1];
	always @(posedge io_in[12]) \mchip.my_chip.async2sync2.metastable  <= io_in[2];
	always @(posedge io_in[12]) \mchip.my_chip.async2sync3.metastable  <= io_in[3];
	always @(posedge io_in[12]) \mchip.my_chip.async2sync4.metastable  <= io_in[4];
	always @(posedge io_in[12]) \mchip.my_chip.async2sync5.metastable  <= io_in[5];
	always @(posedge io_in[12]) \mchip.my_chip.async2sync6.metastable  <= \mchip.my_chip.async2sync6.async ;
	always @(posedge io_in[12])
		if (!_0024_)
			\mchip.my_chip.game.buttondetector.game_over  <= 1'h0;
		else
			\mchip.my_chip.game.buttondetector.game_over  <= _0026_;
	always @(negedge _0025_)
		if (!\mchip.my_chip.async2sync0.sync )
			_0044_ <= 1'h0;
		else
			_0044_ <= _0040_;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[0] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[0]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[0]  <= \mchip.my_chip.game.tilesreg.new_tiles [0];
	assign \mchip.my_chip.game.tilesreg.tiles [0] = \mchip.my_chip.game.tilesreg.tiles_reg[0] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[1] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[1]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[1]  <= \mchip.my_chip.game.tilesreg.new_tiles [1];
	assign \mchip.my_chip.game.tilesreg.tiles [1] = \mchip.my_chip.game.tilesreg.tiles_reg[1] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[2] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[2]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[2]  <= \mchip.my_chip.game.tilesreg.new_tiles [2];
	assign \mchip.my_chip.game.tilesreg.tiles [2] = \mchip.my_chip.game.tilesreg.tiles_reg[2] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[3] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[3]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[3]  <= \mchip.my_chip.game.tilesreg.new_tiles [3];
	assign \mchip.my_chip.game.tilesreg.tiles [3] = \mchip.my_chip.game.tilesreg.tiles_reg[3] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[4] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[4]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[4]  <= \mchip.my_chip.game.tilesreg.tiles [0];
	assign \mchip.my_chip.game.tilesreg.tiles [4] = \mchip.my_chip.game.tilesreg.tiles_reg[4] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[5] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[5]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[5]  <= \mchip.my_chip.game.tilesreg.tiles [1];
	assign \mchip.my_chip.game.tilesreg.tiles [5] = \mchip.my_chip.game.tilesreg.tiles_reg[5] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[6] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[6]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[6]  <= \mchip.my_chip.game.tilesreg.tiles [2];
	assign \mchip.my_chip.game.tilesreg.tiles [6] = \mchip.my_chip.game.tilesreg.tiles_reg[6] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[7] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[7]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[7]  <= \mchip.my_chip.game.tilesreg.tiles [3];
	assign \mchip.my_chip.game.tilesreg.tiles [7] = \mchip.my_chip.game.tilesreg.tiles_reg[7] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[8] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[8]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[8]  <= \mchip.my_chip.game.tilesreg.tiles [4];
	assign \mchip.my_chip.game.tilesreg.tiles [8] = \mchip.my_chip.game.tilesreg.tiles_reg[8] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[9] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[9]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[9]  <= \mchip.my_chip.game.tilesreg.tiles [5];
	assign \mchip.my_chip.game.tilesreg.tiles [9] = \mchip.my_chip.game.tilesreg.tiles_reg[9] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[10] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[10]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[10]  <= \mchip.my_chip.game.tilesreg.tiles [6];
	assign \mchip.my_chip.game.tilesreg.tiles [10] = \mchip.my_chip.game.tilesreg.tiles_reg[10] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[11] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[11]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[11]  <= \mchip.my_chip.game.tilesreg.tiles [7];
	assign \mchip.my_chip.game.tilesreg.tiles [11] = \mchip.my_chip.game.tilesreg.tiles_reg[11] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[12] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[12]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[12]  <= \mchip.my_chip.game.tilesreg.tiles [8];
	assign \mchip.my_chip.game.tilesreg.tiles [12] = \mchip.my_chip.game.tilesreg.tiles_reg[12] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[13] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[13]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[13]  <= \mchip.my_chip.game.tilesreg.tiles [9];
	assign \mchip.my_chip.game.tilesreg.tiles [13] = \mchip.my_chip.game.tilesreg.tiles_reg[13] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[14] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[14]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[14]  <= \mchip.my_chip.game.tilesreg.tiles [10];
	assign \mchip.my_chip.game.tilesreg.tiles [14] = \mchip.my_chip.game.tilesreg.tiles_reg[14] ;
	reg \mchip.my_chip.game.tilesreg.tiles_reg[15] ;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.tilesreg.tiles_reg[15]  <= 1'h0;
		else if (!_0025_)
			\mchip.my_chip.game.tilesreg.tiles_reg[15]  <= \mchip.my_chip.game.tilesreg.tiles [11];
	assign \mchip.my_chip.game.tilesreg.tiles [15] = \mchip.my_chip.game.tilesreg.tiles_reg[15] ;
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.buttondetector.press_reg [0] <= 1'h0;
		else
			\mchip.my_chip.game.buttondetector.press_reg [0] <= _0036_;
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.buttondetector.press_reg [1] <= 1'h0;
		else
			\mchip.my_chip.game.buttondetector.press_reg [1] <= _0037_;
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.buttondetector.press_reg [2] <= 1'h0;
		else
			\mchip.my_chip.game.buttondetector.press_reg [2] <= _0038_;
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.buttondetector.press_reg [3] <= 1'h0;
		else
			\mchip.my_chip.game.buttondetector.press_reg [3] <= _0039_;
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [0] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [0] <= _0509_[0];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [1] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [1] <= _0510_[1];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [2] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [2] <= _0510_[2];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [3] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [3] <= _0510_[3];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [4] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [4] <= _0510_[4];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [5] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [5] <= _0510_[5];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [6] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [6] <= _0510_[6];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [7] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [7] <= _0510_[7];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [8] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [8] <= _0510_[8];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [9] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [9] <= _0510_[9];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [10] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [10] <= _0510_[10];
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.my_chip.game.count [11] <= 1'h0;
		else if (_0035_)
			\mchip.my_chip.game.count [11] <= _0510_[11];
	always @(posedge io_in[12]) \mchip.my_chip.game.pframe  <= \mchip.my_chip.game.frame ;
	always @(negedge _0025_)
		if (!\mchip.my_chip.async2sync0.sync )
			_0045_ <= 1'h0;
		else
			_0045_ <= _0030_;
	always @(negedge _0025_)
		if (!\mchip.my_chip.async2sync0.sync )
			_0046_ <= 1'h0;
		else
			_0046_ <= _0031_;
	always @(negedge _0025_)
		if (!\mchip.my_chip.async2sync0.sync )
			_0047_ <= 1'h0;
		else
			_0047_ <= _0032_;
	always @(negedge _0025_)
		if (!\mchip.my_chip.async2sync0.sync )
			_0048_ <= 1'h0;
		else
			_0048_ <= _0033_;
	always @(negedge _0025_)
		if (!\mchip.my_chip.async2sync0.sync )
			_0049_ <= 1'h0;
		else
			_0049_ <= _0034_;
	always @(negedge _0025_)
		if (!\mchip.my_chip.async2sync0.sync )
			_0050_ <= 1'h0;
		else
			_0050_ <= _0027_;
	always @(negedge _0025_)
		if (!\mchip.my_chip.async2sync0.sync )
			_0051_ <= 1'h0;
		else
			_0051_ <= _0028_;
	always @(negedge _0025_)
		if (!\mchip.my_chip.async2sync0.sync )
			_0052_ <= 1'h0;
		else
			_0052_ <= _0029_;
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.my_chip.spi.count [0] <= 1'h0;
		else
			\mchip.my_chip.spi.count [0] <= _0511_[0];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.my_chip.spi.count [1] <= 1'h0;
		else
			\mchip.my_chip.spi.count [1] <= _0512_[1];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.my_chip.spi.count [2] <= 1'h0;
		else
			\mchip.my_chip.spi.count [2] <= _0512_[2];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.my_chip.spi.count [3] <= 1'h0;
		else
			\mchip.my_chip.spi.count [3] <= _0512_[3];
	always @(posedge io_in[12])
		if (_0020_)
			\mchip.my_chip.spi.count [4] <= 1'h0;
		else
			\mchip.my_chip.spi.count [4] <= _0512_[4];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [0] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [0] <= \mchip.my_chip.game.random.random_reg [1];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [1] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [1] <= \mchip.my_chip.game.random.random_reg [2];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [2] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [2] <= \mchip.my_chip.game.random.random_reg [3];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [3] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [3] <= \mchip.my_chip.game.random.random_reg [4];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [4] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [4] <= \mchip.my_chip.game.random.random_reg [5];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [5] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [5] <= \mchip.my_chip.game.random.random_reg [6];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [6] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [6] <= \mchip.my_chip.game.random.random_reg [7];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [7] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [7] <= \mchip.my_chip.game.random.random_reg [8];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [8] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [8] <= \mchip.my_chip.game.random.random_reg [9];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [9] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [9] <= \mchip.my_chip.game.random.random_reg [10];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [10] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [10] <= \mchip.my_chip.game.random.random_reg [11];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [11] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [11] <= \mchip.my_chip.game.random.random_reg [12];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [12] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [12] <= \mchip.my_chip.game.random.random_reg [13];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [13] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [13] <= \mchip.my_chip.game.random.random_reg [14];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [14] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [14] <= \mchip.my_chip.game.random.random_reg [15];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [15] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [15] <= \mchip.my_chip.game.random.random_reg [16];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [16] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [16] <= \mchip.my_chip.game.random.random_reg [17];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [17] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [17] <= \mchip.my_chip.game.random.random_reg [18];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [18] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [18] <= \mchip.my_chip.game.random.random_reg [19];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [19] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [19] <= \mchip.my_chip.game.random.random_reg [20];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [20] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [20] <= \mchip.my_chip.game.random.random_reg [21];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [21] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [21] <= \mchip.my_chip.game.random.random_reg [22];
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [22] <= 1'h1;
		else
			\mchip.my_chip.game.random.random_reg [22] <= _0041_;
	always @(posedge io_in[12])
		if (!\mchip.my_chip.async2sync0.sync )
			\mchip.my_chip.game.random.random_reg [23] <= 1'h0;
		else
			\mchip.my_chip.game.random.random_reg [23] <= \mchip.my_chip.game.random.next_bit ;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.my_chip.spi.col [0] <= 1'h0;
		else if (_0043_)
			\mchip.my_chip.spi.col [0] <= _0514_[0];
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.my_chip.spi.col [1] <= 1'h0;
		else if (_0043_)
			\mchip.my_chip.spi.col [1] <= _0515_[1];
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.my_chip.spi.col [2] <= 1'h0;
		else if (_0043_)
			\mchip.my_chip.spi.col [2] <= _0515_[2];
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.my_chip.spi.col [3] <= 1'h0;
		else if (_0043_)
			\mchip.my_chip.spi.col [3] <= _0515_[3];
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.my_chip.spi.col [4] <= 1'h0;
		else if (_0043_)
			\mchip.my_chip.spi.col [4] <= _0515_[4];
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.my_chip.spi.col [5] <= 1'h0;
		else if (_0043_)
			\mchip.my_chip.spi.col [5] <= _0515_[5];
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.my_chip.spi.col [6] <= 1'h0;
		else if (_0043_)
			\mchip.my_chip.spi.col [6] <= _0515_[6];
	always @(posedge io_in[12])
		if (_0022_)
			\mchip.my_chip.spi.row [0] <= 1'h0;
		else if (_0042_)
			\mchip.my_chip.spi.row [0] <= \mchip.my_chip.game.displaytiles.horz_mask [7];
	always @(posedge io_in[12])
		if (_0022_)
			\mchip.my_chip.spi.row [1] <= 1'h0;
		else if (_0042_)
			\mchip.my_chip.spi.row [1] <= _0513_[1];
	always @(posedge io_in[12])
		if (_0022_)
			\mchip.my_chip.spi.row [2] <= 1'h0;
		else if (_0042_)
			\mchip.my_chip.spi.row [2] <= _0513_[2];
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [0] <= _0008_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [1] <= _0011_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [2] <= _0012_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [3] <= _0013_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [4] <= _0014_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [5] <= _0015_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [6] <= _0016_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [7] <= _0017_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [8] <= _0018_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [9] <= _0019_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [10] <= _0000_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [11] <= _0009_;
	always @(posedge io_in[12]) \mchip.my_chip.spi.state [12] <= _0010_;
	always @(posedge io_in[12]) \mchip.my_chip.async2sync0.sync  <= \mchip.my_chip.async2sync0.metastable ;
	assign _0509_[11:1] = \mchip.my_chip.game.count [11:1];
	assign _0510_[0] = _0509_[0];
	assign _0511_[4:1] = \mchip.my_chip.spi.count [4:1];
	assign _0512_[0] = _0511_[0];
	assign _0513_[0] = \mchip.my_chip.game.displaytiles.horz_mask [7];
	assign _0514_[6:1] = \mchip.my_chip.spi.col [6:1];
	assign _0515_[0] = _0514_[0];
	assign io_out = {2'h0, \mchip.my_chip.oled_clk , \mchip.my_chip.oled_mosi , \mchip.my_chip.spi.state [3], \mchip.my_chip.async2sync0.sync , 8'h00};
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.my_chip.oled_clk , \mchip.my_chip.oled_mosi , \mchip.my_chip.spi.state [3], \mchip.my_chip.async2sync0.sync , 8'h00};
	assign \mchip.my_chip.async2sync0.async  = io_in[0];
	assign \mchip.my_chip.async2sync0.clk  = io_in[12];
	assign \mchip.my_chip.async2sync1.async  = io_in[1];
	assign \mchip.my_chip.async2sync1.clk  = io_in[12];
	assign \mchip.my_chip.async2sync2.async  = io_in[2];
	assign \mchip.my_chip.async2sync2.clk  = io_in[12];
	assign \mchip.my_chip.async2sync3.async  = io_in[3];
	assign \mchip.my_chip.async2sync3.clk  = io_in[12];
	assign \mchip.my_chip.async2sync4.async  = io_in[4];
	assign \mchip.my_chip.async2sync4.clk  = io_in[12];
	assign \mchip.my_chip.async2sync5.async  = io_in[5];
	assign \mchip.my_chip.async2sync5.clk  = io_in[12];
	assign \mchip.my_chip.async2sync6.clk  = io_in[12];
	assign \mchip.my_chip.btn  = {\mchip.my_chip.async2sync6.async , io_in[5:0]};
	assign \mchip.my_chip.clk  = io_in[12];
	assign \mchip.my_chip.col  = \mchip.my_chip.spi.col ;
	assign \mchip.my_chip.game.btn  = {\mchip.my_chip.async2sync6.sync , \mchip.my_chip.async2sync5.sync , \mchip.my_chip.async2sync4.sync , \mchip.my_chip.async2sync3.sync , \mchip.my_chip.async2sync2.sync , \mchip.my_chip.async2sync1.sync };
	assign \mchip.my_chip.game.buttondetector.btn  = {\mchip.my_chip.async2sync6.sync , \mchip.my_chip.async2sync4.sync , \mchip.my_chip.async2sync2.sync , \mchip.my_chip.async2sync1.sync };
	assign \mchip.my_chip.game.buttondetector.clk  = io_in[12];
	assign \mchip.my_chip.game.buttondetector.col  = \mchip.my_chip.spi.col ;
	assign \mchip.my_chip.game.buttondetector.mask  = 8'h00;
	assign \mchip.my_chip.game.buttondetector.row  = \mchip.my_chip.spi.row ;
	assign \mchip.my_chip.game.buttondetector.rst_n  = \mchip.my_chip.async2sync0.sync ;
	assign \mchip.my_chip.game.buttondetector.tiles  = \mchip.my_chip.game.tilesreg.tiles [15:12];
	assign \mchip.my_chip.game.clk  = io_in[12];
	assign \mchip.my_chip.game.col  = \mchip.my_chip.spi.col ;
	assign \mchip.my_chip.game.count_end  = 12'h35f;
	assign \mchip.my_chip.game.dc  = \mchip.my_chip.spi.state [3];
	assign \mchip.my_chip.game.displaytext.a  = 64'h2424243c24242418;
	assign \mchip.my_chip.game.displaytext.clk  = io_in[12];
	assign \mchip.my_chip.game.displaytext.col  = \mchip.my_chip.spi.col ;
	assign \mchip.my_chip.game.displaytext.data  = 8'h00;
	assign \mchip.my_chip.game.displaytext.e  = 64'h3c2020382020203c;
	assign \mchip.my_chip.game.displaytext.g  = 64'h1824242c20242418;
	assign \mchip.my_chip.game.displaytext.game_over  = \mchip.my_chip.game.state [3];
	assign \mchip.my_chip.game.displaytext.l  = 64'h3c20202020202020;
	assign \mchip.my_chip.game.displaytext.m  = 64'h4242425a5a666642;
	assign \mchip.my_chip.game.displaytext.o  = 64'h1824242424242418;
	assign \mchip.my_chip.game.displaytext.p  = 64'h2020203824242438;
	assign \mchip.my_chip.game.displaytext.place  = \mchip.my_chip.spi.count [2:0];
	assign \mchip.my_chip.game.displaytext.r  = 64'h2424243824242438;
	assign \mchip.my_chip.game.displaytext.row  = \mchip.my_chip.spi.row ;
	assign \mchip.my_chip.game.displaytext.rst_n  = \mchip.my_chip.async2sync0.sync ;
	assign \mchip.my_chip.game.displaytext.v  = 64'h1824242442424242;
	assign \mchip.my_chip.game.displaytext.y  = 64'h1808081824242424;
	assign \mchip.my_chip.game.displaytiles.clk  = io_in[12];
	assign \mchip.my_chip.game.displaytiles.col  = \mchip.my_chip.spi.col ;
	assign \mchip.my_chip.game.displaytiles.data  = 8'h00;
	assign \mchip.my_chip.game.displaytiles.horz_mask [6:0] = {6'h3f, \mchip.my_chip.spi.row [0]};
	assign \mchip.my_chip.game.displaytiles.place  = \mchip.my_chip.spi.count [2:0];
	assign \mchip.my_chip.game.displaytiles.row  = \mchip.my_chip.spi.row ;
	assign \mchip.my_chip.game.displaytiles.rst_n  = \mchip.my_chip.async2sync0.sync ;
	assign \mchip.my_chip.game.displaytiles.tile_loc  = {1'h0, \mchip.my_chip.spi.col [6:5], \mchip.my_chip.spi.row [2:1]};
	assign \mchip.my_chip.game.displaytiles.tiles  = {4'h0, \mchip.my_chip.game.tilesreg.tiles [15:0]};
	assign \mchip.my_chip.game.displaytiles.vert_mask  = 8'h00;
	assign \mchip.my_chip.game.game_over  = \mchip.my_chip.game.buttondetector.game_over ;
	assign \mchip.my_chip.game.mask  = 8'h00;
	assign \mchip.my_chip.game.new_tiles  = \mchip.my_chip.game.tilesreg.new_tiles ;
	assign \mchip.my_chip.game.place  = \mchip.my_chip.spi.count [2:0];
	assign \mchip.my_chip.game.random.clk  = io_in[12];
	assign \mchip.my_chip.game.random.rst_n  = \mchip.my_chip.async2sync0.sync ;
	assign \mchip.my_chip.game.row  = \mchip.my_chip.spi.row ;
	assign \mchip.my_chip.game.rst_n  = \mchip.my_chip.async2sync0.sync ;
	assign \mchip.my_chip.game.text_data  = 8'h00;
	assign \mchip.my_chip.game.tile_data  = 8'h00;
	assign \mchip.my_chip.game.tiles  = {4'h0, \mchip.my_chip.game.tilesreg.tiles [15:0]};
	assign \mchip.my_chip.game.tilesreg.clk  = io_in[12];
	assign \mchip.my_chip.game.tilesreg.rst_n  = \mchip.my_chip.async2sync0.sync ;
	assign \mchip.my_chip.game.tilesreg.tiles [19:16] = 4'h0;
	assign \mchip.my_chip.oled_cs_n  = 1'h0;
	assign \mchip.my_chip.oled_dc  = \mchip.my_chip.spi.state [3];
	assign \mchip.my_chip.oled_res_n  = \mchip.my_chip.async2sync0.sync ;
	assign \mchip.my_chip.place  = \mchip.my_chip.spi.count [2:0];
	assign \mchip.my_chip.row  = \mchip.my_chip.spi.row ;
	assign \mchip.my_chip.rst_n  = \mchip.my_chip.async2sync0.sync ;
	assign \mchip.my_chip.sbtn  = {\mchip.my_chip.async2sync6.sync , \mchip.my_chip.async2sync5.sync , \mchip.my_chip.async2sync4.sync , \mchip.my_chip.async2sync3.sync , \mchip.my_chip.async2sync2.sync , \mchip.my_chip.async2sync1.sync };
	assign \mchip.my_chip.spi.clk  = io_in[12];
	assign \mchip.my_chip.spi.count_end  = 5'h07;
	assign \mchip.my_chip.spi.dc  = \mchip.my_chip.spi.state [3];
	assign \mchip.my_chip.spi.mosi  = \mchip.my_chip.oled_mosi ;
	assign \mchip.my_chip.spi.out_byte  = 32'd0;
	assign \mchip.my_chip.spi.place  = \mchip.my_chip.spi.count [2:0];
	assign \mchip.my_chip.spi.rst_n  = \mchip.my_chip.async2sync0.sync ;
	assign \mchip.my_chip.spi.spi_clk  = \mchip.my_chip.oled_clk ;
	assign \mchip.reset  = io_in[13];
endmodule
module d16_jaehyun3_bobatc (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire [2:0] _1628_;
	wire [2:0] _1629_;
	wire [2:0] _1630_;
	wire [2:0] _1631_;
	wire [3:0] _1632_;
	wire [2:0] _1633_;
	wire [2:0] _1634_;
	wire [2:0] _1635_;
	wire [2:0] _1636_;
	wire [3:0] _1637_;
	wire [1:0] _1638_;
	wire [1:0] _1639_;
	wire [1:0] _1640_;
	wire [1:0] _1641_;
	wire [2:0] _1642_;
	wire [1:0] _1643_;
	wire [1:0] _1644_;
	wire [1:0] _1645_;
	wire [1:0] _1646_;
	wire [2:0] _1647_;
	wire [3:0] _1648_;
	wire [3:0] _1649_;
	wire [9:0] _1650_;
	wire [9:0] _1651_;
	wire [3:0] _1652_;
	wire [3:0] _1653_;
	wire [9:0] _1654_;
	wire [9:0] _1655_;
	wire [3:0] _1656_;
	wire [3:0] _1657_;
	wire [7:0] _1658_;
	wire [7:0] _1659_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire [15:0] \mchip.top.bobby.all_id ;
	wire [3:0] \mchip.top.bobby.cleared_id_to_lock ;
	wire [3:0] \mchip.top.bobby.cleared_landing_id ;
	wire [3:0] \mchip.top.bobby.cleared_takeoff_id ;
	wire \mchip.top.bobby.clock ;
	reg \mchip.top.bobby.emergency ;
	reg [3:0] \mchip.top.bobby.emergency_id ;
	wire \mchip.top.bobby.emergency_out ;
	wire \mchip.top.bobby.emergency_override ;
	wire [15:0] \mchip.top.bobby.fsm.all_id ;
	wire \mchip.top.bobby.fsm.clock ;
	wire \mchip.top.bobby.fsm.emergency ;
	wire [3:0] \mchip.top.bobby.fsm.emergency_id ;
	wire [1:0] \mchip.top.bobby.fsm.msg_action ;
	wire [2:0] \mchip.top.bobby.fsm.msg_type ;
	wire [3:0] \mchip.top.bobby.fsm.plane_id ;
	wire \mchip.top.bobby.fsm.reset ;
	wire \mchip.top.bobby.fsm.reverse_takeoff_first ;
	wire [9:0] \mchip.top.bobby.fsm.runway ;
	wire [1:0] \mchip.top.bobby.fsm.runway_active ;
	wire \mchip.top.bobby.fsm.set_emergency ;
	reg [7:0] \mchip.top.bobby.fsm.state ;
	reg \mchip.top.bobby.fsm.takeoff_first ;
	wire [7:0] \mchip.top.bobby.fsm.uart_request ;
	wire [15:0] \mchip.top.bobby.id_manager.all_id ;
	wire \mchip.top.bobby.id_manager.clock ;
	wire \mchip.top.bobby.id_manager.reset ;
	reg [15:0] \mchip.top.bobby.id_manager.taken_id ;
	wire \mchip.top.bobby.landing_fifo.clock ;
	reg [3:0] \mchip.top.bobby.landing_fifo.count ;
	wire [3:0] \mchip.top.bobby.landing_fifo.data_in ;
	reg [3:0] \mchip.top.bobby.landing_fifo.data_out ;
	reg [2:0] \mchip.top.bobby.landing_fifo.get_ptr ;
	reg [2:0] \mchip.top.bobby.landing_fifo.put_ptr ;
	reg [31:0] \mchip.top.bobby.landing_fifo.queue ;
	wire \mchip.top.bobby.landing_fifo.reset ;
	wire \mchip.top.bobby.reply_fsm.clock ;
	wire \mchip.top.bobby.reply_fsm.next_state ;
	wire \mchip.top.bobby.reply_fsm.reset ;
	wire \mchip.top.bobby.reply_fsm.send_reply ;
	reg \mchip.top.bobby.reply_fsm.state ;
	wire \mchip.top.bobby.reply_fsm.uart_tx_send ;
	reg [7:0] \mchip.top.bobby.reply_to_send ;
	wire \mchip.top.bobby.reset ;
	wire [9:0] \mchip.top.bobby.runway ;
	wire [1:0] \mchip.top.bobby.runway_active ;
	wire \mchip.top.bobby.runway_manager.clock ;
	wire [3:0] \mchip.top.bobby.runway_manager.plane_id_lock ;
	wire [3:0] \mchip.top.bobby.runway_manager.plane_id_unlock ;
	wire \mchip.top.bobby.runway_manager.reset ;
	reg [9:0] \mchip.top.bobby.runway_manager.runway ;
	wire [1:0] \mchip.top.bobby.runway_manager.runway_active ;
	wire [1:0] \mchip.top.bobby.runway_manager.runway_override ;
	wire [1:0] \mchip.top.bobby.runway_override ;
	wire \mchip.top.bobby.send_reply ;
	wire \mchip.top.bobby.set_emergency ;
	wire \mchip.top.bobby.takeoff_fifo.clock ;
	reg [3:0] \mchip.top.bobby.takeoff_fifo.count ;
	wire [3:0] \mchip.top.bobby.takeoff_fifo.data_in ;
	reg [3:0] \mchip.top.bobby.takeoff_fifo.data_out ;
	reg [2:0] \mchip.top.bobby.takeoff_fifo.get_ptr ;
	reg [2:0] \mchip.top.bobby.takeoff_fifo.put_ptr ;
	reg [31:0] \mchip.top.bobby.takeoff_fifo.queue ;
	wire \mchip.top.bobby.takeoff_fifo.reset ;
	wire \mchip.top.bobby.uart_replies.clock ;
	reg [2:0] \mchip.top.bobby.uart_replies.count ;
	wire [7:0] \mchip.top.bobby.uart_replies.data_in ;
	reg [7:0] \mchip.top.bobby.uart_replies.data_out ;
	reg [1:0] \mchip.top.bobby.uart_replies.get_ptr ;
	reg [1:0] \mchip.top.bobby.uart_replies.put_ptr ;
	reg [31:0] \mchip.top.bobby.uart_replies.queue ;
	wire \mchip.top.bobby.uart_replies.re ;
	wire \mchip.top.bobby.uart_replies.reset ;
	wire [7:0] \mchip.top.bobby.uart_request ;
	wire \mchip.top.bobby.uart_requests.clock ;
	reg [2:0] \mchip.top.bobby.uart_requests.count ;
	wire [7:0] \mchip.top.bobby.uart_requests.data_in ;
	reg [7:0] \mchip.top.bobby.uart_requests.data_out ;
	reg [1:0] \mchip.top.bobby.uart_requests.get_ptr ;
	reg [1:0] \mchip.top.bobby.uart_requests.put_ptr ;
	reg [31:0] \mchip.top.bobby.uart_requests.queue ;
	wire \mchip.top.bobby.uart_requests.reset ;
	wire [7:0] \mchip.top.bobby.uart_rx_data ;
	wire [7:0] \mchip.top.bobby.uart_tx_data ;
	wire \mchip.top.bobby.uart_tx_send ;
	wire \mchip.top.clock ;
	wire \mchip.top.emergency ;
	wire \mchip.top.emergency_override ;
	reg \mchip.top.eo_sync ;
	reg \mchip.top.eo_temp ;
	wire \mchip.top.framing_error ;
	wire \mchip.top.receiver.clock ;
	wire \mchip.top.receiver.conductor.clock ;
	reg [9:0] \mchip.top.receiver.conductor.clockCount ;
	wire \mchip.top.receiver.conductor.reset ;
	wire \mchip.top.receiver.conductor.start_tx ;
	reg [7:0] \mchip.top.receiver.data ;
	reg [3:0] \mchip.top.receiver.data_counter ;
	wire \mchip.top.receiver.framing_error ;
	wire \mchip.top.receiver.fsm.clock ;
	wire \mchip.top.receiver.fsm.framing_error ;
	wire \mchip.top.receiver.fsm.receiving ;
	wire \mchip.top.receiver.fsm.reset ;
	wire \mchip.top.receiver.fsm.rx ;
	reg [3:0] \mchip.top.receiver.fsm.state ;
	wire \mchip.top.receiver.receiving ;
	wire \mchip.top.receiver.reset ;
	wire \mchip.top.receiver.rx ;
	wire \mchip.top.receiving ;
	wire \mchip.top.reset ;
	reg [1:0] \mchip.top.ro_sync ;
	reg [1:0] \mchip.top.ro_temp ;
	wire [1:0] \mchip.top.runway_active ;
	wire [1:0] \mchip.top.runway_override ;
	wire \mchip.top.rx ;
	wire \mchip.top.sending ;
	wire \mchip.top.transmitter.clock ;
	wire \mchip.top.transmitter.conductor.clock ;
	reg [9:0] \mchip.top.transmitter.conductor.clockCount ;
	wire \mchip.top.transmitter.conductor.reset ;
	wire \mchip.top.transmitter.conductor.start_rx ;
	wire [7:0] \mchip.top.transmitter.data ;
	reg \mchip.top.transmitter.data_bit ;
	reg [3:0] \mchip.top.transmitter.data_counter ;
	wire \mchip.top.transmitter.fsm.clock ;
	wire \mchip.top.transmitter.fsm.reset ;
	wire \mchip.top.transmitter.fsm.send ;
	wire \mchip.top.transmitter.fsm.sending ;
	reg [3:0] \mchip.top.transmitter.fsm.state ;
	wire \mchip.top.transmitter.reset ;
	reg [7:0] \mchip.top.transmitter.saved_data ;
	wire \mchip.top.transmitter.send ;
	wire \mchip.top.transmitter.sending ;
	reg \mchip.top.transmitter.tx ;
	wire \mchip.top.tx ;
	wire [7:0] \mchip.top.uart_rx_data ;
	wire [7:0] \mchip.top.uart_tx_data ;
	wire \mchip.top.uart_tx_send ;
	assign _1652_[0] = ~\mchip.top.transmitter.data_counter [0];
	assign _1650_[0] = ~\mchip.top.receiver.conductor.clockCount [0];
	assign _1643_[0] = ~\mchip.top.bobby.uart_requests.get_ptr [0];
	assign io_out[2] = \mchip.top.bobby.runway_manager.runway [0] | \mchip.top.ro_sync [0];
	assign io_out[3] = \mchip.top.bobby.runway_manager.runway [5] | \mchip.top.ro_sync [1];
	assign _1648_[0] = ~\mchip.top.receiver.data_counter [0];
	assign _1633_[0] = ~\mchip.top.bobby.takeoff_fifo.get_ptr [0];
	assign _1647_[0] = ~\mchip.top.bobby.uart_requests.count [0];
	assign _0038_ = ~\mchip.top.bobby.fsm.takeoff_first ;
	assign _1637_[0] = ~\mchip.top.bobby.takeoff_fifo.count [0];
	assign _1285_ = \mchip.top.bobby.fsm.state [7] | \mchip.top.bobby.fsm.state [6];
	assign _1286_ = \mchip.top.bobby.fsm.state [3] | \mchip.top.bobby.fsm.state [4];
	assign _1287_ = \mchip.top.bobby.fsm.state [2] | \mchip.top.bobby.fsm.state [0];
	assign _1288_ = _1287_ | _1286_;
	assign _1289_ = ~(_1288_ | _1285_);
	assign _1290_ = io_out[3] & io_out[2];
	assign _1291_ = _1289_ & ~_1290_;
	assign _1292_ = ~\mchip.top.bobby.uart_requests.data_out [7];
	assign _1293_ = ~\mchip.top.bobby.uart_requests.data_out [6];
	assign _1294_ = ~\mchip.top.bobby.uart_requests.data_out [5];
	assign _1295_ = (\mchip.top.bobby.uart_requests.data_out [4] ? \mchip.top.bobby.id_manager.taken_id [1] : \mchip.top.bobby.id_manager.taken_id [0]);
	assign _1296_ = (\mchip.top.bobby.uart_requests.data_out [4] ? \mchip.top.bobby.id_manager.taken_id [3] : \mchip.top.bobby.id_manager.taken_id [2]);
	assign _1297_ = (\mchip.top.bobby.uart_requests.data_out [5] ? _1296_ : _1295_);
	assign _1298_ = (\mchip.top.bobby.uart_requests.data_out [4] ? \mchip.top.bobby.id_manager.taken_id [5] : \mchip.top.bobby.id_manager.taken_id [4]);
	assign _1299_ = (\mchip.top.bobby.uart_requests.data_out [4] ? \mchip.top.bobby.id_manager.taken_id [7] : \mchip.top.bobby.id_manager.taken_id [6]);
	assign _1300_ = (\mchip.top.bobby.uart_requests.data_out [5] ? _1299_ : _1298_);
	assign _1301_ = (\mchip.top.bobby.uart_requests.data_out [6] ? _1300_ : _1297_);
	assign _1302_ = (\mchip.top.bobby.uart_requests.data_out [4] ? \mchip.top.bobby.id_manager.taken_id [9] : \mchip.top.bobby.id_manager.taken_id [8]);
	assign _1303_ = (\mchip.top.bobby.uart_requests.data_out [4] ? \mchip.top.bobby.id_manager.taken_id [11] : \mchip.top.bobby.id_manager.taken_id [10]);
	assign _1304_ = (\mchip.top.bobby.uart_requests.data_out [5] ? _1303_ : _1302_);
	assign _1305_ = (\mchip.top.bobby.uart_requests.data_out [4] ? \mchip.top.bobby.id_manager.taken_id [13] : \mchip.top.bobby.id_manager.taken_id [12]);
	assign _1306_ = (\mchip.top.bobby.uart_requests.data_out [4] ? \mchip.top.bobby.id_manager.taken_id [15] : \mchip.top.bobby.id_manager.taken_id [14]);
	assign _1307_ = (\mchip.top.bobby.uart_requests.data_out [5] ? _1306_ : _1305_);
	assign _1308_ = (\mchip.top.bobby.uart_requests.data_out [6] ? _1307_ : _1304_);
	assign _1309_ = (\mchip.top.bobby.uart_requests.data_out [7] ? _1308_ : _1301_);
	assign _1310_ = ~\mchip.top.bobby.uart_requests.data_out [3];
	assign _1311_ = \mchip.top.bobby.uart_requests.data_out [2] | ~\mchip.top.bobby.uart_requests.data_out [1];
	assign _1312_ = _1310_ & ~_1311_;
	assign _1313_ = _1312_ & _1309_;
	assign _1314_ = \mchip.top.bobby.uart_requests.data_out [1] | \mchip.top.bobby.uart_requests.data_out [2];
	assign _1315_ = _1310_ & ~_1314_;
	assign _1316_ = _1313_ & ~_1315_;
	assign _1317_ = \mchip.top.bobby.fsm.state [5] | \mchip.top.bobby.fsm.state [6];
	assign _1318_ = _1317_ | \mchip.top.bobby.fsm.state [7];
	assign _1319_ = \mchip.top.bobby.fsm.state [3] | \mchip.top.bobby.fsm.state [2];
	assign _1320_ = \mchip.top.bobby.fsm.state [1] | \mchip.top.bobby.fsm.state [0];
	assign _1321_ = _1320_ | _1319_;
	assign _1322_ = ~(_1321_ | _1318_);
	assign _1323_ = _1322_ & _1316_;
	assign _0040_ = _1291_ & ~_1323_;
	assign _1324_ = \mchip.top.bobby.fsm.state [5] & ~_1290_;
	assign _1325_ = ~\mchip.top.bobby.fsm.state [5];
	assign _1326_ = ~(_1289_ & _1325_);
	assign _1327_ = ~(_1326_ | _1290_);
	assign _1328_ = _1327_ ^ _1324_;
	assign _0039_ = ~_1328_;
	assign _1632_[0] = ~\mchip.top.bobby.landing_fifo.count [0];
	assign _1642_[0] = ~\mchip.top.bobby.uart_replies.count [0];
	assign _1329_ = ~(\mchip.top.bobby.emergency  | \mchip.top.eo_sync );
	assign \mchip.top.bobby.emergency_out  = ~_1329_;
	assign _1330_ = \mchip.top.bobby.uart_requests.count [1] | \mchip.top.bobby.uart_requests.count [0];
	assign _1331_ = _1330_ | \mchip.top.bobby.uart_requests.count [2];
	assign _1332_ = _1331_ | _1329_;
	assign _1333_ = ~io_in[13];
	assign _1334_ = ~(\mchip.top.bobby.landing_fifo.count [1] | \mchip.top.bobby.landing_fifo.count [0]);
	assign _1335_ = \mchip.top.bobby.landing_fifo.count [3] | \mchip.top.bobby.landing_fifo.count [2];
	assign _1336_ = _1334_ & ~_1335_;
	assign _1337_ = ~(_1336_ & _1333_);
	assign _1338_ = _1337_ | _1332_;
	assign _1339_ = \mchip.top.bobby.fsm.state [0] & ~_1338_;
	assign _1340_ = ~(\mchip.top.bobby.takeoff_fifo.count [1] | \mchip.top.bobby.takeoff_fifo.count [0]);
	assign _1341_ = \mchip.top.bobby.takeoff_fifo.count [3] | \mchip.top.bobby.takeoff_fifo.count [2];
	assign _1342_ = _1340_ & ~_1341_;
	assign _1343_ = ~(_1342_ | _1336_);
	assign _1344_ = _1343_ | _1290_;
	assign _1345_ = _1344_ | _1331_;
	assign _1346_ = ~(_1336_ & _1329_);
	assign _1347_ = ~(_1342_ & _1333_);
	assign _1348_ = _1347_ | _1346_;
	assign _1349_ = _1348_ | _1345_;
	assign _1350_ = \mchip.top.bobby.fsm.state [0] & ~_1349_;
	assign _1351_ = _1348_ | _1344_;
	assign _1352_ = \mchip.top.bobby.fsm.state [6] & ~_1351_;
	assign _1353_ = _1352_ | _1350_;
	assign _1354_ = ~(_1329_ & _1333_);
	assign _1355_ = _1354_ | ~_1290_;
	assign _1356_ = \mchip.top.bobby.fsm.state [6] & ~_1355_;
	assign _1357_ = _1356_ | \mchip.top.bobby.fsm.state [7];
	assign _1358_ = _1357_ | _1353_;
	assign _1359_ = _1331_ | ~_1290_;
	assign _1360_ = _1359_ | _1354_;
	assign _1361_ = \mchip.top.bobby.fsm.state [0] & ~_1360_;
	assign _1362_ = \mchip.top.bobby.uart_requests.data_out [2] & ~\mchip.top.bobby.uart_requests.data_out [1];
	assign _1363_ = _1362_ & ~\mchip.top.bobby.uart_requests.data_out [3];
	assign _1364_ = ~(_1363_ & \mchip.top.bobby.uart_requests.data_out [0]);
	assign _1365_ = ~(\mchip.top.bobby.uart_requests.data_out [2] | \mchip.top.bobby.uart_requests.data_out [3]);
	assign _1366_ = _1365_ | _1337_;
	assign _1367_ = _1366_ | _1364_;
	assign _1368_ = \mchip.top.bobby.fsm.state [4] & ~_1367_;
	assign _1369_ = _1368_ | _1361_;
	assign _1370_ = _1337_ | _1329_;
	assign _1371_ = \mchip.top.bobby.fsm.state [6] & ~_1370_;
	assign _1372_ = _1371_ | io_in[13];
	assign _1373_ = _1372_ | _1369_;
	assign _1374_ = _1373_ | _1358_;
	assign _0002_ = _1374_ | _1339_;
	assign _1375_ = \mchip.top.bobby.uart_replies.count [1] | \mchip.top.bobby.uart_replies.count [0];
	assign _1376_ = \mchip.top.bobby.uart_replies.count [2] & ~_1375_;
	assign _1377_ = _1376_ | io_in[13];
	assign _1378_ = \mchip.top.bobby.fsm.state [2] & ~_1377_;
	assign _1379_ = _1315_ | io_in[13];
	assign _1380_ = _1379_ | ~_1312_;
	assign _1381_ = \mchip.top.bobby.fsm.state [4] & ~_1380_;
	assign _1382_ = _1381_ | _1378_;
	assign _1383_ = _1315_ & ~io_in[13];
	assign _1384_ = _1309_ | ~_1383_;
	assign _1385_ = \mchip.top.bobby.fsm.state [4] & ~_1384_;
	assign _1386_ = _1312_ | ~_1363_;
	assign _1387_ = _1386_ | _1379_;
	assign _1388_ = _1387_ | \mchip.top.bobby.uart_requests.data_out [0];
	assign _1389_ = \mchip.top.bobby.fsm.state [4] & ~_1388_;
	assign _1390_ = _1389_ | _1385_;
	assign _0007_ = _1390_ | _1382_;
	assign _1391_ = ~io_in[0];
	assign _1392_ = \mchip.top.receiver.conductor.clockCount [8] | \mchip.top.receiver.conductor.clockCount [9];
	assign _1393_ = ~(\mchip.top.receiver.conductor.clockCount [6] & \mchip.top.receiver.conductor.clockCount [7]);
	assign _1394_ = \mchip.top.receiver.conductor.clockCount [5] | ~\mchip.top.receiver.conductor.clockCount [4];
	assign _1395_ = _1394_ | _1393_;
	assign _1396_ = \mchip.top.receiver.conductor.clockCount [2] | ~\mchip.top.receiver.conductor.clockCount [3];
	assign _1397_ = \mchip.top.receiver.conductor.clockCount [1] | ~\mchip.top.receiver.conductor.clockCount [0];
	assign _1398_ = _1397_ | _1396_;
	assign _1399_ = _1398_ | _1395_;
	assign _1400_ = _1399_ | _1392_;
	assign _1401_ = _1400_ | _1391_;
	assign _1402_ = _1333_ & ~_1401_;
	assign _1403_ = ~(\mchip.top.receiver.fsm.state [2] | \mchip.top.receiver.fsm.state [3]);
	assign _1404_ = _1402_ & ~_1403_;
	assign _1405_ = ~(\mchip.top.receiver.data_counter [1] | \mchip.top.receiver.data_counter [0]);
	assign _1406_ = \mchip.top.receiver.data_counter [2] | ~\mchip.top.receiver.data_counter [3];
	assign _1407_ = _1405_ & ~_1406_;
	assign _1408_ = _1400_ | ~_1407_;
	assign _1409_ = io_in[13] | ~io_in[0];
	assign _1410_ = _1409_ | _1408_;
	assign _1411_ = \mchip.top.receiver.fsm.state [1] & ~_1410_;
	assign _1412_ = _1391_ & ~_1400_;
	assign _1413_ = ~(_1401_ & _1333_);
	assign _1414_ = _1413_ | _1412_;
	assign _1415_ = \mchip.top.receiver.fsm.state [3] & ~_1414_;
	assign _1416_ = _1415_ | _1411_;
	assign _1417_ = \mchip.top.receiver.fsm.state [0] & ~_1409_;
	assign _1418_ = _1417_ | io_in[13];
	assign _1419_ = _1418_ | _1416_;
	assign _0008_ = _1419_ | _1404_;
	assign _1420_ = \mchip.top.transmitter.fsm.state [1] | \mchip.top.transmitter.fsm.state [2];
	assign \mchip.top.sending  = _1420_ | \mchip.top.transmitter.fsm.state [3];
	assign _1421_ = \mchip.top.bobby.reply_fsm.state  & ~\mchip.top.sending ;
	assign _1422_ = \mchip.top.transmitter.conductor.clockCount [0] & ~\mchip.top.transmitter.conductor.clockCount [1];
	assign _1423_ = \mchip.top.transmitter.conductor.clockCount [2] | ~\mchip.top.transmitter.conductor.clockCount [3];
	assign _1424_ = _1422_ & ~_1423_;
	assign _1425_ = ~(\mchip.top.transmitter.conductor.clockCount [6] & \mchip.top.transmitter.conductor.clockCount [7]);
	assign _1426_ = \mchip.top.transmitter.conductor.clockCount [5] | ~\mchip.top.transmitter.conductor.clockCount [4];
	assign _1427_ = _1426_ | _1425_;
	assign _1428_ = _1424_ & ~_1427_;
	assign _1429_ = \mchip.top.transmitter.conductor.clockCount [8] | \mchip.top.transmitter.conductor.clockCount [9];
	assign _1430_ = _1428_ & ~_1429_;
	assign _1431_ = _1430_ | io_in[13];
	assign _0036_ = _1431_ | _1421_;
	assign _0198_ = ~(_1400_ & _1333_);
	assign _1432_ = \mchip.top.receiver.fsm.state [2] | \mchip.top.receiver.fsm.state [1];
	assign _1433_ = _1432_ | \mchip.top.receiver.fsm.state [3];
	assign _1434_ = _1391_ & ~_1433_;
	assign _0037_ = _1434_ | _0198_;
	assign _1435_ = ~(_1407_ | _1400_);
	assign _1436_ = ~(_1435_ & _1333_);
	assign _1437_ = \mchip.top.receiver.fsm.state [1] & ~_1436_;
	assign _1438_ = \mchip.top.receiver.fsm.state [1] & ~_0198_;
	assign _1439_ = _1413_ | ~_1412_;
	assign _1440_ = \mchip.top.receiver.fsm.state [2] & ~_1439_;
	assign _1441_ = _1440_ | _1438_;
	assign _0009_ = _1441_ | _1437_;
	assign _1442_ = \mchip.top.receiver.fsm.state [2] & ~_1414_;
	assign _1443_ = io_in[0] | io_in[13];
	assign _1444_ = \mchip.top.receiver.fsm.state [0] & ~_1443_;
	assign _0010_ = _1444_ | _1442_;
	assign _1445_ = \mchip.top.receiver.fsm.state [3] & ~_1439_;
	assign _1446_ = _1443_ | _1408_;
	assign _1447_ = \mchip.top.receiver.fsm.state [1] & ~_1446_;
	assign _0011_ = _1447_ | _1445_;
	assign _1448_ = ~_1430_;
	assign _1449_ = ~\mchip.top.transmitter.fsm.state [1];
	assign _1450_ = \mchip.top.transmitter.data_counter [2] | ~\mchip.top.transmitter.data_counter [3];
	assign _1451_ = \mchip.top.transmitter.data_counter [1] | \mchip.top.transmitter.data_counter [0];
	assign _1452_ = _1451_ | _1450_;
	assign _1453_ = _1430_ & ~_1452_;
	assign _1454_ = _1453_ | _1449_;
	assign _1455_ = \mchip.top.transmitter.fsm.state [0] | \mchip.top.transmitter.fsm.state [3];
	assign _1456_ = _1449_ & ~_1455_;
	assign _1457_ = (_1456_ ? _1448_ : _1454_);
	assign _0199_ = _1430_ & ~_1457_;
	assign _0016_ = _0199_ | _1421_;
	assign _1458_ = \mchip.top.bobby.reply_fsm.state  | io_in[13];
	assign _1459_ = \mchip.top.transmitter.fsm.state [0] & ~_1458_;
	assign _1460_ = ~(_1430_ & _1333_);
	assign _1461_ = \mchip.top.transmitter.fsm.state [3] & ~_1460_;
	assign _1462_ = _1461_ | io_in[13];
	assign _0012_ = _1462_ | _1459_;
	assign _1463_ = \mchip.top.transmitter.fsm.state [2] & ~_1460_;
	assign _1464_ = _1453_ | io_in[13];
	assign _1465_ = \mchip.top.transmitter.fsm.state [1] & ~_1464_;
	assign _0013_ = _1465_ | _1463_;
	assign _1466_ = io_in[13] | ~\mchip.top.bobby.reply_fsm.state ;
	assign _1467_ = \mchip.top.transmitter.fsm.state [0] & ~_1466_;
	assign _1468_ = \mchip.top.transmitter.fsm.state [2] & ~_1431_;
	assign _0014_ = _1468_ | _1467_;
	assign _1469_ = \mchip.top.transmitter.fsm.state [3] & ~_1431_;
	assign _1470_ = ~(_1453_ & _1333_);
	assign _1471_ = \mchip.top.transmitter.fsm.state [1] & ~_1470_;
	assign _0015_ = _1471_ | _1469_;
	assign _1472_ = ~(\mchip.top.receiver.fsm.state [2] | \mchip.top.receiver.fsm.state [0]);
	assign \mchip.top.receiver.fsm.receiving  = _1472_ & ~\mchip.top.receiver.fsm.state [3];
	assign _1473_ = \mchip.top.bobby.fsm.state [1] | \mchip.top.bobby.fsm.state [2];
	assign _1474_ = _1473_ | _1286_;
	assign _1475_ = _1474_ | _1318_;
	assign _1476_ = _1331_ & ~_1475_;
	assign _1477_ = _1408_ | _1391_;
	assign _1478_ = _1477_ | _1435_;
	assign _1479_ = \mchip.top.receiver.fsm.receiving  & ~_1478_;
	assign _1480_ = \mchip.top.bobby.uart_requests.count [2] & ~_1330_;
	assign _1481_ = _1479_ & ~_1480_;
	assign _0019_ = (_1476_ ? _1479_ : _1481_);
	assign _1482_ = ~_1479_;
	assign _0020_ = (_1476_ ? _1482_ : _1481_);
	assign _1483_ = _1479_ | ~_1476_;
	assign _1484_ = ~(_1481_ | _1476_);
	assign _1485_ = _1484_ | io_in[13];
	assign _0021_ = _1483_ & ~_1485_;
	assign _1486_ = ~(_1430_ & \mchip.top.transmitter.fsm.state [3]);
	assign _1487_ = (\mchip.top.sending  ? _1486_ : \mchip.top.bobby.reply_fsm.state );
	assign _1488_ = ~(_1375_ | \mchip.top.bobby.uart_replies.count [2]);
	assign _1489_ = _1488_ | _1487_;
	assign \mchip.top.bobby.reply_fsm.next_state  = ~(_1489_ | \mchip.top.bobby.reply_fsm.state );
	assign _1490_ = \mchip.top.bobby.reply_fsm.next_state  & ~_1488_;
	assign _1491_ = ~_1376_;
	assign _1492_ = _1320_ | _1286_;
	assign _1493_ = _1492_ | _1317_;
	assign _1494_ = _1493_ | \mchip.top.bobby.fsm.state [7];
	assign _1495_ = (_1494_ ? \mchip.top.bobby.fsm.state [7] : _1491_);
	assign _1496_ = _1495_ & ~_1376_;
	assign _0022_ = (_1490_ ? _1495_ : _1496_);
	assign _1497_ = ~_1495_;
	assign _0023_ = (_1490_ ? _1497_ : _1496_);
	assign _1498_ = _1495_ | ~_1490_;
	assign _1499_ = ~(_1496_ | _1490_);
	assign _1500_ = _1499_ | io_in[13];
	assign _0024_ = _1498_ & ~_1500_;
	assign _1501_ = (_1343_ ? _0038_ : _1342_);
	assign _1502_ = _1501_ | _1290_;
	assign _1503_ = _1502_ | \mchip.top.bobby.emergency_out ;
	assign _1504_ = ~\mchip.top.bobby.fsm.state [6];
	assign _1505_ = \mchip.top.bobby.fsm.state [5] | \mchip.top.bobby.fsm.state [7];
	assign _1506_ = _1505_ | _1474_;
	assign _1507_ = _1506_ | \mchip.top.bobby.fsm.state [6];
	assign _1508_ = (_1507_ ? _1504_ : _1331_);
	assign _1509_ = _1508_ | _1503_;
	assign _1510_ = ~(_1509_ | _1342_);
	assign _1511_ = ~\mchip.top.bobby.uart_requests.data_out [0];
	assign _1512_ = \mchip.top.bobby.takeoff_fifo.count [2] | ~\mchip.top.bobby.takeoff_fifo.count [3];
	assign _1513_ = _1340_ & ~_1512_;
	assign _1514_ = _1511_ & ~_1513_;
	assign _1515_ = _1514_ & _1309_;
	assign _1516_ = ~(_1515_ & _1315_);
	assign _1517_ = _1322_ & ~_1516_;
	assign _1518_ = _1517_ & ~_1513_;
	assign _0025_ = (_1510_ ? _1517_ : _1518_);
	assign _1519_ = ~_1517_;
	assign _0026_ = (_1510_ ? _1519_ : _1518_);
	assign _1520_ = ~(_1519_ & _1510_);
	assign _1521_ = ~(_1518_ | _1510_);
	assign _1522_ = _1521_ | io_in[13];
	assign _0027_ = _1520_ & ~_1522_;
	assign _1523_ = io_out[2] & ~io_out[3];
	assign _1524_ = ~(\mchip.top.bobby.fsm.state [5] | \mchip.top.bobby.fsm.state [1]);
	assign _1525_ = _1523_ & ~_1524_;
	assign _1526_ = \mchip.top.bobby.fsm.state [6] | \mchip.top.bobby.fsm.state [3];
	assign _1527_ = _1526_ | _1287_;
	assign _1528_ = ~(_1527_ | \mchip.top.bobby.fsm.state [7]);
	assign _1529_ = ~(_1528_ & _1524_);
	assign _1530_ = ~(_1309_ & \mchip.top.bobby.uart_requests.data_out [0]);
	assign _1531_ = _1530_ | ~_1312_;
	assign _1532_ = ~(_1531_ | _1315_);
	assign _1533_ = (_1529_ ? _1525_ : _1532_);
	assign _0028_ = _0040_ & ~_1533_;
	assign _0029_ = _1533_ & _0040_;
	assign _1534_ = _1291_ | ~_1323_;
	assign _1535_ = \mchip.top.bobby.runway_manager.runway [6] ^ \mchip.top.bobby.uart_requests.data_out [4];
	assign _1536_ = \mchip.top.bobby.runway_manager.runway [7] ^ \mchip.top.bobby.uart_requests.data_out [5];
	assign _1537_ = ~(_1536_ | _1535_);
	assign _1538_ = \mchip.top.bobby.runway_manager.runway [9] ^ \mchip.top.bobby.uart_requests.data_out [7];
	assign _1539_ = \mchip.top.bobby.runway_manager.runway [8] ^ \mchip.top.bobby.uart_requests.data_out [6];
	assign _1540_ = _1539_ | _1538_;
	assign _1541_ = _1537_ & ~_1540_;
	assign _1542_ = _1541_ | ~_1533_;
	assign _1543_ = (_1534_ ? _0040_ : _1542_);
	assign _1544_ = ~(_1534_ | _1533_);
	assign _1545_ = _1544_ | _0028_;
	assign _0030_ = _1543_ & ~_1545_;
	assign _1546_ = \mchip.top.bobby.runway_manager.runway [1] ^ \mchip.top.bobby.uart_requests.data_out [4];
	assign _1547_ = \mchip.top.bobby.runway_manager.runway [2] ^ \mchip.top.bobby.uart_requests.data_out [5];
	assign _1548_ = ~(_1547_ | _1546_);
	assign _1549_ = \mchip.top.bobby.runway_manager.runway [4] ^ \mchip.top.bobby.uart_requests.data_out [7];
	assign _1550_ = \mchip.top.bobby.runway_manager.runway [3] ^ \mchip.top.bobby.uart_requests.data_out [6];
	assign _1551_ = _1550_ | _1549_;
	assign _1552_ = _1548_ & ~_1551_;
	assign _1553_ = _1552_ | _1533_;
	assign _1554_ = (_1534_ ? _0040_ : _1553_);
	assign _1555_ = _1533_ & ~_1534_;
	assign _1556_ = _1555_ | _0029_;
	assign _0031_ = _1554_ & ~_1556_;
	assign _1557_ = _1336_ | ~_1342_;
	assign _1558_ = (_1343_ ? \mchip.top.bobby.fsm.takeoff_first  : _1557_);
	assign _1559_ = _1558_ | _1290_;
	assign _1560_ = (_1329_ ? _1559_ : _1336_);
	assign _1561_ = _1560_ | _1504_;
	assign _1562_ = ~_1363_;
	assign _1563_ = _1336_ | _1511_;
	assign _1564_ = _1563_ | _1562_;
	assign _1565_ = _1564_ | _1312_;
	assign _1566_ = _1565_ | _1315_;
	assign _1567_ = \mchip.top.bobby.fsm.state [4] & ~_1566_;
	assign _1568_ = _1561_ & ~_1567_;
	assign _1569_ = \mchip.top.bobby.fsm.state [5] | \mchip.top.bobby.fsm.state [3];
	assign _1570_ = _1569_ | _1473_;
	assign _1571_ = _1570_ | \mchip.top.bobby.fsm.state [7];
	assign _1572_ = _1571_ | \mchip.top.bobby.fsm.state [6];
	assign _1573_ = _1572_ | \mchip.top.bobby.fsm.state [4];
	assign _1574_ = _1560_ | _1331_;
	assign _1575_ = (_1573_ ? _1568_ : _1574_);
	assign _1576_ = ~(_1575_ | _1336_);
	assign _1577_ = \mchip.top.bobby.landing_fifo.count [2] | ~\mchip.top.bobby.landing_fifo.count [3];
	assign _1578_ = _1334_ & ~_1577_;
	assign _1579_ = _1578_ | \mchip.top.bobby.emergency_out ;
	assign _1580_ = \mchip.top.bobby.uart_requests.data_out [0] & ~_1579_;
	assign _1581_ = ~(_1580_ & _1309_);
	assign _1582_ = _1581_ | ~_1315_;
	assign _1583_ = _1322_ & ~_1582_;
	assign _1584_ = _1583_ & ~_1578_;
	assign _0032_ = (_1576_ ? _1583_ : _1584_);
	assign _1585_ = ~_1583_;
	assign _0033_ = (_1576_ ? _1585_ : _1584_);
	assign _1586_ = ~(_1585_ & _1576_);
	assign _1587_ = ~(_1584_ | _1576_);
	assign _1588_ = _1587_ | io_in[13];
	assign _0034_ = _1586_ & ~_1588_;
	assign _1589_ = ~(\mchip.top.bobby.id_manager.taken_id [15] & \mchip.top.bobby.id_manager.taken_id [14]);
	assign _1590_ = ~(\mchip.top.bobby.id_manager.taken_id [13] & \mchip.top.bobby.id_manager.taken_id [12]);
	assign _1591_ = _1590_ | _1589_;
	assign _1592_ = ~(\mchip.top.bobby.id_manager.taken_id [11] & \mchip.top.bobby.id_manager.taken_id [10]);
	assign _1593_ = ~(\mchip.top.bobby.id_manager.taken_id [9] & \mchip.top.bobby.id_manager.taken_id [8]);
	assign _1594_ = _1593_ | _1592_;
	assign _1595_ = _1594_ | _1591_;
	assign _1596_ = ~(\mchip.top.bobby.id_manager.taken_id [7] & \mchip.top.bobby.id_manager.taken_id [6]);
	assign _1597_ = ~(\mchip.top.bobby.id_manager.taken_id [5] & \mchip.top.bobby.id_manager.taken_id [4]);
	assign _1598_ = _1597_ | _1596_;
	assign _1599_ = ~(\mchip.top.bobby.id_manager.taken_id [3] & \mchip.top.bobby.id_manager.taken_id [2]);
	assign _1600_ = ~(\mchip.top.bobby.id_manager.taken_id [1] & \mchip.top.bobby.id_manager.taken_id [0]);
	assign _1601_ = _1600_ | _1599_;
	assign _1602_ = _1601_ | _1598_;
	assign _1603_ = _1602_ | _1595_;
	assign _1604_ = \mchip.top.bobby.uart_requests.data_out [1] & \mchip.top.bobby.uart_requests.data_out [2];
	assign _1605_ = ~(_1604_ & \mchip.top.bobby.uart_requests.data_out [3]);
	assign _1606_ = _1605_ | ~_1603_;
	assign _1607_ = _1606_ | ~_1562_;
	assign _1608_ = _1607_ | _1312_;
	assign _1609_ = _1608_ | _1315_;
	assign _1610_ = _1609_ | ~_1322_;
	assign _1611_ = _1603_ & ~_1610_;
	assign _1612_ = _1363_ & ~\mchip.top.bobby.uart_requests.data_out [0];
	assign _1613_ = ~(_1552_ & \mchip.top.bobby.runway_manager.runway [0]);
	assign _1614_ = ~(_1541_ & \mchip.top.bobby.runway_manager.runway [5]);
	assign _1615_ = (\mchip.top.bobby.uart_requests.data_out [0] ? _1614_ : _1613_);
	assign _1616_ = _1309_ & ~_1615_;
	assign _1617_ = (_1312_ ? _1616_ : _1612_);
	assign _1618_ = _1580_ | _1514_;
	assign _1619_ = _1309_ & ~_1618_;
	assign _1620_ = (_1315_ ? _1619_ : _1617_);
	assign _1621_ = \mchip.top.bobby.fsm.state [5] | \mchip.top.bobby.fsm.state [2];
	assign _1622_ = _1621_ | _1320_;
	assign _1623_ = _1622_ | _1285_;
	assign _1624_ = _1623_ | \mchip.top.bobby.fsm.state [3];
	assign _1625_ = (_1624_ ? \mchip.top.bobby.fsm.state [3] : _1620_);
	assign _0017_ = _1625_ | _1611_;
	assign _1626_ = \mchip.top.bobby.fsm.state [4] | \mchip.top.bobby.fsm.state [2];
	assign _1627_ = _1626_ | _1320_;
	assign _0211_ = _1627_ | _1318_;
	assign _0212_ = ~(_0211_ & _1610_);
	assign _0213_ = _0212_ | _1328_;
	assign _0214_ = _1605_ | _1603_;
	assign _0215_ = _0214_ | ~_1562_;
	assign _0216_ = _0215_ | _1312_;
	assign _0217_ = _0216_ | _1315_;
	assign _0218_ = _0217_ | ~_1322_;
	assign _0219_ = ~(_1619_ & _1315_);
	assign _0220_ = _1322_ & ~_0219_;
	assign _0221_ = _0218_ & ~_0220_;
	assign _0222_ = (\mchip.top.bobby.uart_requests.data_out [3] ? _1604_ : _1362_);
	assign _0223_ = _0222_ | _1312_;
	assign _0224_ = _0223_ | _1315_;
	assign _0225_ = _1322_ & ~_0224_;
	assign _0226_ = ~(_1618_ & _1309_);
	assign _0227_ = _0226_ | ~_1315_;
	assign _0228_ = _1322_ & ~_0227_;
	assign _0229_ = ~(_0228_ | _0225_);
	assign _0230_ = ~(_0229_ & _0221_);
	assign _0035_ = _0230_ | _0213_;
	assign _0231_ = _1364_ | _1312_;
	assign _0232_ = _0231_ | _1315_;
	assign \mchip.top.bobby.fsm.set_emergency  = _1322_ & ~_0232_;
	assign _0233_ = \mchip.top.bobby.emergency_id [3] ^ \mchip.top.bobby.uart_requests.data_out [7];
	assign _0234_ = \mchip.top.bobby.emergency_id [2] ^ \mchip.top.bobby.uart_requests.data_out [6];
	assign _0235_ = _0234_ | _0233_;
	assign _0236_ = \mchip.top.bobby.emergency_id [1] ^ \mchip.top.bobby.uart_requests.data_out [5];
	assign _0237_ = \mchip.top.bobby.emergency_id [0] ^ \mchip.top.bobby.uart_requests.data_out [4];
	assign _0238_ = _0237_ | _0236_;
	assign _0239_ = _0238_ | _0235_;
	assign _0240_ = _0239_ | \mchip.top.bobby.uart_requests.data_out [0];
	assign _0241_ = _0240_ | _1562_;
	assign _0242_ = _0241_ | _1312_;
	assign _0243_ = _0242_ | _1315_;
	assign _0244_ = _1322_ & ~_0243_;
	assign _0018_ = _0244_ | \mchip.top.bobby.fsm.set_emergency ;
	assign _1654_[0] = ~\mchip.top.transmitter.conductor.clockCount [0];
	assign _0245_ = _1336_ | \mchip.top.bobby.emergency_out ;
	assign _0246_ = _0245_ | _1347_;
	assign _0247_ = _0246_ | _1345_;
	assign _0248_ = \mchip.top.bobby.fsm.state [0] & ~_0247_;
	assign _0249_ = _0246_ | _1344_;
	assign _0250_ = \mchip.top.bobby.fsm.state [6] & ~_0249_;
	assign _0251_ = _0250_ | _0248_;
	assign _0252_ = _1331_ | ~_1343_;
	assign _0253_ = _1290_ | \mchip.top.bobby.fsm.takeoff_first ;
	assign _0254_ = _0253_ | _1354_;
	assign _0255_ = _0254_ | _0252_;
	assign _0256_ = \mchip.top.bobby.fsm.state [0] & ~_0255_;
	assign _0257_ = ~_1343_;
	assign _0258_ = _0254_ | _0257_;
	assign _0259_ = \mchip.top.bobby.fsm.state [6] & ~_0258_;
	assign _0260_ = _0259_ | _0256_;
	assign _0006_ = _0260_ | _0251_;
	assign _0261_ = _1336_ | io_in[13];
	assign _0262_ = _0261_ | _1332_;
	assign _0263_ = \mchip.top.bobby.fsm.state [0] & ~_0262_;
	assign _0264_ = _0261_ | _1329_;
	assign _0265_ = \mchip.top.bobby.fsm.state [6] & ~_0264_;
	assign _0266_ = _0261_ | _1365_;
	assign _0267_ = _0266_ | _1364_;
	assign _0268_ = \mchip.top.bobby.fsm.state [4] & ~_0267_;
	assign _0269_ = _0268_ | _0265_;
	assign _0005_ = _0269_ | _0263_;
	assign _0270_ = ~(_1376_ & _1333_);
	assign _0271_ = \mchip.top.bobby.fsm.state [2] & ~_0270_;
	assign _0272_ = _1363_ | _1312_;
	assign _0273_ = _0272_ | _1379_;
	assign _0274_ = \mchip.top.bobby.fsm.state [4] & ~_0273_;
	assign _0275_ = ~(_1383_ & _1309_);
	assign _0276_ = \mchip.top.bobby.fsm.state [4] & ~_0275_;
	assign _0277_ = _0276_ | _0274_;
	assign _0004_ = _0277_ | _0271_;
	assign _0278_ = _1290_ | _0038_;
	assign _0279_ = _0278_ | _1354_;
	assign _0280_ = _0279_ | _0257_;
	assign _0281_ = \mchip.top.bobby.fsm.state [6] & ~_0280_;
	assign _0282_ = _0279_ | _0252_;
	assign _0283_ = \mchip.top.bobby.fsm.state [0] & ~_0282_;
	assign _0284_ = _0283_ | _0281_;
	assign _0285_ = \mchip.top.bobby.emergency_out  | _1290_;
	assign _0286_ = _1342_ | io_in[13];
	assign _0287_ = _0286_ | _0285_;
	assign _0288_ = _0287_ | _1343_;
	assign _0289_ = \mchip.top.bobby.fsm.state [6] & ~_0288_;
	assign _0290_ = _1343_ | _1331_;
	assign _0291_ = _0290_ | _0287_;
	assign _0292_ = \mchip.top.bobby.fsm.state [0] & ~_0291_;
	assign _0293_ = _0292_ | _0289_;
	assign _0003_ = _0293_ | _0284_;
	assign _0294_ = \mchip.top.receiver.fsm.state [1] & ~_1478_;
	assign _0295_ = \mchip.top.receiver.fsm.state [3] & ~_1401_;
	assign _0296_ = _0295_ | _0294_;
	assign _0297_ = ~(\mchip.top.receiver.fsm.state [1] | \mchip.top.receiver.fsm.state [3]);
	assign _0298_ = _0296_ & ~_0297_;
	assign _0197_ = _0298_ | io_in[13];
	assign _0299_ = ~(\mchip.top.receiver.fsm.receiving  & _1435_);
	assign _0196_ = ~(_0299_ | _1400_);
	assign _0201_ = _1421_ | io_in[13];
	assign _0300_ = \mchip.top.transmitter.fsm.state [0] | \mchip.top.transmitter.fsm.state [2];
	assign _0301_ = _0300_ | \mchip.top.transmitter.fsm.state [3];
	assign _0302_ = _1453_ & ~_0301_;
	assign _0200_ = _0302_ | io_in[13];
	assign _0303_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [4] : \mchip.top.bobby.takeoff_fifo.queue [0]);
	assign _0304_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [12] : \mchip.top.bobby.takeoff_fifo.queue [8]);
	assign _0305_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [1] ? _0304_ : _0303_);
	assign _0306_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [20] : \mchip.top.bobby.takeoff_fifo.queue [16]);
	assign _0307_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [28] : \mchip.top.bobby.takeoff_fifo.queue [24]);
	assign _0308_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [1] ? _0307_ : _0306_);
	assign _1657_[0] = (\mchip.top.bobby.takeoff_fifo.get_ptr [2] ? _0308_ : _0305_);
	assign _0309_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [5] : \mchip.top.bobby.takeoff_fifo.queue [1]);
	assign _0310_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [13] : \mchip.top.bobby.takeoff_fifo.queue [9]);
	assign _0311_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [1] ? _0310_ : _0309_);
	assign _0312_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [21] : \mchip.top.bobby.takeoff_fifo.queue [17]);
	assign _0313_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [29] : \mchip.top.bobby.takeoff_fifo.queue [25]);
	assign _0314_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [1] ? _0313_ : _0312_);
	assign _1657_[1] = (\mchip.top.bobby.takeoff_fifo.get_ptr [2] ? _0314_ : _0311_);
	assign _0315_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [6] : \mchip.top.bobby.takeoff_fifo.queue [2]);
	assign _0316_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [14] : \mchip.top.bobby.takeoff_fifo.queue [10]);
	assign _0317_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [1] ? _0316_ : _0315_);
	assign _0318_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [22] : \mchip.top.bobby.takeoff_fifo.queue [18]);
	assign _0319_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [30] : \mchip.top.bobby.takeoff_fifo.queue [26]);
	assign _0320_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [1] ? _0319_ : _0318_);
	assign _1657_[2] = (\mchip.top.bobby.takeoff_fifo.get_ptr [2] ? _0320_ : _0317_);
	assign _0321_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [7] : \mchip.top.bobby.takeoff_fifo.queue [3]);
	assign _0322_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [15] : \mchip.top.bobby.takeoff_fifo.queue [11]);
	assign _0323_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [1] ? _0322_ : _0321_);
	assign _0324_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [23] : \mchip.top.bobby.takeoff_fifo.queue [19]);
	assign _0325_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [0] ? \mchip.top.bobby.takeoff_fifo.queue [31] : \mchip.top.bobby.takeoff_fifo.queue [27]);
	assign _0326_ = (\mchip.top.bobby.takeoff_fifo.get_ptr [1] ? _0325_ : _0324_);
	assign _1657_[3] = (\mchip.top.bobby.takeoff_fifo.get_ptr [2] ? _0326_ : _0323_);
	assign _0327_ = _1408_ | io_in[0];
	assign _0328_ = _0327_ | _1435_;
	assign _0329_ = \mchip.top.receiver.fsm.state [1] & ~_0328_;
	assign _0330_ = _0329_ | \mchip.top.receiver.fsm.state [3];
	assign \mchip.top.framing_error  = _0330_ & ~_0297_;
	assign _0331_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [4] : \mchip.top.bobby.landing_fifo.queue [0]);
	assign _0332_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [12] : \mchip.top.bobby.landing_fifo.queue [8]);
	assign _0333_ = (\mchip.top.bobby.landing_fifo.get_ptr [1] ? _0332_ : _0331_);
	assign _0334_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [20] : \mchip.top.bobby.landing_fifo.queue [16]);
	assign _0335_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [28] : \mchip.top.bobby.landing_fifo.queue [24]);
	assign _0336_ = (\mchip.top.bobby.landing_fifo.get_ptr [1] ? _0335_ : _0334_);
	assign _1656_[0] = (\mchip.top.bobby.landing_fifo.get_ptr [2] ? _0336_ : _0333_);
	assign _0337_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [5] : \mchip.top.bobby.landing_fifo.queue [1]);
	assign _0338_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [13] : \mchip.top.bobby.landing_fifo.queue [9]);
	assign _0339_ = (\mchip.top.bobby.landing_fifo.get_ptr [1] ? _0338_ : _0337_);
	assign _0340_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [21] : \mchip.top.bobby.landing_fifo.queue [17]);
	assign _0341_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [29] : \mchip.top.bobby.landing_fifo.queue [25]);
	assign _0342_ = (\mchip.top.bobby.landing_fifo.get_ptr [1] ? _0341_ : _0340_);
	assign _1656_[1] = (\mchip.top.bobby.landing_fifo.get_ptr [2] ? _0342_ : _0339_);
	assign _0343_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [6] : \mchip.top.bobby.landing_fifo.queue [2]);
	assign _0344_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [14] : \mchip.top.bobby.landing_fifo.queue [10]);
	assign _0345_ = (\mchip.top.bobby.landing_fifo.get_ptr [1] ? _0344_ : _0343_);
	assign _0346_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [22] : \mchip.top.bobby.landing_fifo.queue [18]);
	assign _0347_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [30] : \mchip.top.bobby.landing_fifo.queue [26]);
	assign _0348_ = (\mchip.top.bobby.landing_fifo.get_ptr [1] ? _0347_ : _0346_);
	assign _1656_[2] = (\mchip.top.bobby.landing_fifo.get_ptr [2] ? _0348_ : _0345_);
	assign _0349_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [7] : \mchip.top.bobby.landing_fifo.queue [3]);
	assign _0350_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [15] : \mchip.top.bobby.landing_fifo.queue [11]);
	assign _0351_ = (\mchip.top.bobby.landing_fifo.get_ptr [1] ? _0350_ : _0349_);
	assign _0352_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [23] : \mchip.top.bobby.landing_fifo.queue [19]);
	assign _0353_ = (\mchip.top.bobby.landing_fifo.get_ptr [0] ? \mchip.top.bobby.landing_fifo.queue [31] : \mchip.top.bobby.landing_fifo.queue [27]);
	assign _0354_ = (\mchip.top.bobby.landing_fifo.get_ptr [1] ? _0353_ : _0352_);
	assign _1656_[3] = (\mchip.top.bobby.landing_fifo.get_ptr [2] ? _0354_ : _0351_);
	assign _0355_ = \mchip.top.receiver.conductor.clockCount [1] & \mchip.top.receiver.conductor.clockCount [0];
	assign _0356_ = _0355_ ^ \mchip.top.receiver.conductor.clockCount [2];
	assign _0041_ = _0356_ | _1434_;
	assign _0357_ = _0355_ & \mchip.top.receiver.conductor.clockCount [2];
	assign _0358_ = _0357_ ^ \mchip.top.receiver.conductor.clockCount [3];
	assign _0042_ = _0358_ | _1434_;
	assign _0359_ = ~(\mchip.top.receiver.conductor.clockCount [3] & \mchip.top.receiver.conductor.clockCount [2]);
	assign _0360_ = _0355_ & ~_0359_;
	assign _0361_ = _0360_ & \mchip.top.receiver.conductor.clockCount [4];
	assign _0362_ = _0361_ ^ \mchip.top.receiver.conductor.clockCount [5];
	assign _0043_ = _0362_ | _1434_;
	assign _0363_ = ~(\mchip.top.receiver.conductor.clockCount [4] & \mchip.top.receiver.conductor.clockCount [5]);
	assign _0364_ = _0360_ & ~_0363_;
	assign _0365_ = _0364_ ^ \mchip.top.receiver.conductor.clockCount [6];
	assign _0044_ = _0365_ | _1434_;
	assign _0203_ = (_1421_ ? \mchip.top.bobby.uart_replies.data_out [0] : \mchip.top.transmitter.saved_data [1]);
	assign _0204_ = (_1421_ ? \mchip.top.bobby.uart_replies.data_out [1] : \mchip.top.transmitter.saved_data [2]);
	assign _0205_ = (_1421_ ? \mchip.top.bobby.uart_replies.data_out [2] : \mchip.top.transmitter.saved_data [3]);
	assign _0206_ = (_1421_ ? \mchip.top.bobby.uart_replies.data_out [3] : \mchip.top.transmitter.saved_data [4]);
	assign _0207_ = (_1421_ ? \mchip.top.bobby.uart_replies.data_out [4] : \mchip.top.transmitter.saved_data [5]);
	assign _0208_ = (_1421_ ? \mchip.top.bobby.uart_replies.data_out [5] : \mchip.top.transmitter.saved_data [6]);
	assign _0209_ = (_1421_ ? \mchip.top.bobby.uart_replies.data_out [6] : \mchip.top.transmitter.saved_data [7]);
	assign _0210_ = _1421_ & \mchip.top.bobby.uart_replies.data_out [7];
	assign _0366_ = _1457_ | \mchip.top.transmitter.data_bit ;
	assign _0367_ = \mchip.top.transmitter.fsm.state [2] & ~_1430_;
	assign _0368_ = ~(\mchip.top.transmitter.fsm.state [3] | \mchip.top.transmitter.fsm.state [1]);
	assign _0369_ = _0368_ & ~\mchip.top.transmitter.fsm.state [2];
	assign _0370_ = (_0369_ ? \mchip.top.bobby.reply_fsm.state  : _0367_);
	assign _0202_ = _0366_ & ~_0370_;
	assign _0371_ = _1290_ | ~_1343_;
	assign _0372_ = _1329_ & ~_0371_;
	assign _0373_ = \mchip.top.bobby.fsm.state [5] | \mchip.top.bobby.fsm.state [4];
	assign _0374_ = _0373_ | \mchip.top.bobby.fsm.state [7];
	assign _0375_ = _0374_ | _1321_;
	assign \mchip.top.bobby.fsm.reverse_takeoff_first  = _0372_ & ~_0375_;
	assign _0376_ = (_0211_ ? \mchip.top.bobby.uart_requests.data_out [4] : \mchip.top.bobby.landing_fifo.data_out [0]);
	assign _0377_ = (_0211_ ? \mchip.top.bobby.uart_requests.data_out [5] : \mchip.top.bobby.landing_fifo.data_out [1]);
	assign _0378_ = ~(_0377_ | _0376_);
	assign _0379_ = ~\mchip.top.bobby.landing_fifo.data_out [2];
	assign _0380_ = (_0211_ ? _1293_ : _0379_);
	assign _0381_ = (_0211_ ? \mchip.top.bobby.uart_requests.data_out [7] : \mchip.top.bobby.landing_fifo.data_out [3]);
	assign _0382_ = _0381_ | ~_0380_;
	assign _0383_ = _0382_ | ~_0378_;
	assign _0384_ = _0380_ & _0378_;
	assign _0385_ = ~(_0384_ ^ _0381_);
	assign _0386_ = _0380_ ^ _0378_;
	assign _0387_ = _0377_ ^ _0376_;
	assign _0388_ = _0383_ | _0376_;
	assign _0389_ = _0388_ | _0387_;
	assign _0390_ = _0389_ | _0386_;
	assign _0391_ = _0390_ | _0385_;
	assign _0392_ = ~(_0391_ | _0383_);
	assign _0393_ = \mchip.top.bobby.id_manager.taken_id [0] & ~_0392_;
	assign _0394_ = ~\mchip.top.bobby.id_manager.taken_id [0];
	assign _0395_ = ~\mchip.top.bobby.id_manager.taken_id [1];
	assign _0396_ = ~\mchip.top.bobby.id_manager.taken_id [2];
	assign _0397_ = ~\mchip.top.bobby.id_manager.taken_id [3];
	assign _0398_ = ~\mchip.top.bobby.id_manager.taken_id [6];
	assign _0399_ = ~\mchip.top.bobby.id_manager.taken_id [7];
	assign _0400_ = ~\mchip.top.bobby.id_manager.taken_id [9];
	assign _0401_ = ~\mchip.top.bobby.id_manager.taken_id [10];
	assign _0402_ = _1589_ | ~\mchip.top.bobby.id_manager.taken_id [13];
	assign _0403_ = \mchip.top.bobby.id_manager.taken_id [12] & ~_0402_;
	assign _0404_ = ~(_0403_ & \mchip.top.bobby.id_manager.taken_id [11]);
	assign _0405_ = _0404_ | _0401_;
	assign _0406_ = _0405_ | _0400_;
	assign _0407_ = \mchip.top.bobby.id_manager.taken_id [8] & ~_0406_;
	assign _0408_ = _0407_ | _0399_;
	assign _0409_ = _0408_ | _0398_;
	assign _0410_ = \mchip.top.bobby.id_manager.taken_id [5] & ~_0409_;
	assign _0411_ = ~(_0410_ & \mchip.top.bobby.id_manager.taken_id [4]);
	assign _0412_ = _0411_ | _0397_;
	assign _0413_ = _0412_ | _0396_;
	assign _0414_ = _0413_ | _0395_;
	assign _0415_ = _0414_ | _0394_;
	assign _0416_ = _0415_ | \mchip.top.bobby.id_manager.taken_id [0];
	assign _0052_ = (_1625_ ? _0393_ : _0416_);
	assign _0417_ = ~_0385_;
	assign _0418_ = ~_0376_;
	assign _0419_ = _0383_ & ~_0418_;
	assign _0420_ = ~(_0419_ & _0387_);
	assign _0421_ = _0420_ | ~_0386_;
	assign _0422_ = _0421_ | _0417_;
	assign _0423_ = _0383_ & ~_0422_;
	assign _0424_ = \mchip.top.bobby.id_manager.taken_id [1] & ~_0423_;
	assign _0425_ = \mchip.top.bobby.id_manager.taken_id [14] & ~\mchip.top.bobby.id_manager.taken_id [15];
	assign _0426_ = \mchip.top.bobby.id_manager.taken_id [13] & ~_0425_;
	assign _0427_ = \mchip.top.bobby.id_manager.taken_id [12] & ~_0426_;
	assign _0428_ = \mchip.top.bobby.id_manager.taken_id [11] & ~_0427_;
	assign _0429_ = \mchip.top.bobby.id_manager.taken_id [10] & ~_0428_;
	assign _0430_ = \mchip.top.bobby.id_manager.taken_id [9] & ~_0429_;
	assign _0431_ = \mchip.top.bobby.id_manager.taken_id [8] & ~_0430_;
	assign _0432_ = \mchip.top.bobby.id_manager.taken_id [7] & ~_0431_;
	assign _0433_ = \mchip.top.bobby.id_manager.taken_id [6] & ~_0432_;
	assign _0434_ = \mchip.top.bobby.id_manager.taken_id [5] & ~_0433_;
	assign _0435_ = \mchip.top.bobby.id_manager.taken_id [4] & ~_0434_;
	assign _0436_ = \mchip.top.bobby.id_manager.taken_id [3] & ~_0435_;
	assign _0437_ = \mchip.top.bobby.id_manager.taken_id [2] & ~_0436_;
	assign _0438_ = \mchip.top.bobby.id_manager.taken_id [1] & ~_0437_;
	assign _0439_ = _0438_ | _0394_;
	assign _0440_ = ~\mchip.top.bobby.id_manager.taken_id [5];
	assign _0441_ = ~\mchip.top.bobby.id_manager.taken_id [11];
	assign _0442_ = ~(_1589_ & \mchip.top.bobby.id_manager.taken_id [13]);
	assign _0443_ = \mchip.top.bobby.id_manager.taken_id [12] & ~_0442_;
	assign _0444_ = _0443_ | _0441_;
	assign _0445_ = \mchip.top.bobby.id_manager.taken_id [10] & ~_0444_;
	assign _0446_ = _0445_ | _0400_;
	assign _0447_ = \mchip.top.bobby.id_manager.taken_id [8] & ~_0446_;
	assign _0448_ = _0447_ | _0399_;
	assign _0449_ = \mchip.top.bobby.id_manager.taken_id [6] & ~_0448_;
	assign _0450_ = _0449_ | _0440_;
	assign _0451_ = \mchip.top.bobby.id_manager.taken_id [4] & ~_0450_;
	assign _0452_ = _0451_ | _0397_;
	assign _0453_ = \mchip.top.bobby.id_manager.taken_id [2] & ~_0452_;
	assign _0454_ = _0453_ | _0395_;
	assign _0455_ = \mchip.top.bobby.id_manager.taken_id [0] & ~_0454_;
	assign _0456_ = _0439_ & ~_0455_;
	assign _0457_ = _0403_ | _0441_;
	assign _0458_ = _0457_ | _0401_;
	assign _0459_ = _0458_ | _0400_;
	assign _0460_ = \mchip.top.bobby.id_manager.taken_id [8] & ~_0459_;
	assign _0461_ = _0460_ | _0399_;
	assign _0462_ = _0461_ | _0398_;
	assign _0463_ = _0462_ | _0440_;
	assign _0464_ = \mchip.top.bobby.id_manager.taken_id [4] & ~_0463_;
	assign _0465_ = _0464_ | _0397_;
	assign _0466_ = _0465_ | _0396_;
	assign _0467_ = _0466_ | _0395_;
	assign _0468_ = \mchip.top.bobby.id_manager.taken_id [0] & ~_0467_;
	assign _0469_ = _0415_ & ~_0468_;
	assign _0470_ = ~(_0469_ & _0456_);
	assign _0471_ = _0455_ | _0439_;
	assign _0472_ = ~(_0468_ ^ _0456_);
	assign _0473_ = _0471_ | ~_0472_;
	assign _0474_ = _0456_ & ~_0468_;
	assign _0475_ = ~(_0474_ ^ _0415_);
	assign _0476_ = _0475_ | _0473_;
	assign _0477_ = _0470_ & ~_0476_;
	assign _0478_ = _0477_ | \mchip.top.bobby.id_manager.taken_id [1];
	assign _0059_ = (_1625_ ? _0424_ : _0478_);
	assign _0479_ = ~(_0383_ & _0418_);
	assign _0480_ = _0479_ | ~_0387_;
	assign _0481_ = _0480_ | ~_0386_;
	assign _0482_ = _0481_ | _0417_;
	assign _0483_ = _0383_ & ~_0482_;
	assign _0484_ = \mchip.top.bobby.id_manager.taken_id [2] & ~_0483_;
	assign _0485_ = ~(_0455_ & _0439_);
	assign _0486_ = _0485_ | ~_0472_;
	assign _0487_ = _0486_ | _0475_;
	assign _0488_ = _0470_ & ~_0487_;
	assign _0489_ = _0488_ | \mchip.top.bobby.id_manager.taken_id [2];
	assign _0060_ = (_1625_ ? _0484_ : _0489_);
	assign _0490_ = _0387_ | ~_0419_;
	assign _0491_ = _0490_ | ~_0386_;
	assign _0492_ = _0491_ | _0417_;
	assign _0493_ = _0383_ & ~_0492_;
	assign _0494_ = \mchip.top.bobby.id_manager.taken_id [3] & ~_0493_;
	assign _0495_ = _0439_ | ~_0455_;
	assign _0496_ = _0495_ | ~_0472_;
	assign _0497_ = _0496_ | _0475_;
	assign _0498_ = _0470_ & ~_0497_;
	assign _0499_ = _0498_ | \mchip.top.bobby.id_manager.taken_id [3];
	assign _0061_ = (_1625_ ? _0494_ : _0499_);
	assign _0500_ = _0479_ | _0387_;
	assign _0501_ = _0500_ | ~_0386_;
	assign _0502_ = _0501_ | _0417_;
	assign _0503_ = _0383_ & ~_0502_;
	assign _0504_ = \mchip.top.bobby.id_manager.taken_id [4] & ~_0503_;
	assign _0505_ = ~(_0455_ ^ _0439_);
	assign _0506_ = ~(_0470_ & _0439_);
	assign _0507_ = _0506_ | _0505_;
	assign _0508_ = _0507_ | ~_0472_;
	assign _0509_ = _0508_ | _0475_;
	assign _0510_ = _0470_ & ~_0509_;
	assign _0511_ = _0510_ | \mchip.top.bobby.id_manager.taken_id [4];
	assign _0062_ = (_1625_ ? _0504_ : _0511_);
	assign _0512_ = _0420_ | _0386_;
	assign _0513_ = _0512_ | _0417_;
	assign _0514_ = _0383_ & ~_0513_;
	assign _0515_ = \mchip.top.bobby.id_manager.taken_id [5] & ~_0514_;
	assign _0516_ = _0472_ | _0471_;
	assign _0517_ = _0516_ | _0475_;
	assign _0518_ = _0470_ & ~_0517_;
	assign _0519_ = _0518_ | \mchip.top.bobby.id_manager.taken_id [5];
	assign _0063_ = (_1625_ ? _0515_ : _0519_);
	assign _0520_ = _0480_ | _0386_;
	assign _0521_ = _0520_ | _0417_;
	assign _0522_ = _0383_ & ~_0521_;
	assign _0523_ = \mchip.top.bobby.id_manager.taken_id [6] & ~_0522_;
	assign _0524_ = _0485_ | _0472_;
	assign _0525_ = _0524_ | _0475_;
	assign _0526_ = _0470_ & ~_0525_;
	assign _0527_ = _0526_ | \mchip.top.bobby.id_manager.taken_id [6];
	assign _0064_ = (_1625_ ? _0523_ : _0527_);
	assign _0528_ = _0490_ | _0386_;
	assign _0529_ = _0528_ | _0417_;
	assign _0530_ = _0383_ & ~_0529_;
	assign _0531_ = \mchip.top.bobby.id_manager.taken_id [7] & ~_0530_;
	assign _0532_ = _0495_ | _0472_;
	assign _0533_ = _0532_ | _0475_;
	assign _0534_ = _0470_ & ~_0533_;
	assign _0535_ = _0534_ | \mchip.top.bobby.id_manager.taken_id [7];
	assign _0065_ = (_1625_ ? _0531_ : _0535_);
	assign _0536_ = _0500_ | _0386_;
	assign _0537_ = _0536_ | _0417_;
	assign _0538_ = _0383_ & ~_0537_;
	assign _0539_ = \mchip.top.bobby.id_manager.taken_id [8] & ~_0538_;
	assign _0540_ = _0507_ | _0472_;
	assign _0541_ = _0540_ | _0475_;
	assign _0542_ = _0470_ & ~_0541_;
	assign _0543_ = _0542_ | \mchip.top.bobby.id_manager.taken_id [8];
	assign _0066_ = (_1625_ ? _0539_ : _0543_);
	assign _0544_ = _0421_ | _0385_;
	assign _0545_ = _0383_ & ~_0544_;
	assign _0546_ = \mchip.top.bobby.id_manager.taken_id [9] & ~_0545_;
	assign _0547_ = _0473_ | ~_0475_;
	assign _0548_ = _0470_ & ~_0547_;
	assign _0549_ = _0548_ | \mchip.top.bobby.id_manager.taken_id [9];
	assign _0067_ = (_1625_ ? _0546_ : _0549_);
	assign _0550_ = _0481_ | _0385_;
	assign _0551_ = _0383_ & ~_0550_;
	assign _0552_ = \mchip.top.bobby.id_manager.taken_id [10] & ~_0551_;
	assign _0553_ = _0486_ | ~_0475_;
	assign _0554_ = _0470_ & ~_0553_;
	assign _0555_ = _0554_ | \mchip.top.bobby.id_manager.taken_id [10];
	assign _0053_ = (_1625_ ? _0552_ : _0555_);
	assign _0556_ = _0491_ | _0385_;
	assign _0557_ = _0383_ & ~_0556_;
	assign _0558_ = \mchip.top.bobby.id_manager.taken_id [11] & ~_0557_;
	assign _0559_ = _0496_ | ~_0475_;
	assign _0560_ = _0470_ & ~_0559_;
	assign _0561_ = _0560_ | \mchip.top.bobby.id_manager.taken_id [11];
	assign _0054_ = (_1625_ ? _0558_ : _0561_);
	assign _0562_ = _0501_ | _0385_;
	assign _0563_ = _0383_ & ~_0562_;
	assign _0564_ = \mchip.top.bobby.id_manager.taken_id [12] & ~_0563_;
	assign _0565_ = _0508_ | ~_0475_;
	assign _0566_ = _0470_ & ~_0565_;
	assign _0567_ = _0566_ | \mchip.top.bobby.id_manager.taken_id [12];
	assign _0055_ = (_1625_ ? _0564_ : _0567_);
	assign _0568_ = _0512_ | _0385_;
	assign _0569_ = _0383_ & ~_0568_;
	assign _0570_ = \mchip.top.bobby.id_manager.taken_id [13] & ~_0569_;
	assign _0571_ = _0516_ | ~_0475_;
	assign _0572_ = _0470_ & ~_0571_;
	assign _0573_ = _0572_ | \mchip.top.bobby.id_manager.taken_id [13];
	assign _0056_ = (_1625_ ? _0570_ : _0573_);
	assign _0574_ = _0520_ | _0385_;
	assign _0575_ = _0383_ & ~_0574_;
	assign _0576_ = \mchip.top.bobby.id_manager.taken_id [14] & ~_0575_;
	assign _0577_ = _0524_ | ~_0475_;
	assign _0578_ = _0470_ & ~_0577_;
	assign _0579_ = _0578_ | \mchip.top.bobby.id_manager.taken_id [14];
	assign _0057_ = (_1625_ ? _0576_ : _0579_);
	assign _0580_ = _0528_ | _0385_;
	assign _0581_ = _0383_ & ~_0580_;
	assign _0582_ = \mchip.top.bobby.id_manager.taken_id [15] & ~_0581_;
	assign _0583_ = _0532_ | ~_0475_;
	assign _0584_ = _0470_ & ~_0583_;
	assign _0585_ = _0584_ | \mchip.top.bobby.id_manager.taken_id [15];
	assign _0058_ = (_1625_ ? _0582_ : _0585_);
	assign _0586_ = (_1327_ ? \mchip.top.bobby.takeoff_fifo.data_out [0] : \mchip.top.bobby.landing_fifo.data_out [0]);
	assign _0587_ = _0218_ & ~_0439_;
	assign _0588_ = (_0211_ ? _0587_ : \mchip.top.bobby.landing_fifo.data_out [0]);
	assign _0589_ = (_0220_ ? \mchip.top.bobby.uart_requests.data_out [4] : _0588_);
	assign _0590_ = (_0225_ ? \mchip.top.bobby.uart_requests.data_out [4] : _0589_);
	assign _0591_ = (_0228_ ? \mchip.top.bobby.uart_requests.data_out [4] : _0590_);
	assign _0048_ = (_1328_ ? _0586_ : _0591_);
	assign _0592_ = (_1327_ ? \mchip.top.bobby.takeoff_fifo.data_out [1] : \mchip.top.bobby.landing_fifo.data_out [1]);
	assign _0593_ = _0455_ & _0218_;
	assign _0594_ = (_0211_ ? _0593_ : \mchip.top.bobby.landing_fifo.data_out [1]);
	assign _0595_ = (_0220_ ? \mchip.top.bobby.uart_requests.data_out [5] : _0594_);
	assign _0596_ = (_0225_ ? \mchip.top.bobby.uart_requests.data_out [5] : _0595_);
	assign _0597_ = (_0228_ ? \mchip.top.bobby.uart_requests.data_out [5] : _0596_);
	assign _0049_ = (_1328_ ? _0592_ : _0597_);
	assign _0598_ = (_1327_ ? \mchip.top.bobby.takeoff_fifo.data_out [2] : \mchip.top.bobby.landing_fifo.data_out [2]);
	assign _0599_ = _0468_ & _0218_;
	assign _0600_ = (_0211_ ? _0599_ : \mchip.top.bobby.landing_fifo.data_out [2]);
	assign _0601_ = (_0220_ ? \mchip.top.bobby.uart_requests.data_out [6] : _0600_);
	assign _0602_ = (_0225_ ? \mchip.top.bobby.uart_requests.data_out [6] : _0601_);
	assign _0603_ = (_0228_ ? \mchip.top.bobby.uart_requests.data_out [6] : _0602_);
	assign _0050_ = (_1328_ ? _0598_ : _0603_);
	assign _0604_ = (_1327_ ? \mchip.top.bobby.takeoff_fifo.data_out [3] : \mchip.top.bobby.landing_fifo.data_out [3]);
	assign _0605_ = _0218_ & ~_0415_;
	assign _0606_ = (_0211_ ? _0605_ : \mchip.top.bobby.landing_fifo.data_out [3]);
	assign _0607_ = (_0220_ ? \mchip.top.bobby.uart_requests.data_out [7] : _0606_);
	assign _0608_ = (_0225_ ? \mchip.top.bobby.uart_requests.data_out [7] : _0607_);
	assign _0609_ = (_0228_ ? \mchip.top.bobby.uart_requests.data_out [7] : _0608_);
	assign _0051_ = (_1328_ ? _0604_ : _0609_);
	assign _0610_ = _0218_ | ~_0211_;
	assign _0611_ = _0610_ | _0220_;
	assign _0612_ = _0611_ | _0225_;
	assign _0613_ = ~(_0612_ | _0228_);
	assign _0047_ = (_1328_ ? _1533_ : _0613_);
	assign _0614_ = _0211_ & ~_0220_;
	assign _0615_ = ~(_0614_ | _0225_);
	assign _0616_ = ~(_0615_ | _0228_);
	assign _0045_ = _0616_ | _1328_;
	assign _0046_ = _0229_ | _1328_;
	assign _0617_ = _1318_ | _1288_;
	assign \mchip.top.bobby.runway_manager.plane_id_lock [0] = (_0617_ ? \mchip.top.bobby.landing_fifo.data_out [0] : \mchip.top.bobby.takeoff_fifo.data_out [0]);
	assign \mchip.top.bobby.runway_manager.plane_id_lock [1] = (_0617_ ? \mchip.top.bobby.landing_fifo.data_out [1] : \mchip.top.bobby.takeoff_fifo.data_out [1]);
	assign \mchip.top.bobby.runway_manager.plane_id_lock [2] = (_0617_ ? \mchip.top.bobby.landing_fifo.data_out [2] : \mchip.top.bobby.takeoff_fifo.data_out [2]);
	assign \mchip.top.bobby.runway_manager.plane_id_lock [3] = (_0617_ ? \mchip.top.bobby.landing_fifo.data_out [3] : \mchip.top.bobby.takeoff_fifo.data_out [3]);
	assign _0618_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [8] : \mchip.top.bobby.uart_requests.queue [0]);
	assign _0619_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [24] : \mchip.top.bobby.uart_requests.queue [16]);
	assign _1659_[0] = (\mchip.top.bobby.uart_requests.get_ptr [1] ? _0619_ : _0618_);
	assign _0620_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [9] : \mchip.top.bobby.uart_requests.queue [1]);
	assign _0621_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [25] : \mchip.top.bobby.uart_requests.queue [17]);
	assign _1659_[1] = (\mchip.top.bobby.uart_requests.get_ptr [1] ? _0621_ : _0620_);
	assign _0622_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [10] : \mchip.top.bobby.uart_requests.queue [2]);
	assign _0623_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [26] : \mchip.top.bobby.uart_requests.queue [18]);
	assign _1659_[2] = (\mchip.top.bobby.uart_requests.get_ptr [1] ? _0623_ : _0622_);
	assign _0624_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [11] : \mchip.top.bobby.uart_requests.queue [3]);
	assign _0625_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [27] : \mchip.top.bobby.uart_requests.queue [19]);
	assign _1659_[3] = (\mchip.top.bobby.uart_requests.get_ptr [1] ? _0625_ : _0624_);
	assign _0626_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [12] : \mchip.top.bobby.uart_requests.queue [4]);
	assign _0627_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [28] : \mchip.top.bobby.uart_requests.queue [20]);
	assign _1659_[4] = (\mchip.top.bobby.uart_requests.get_ptr [1] ? _0627_ : _0626_);
	assign _0628_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [13] : \mchip.top.bobby.uart_requests.queue [5]);
	assign _0629_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [29] : \mchip.top.bobby.uart_requests.queue [21]);
	assign _1659_[5] = (\mchip.top.bobby.uart_requests.get_ptr [1] ? _0629_ : _0628_);
	assign _0630_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [14] : \mchip.top.bobby.uart_requests.queue [6]);
	assign _0631_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [30] : \mchip.top.bobby.uart_requests.queue [22]);
	assign _1659_[6] = (\mchip.top.bobby.uart_requests.get_ptr [1] ? _0631_ : _0630_);
	assign _0632_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [15] : \mchip.top.bobby.uart_requests.queue [7]);
	assign _0633_ = (\mchip.top.bobby.uart_requests.get_ptr [0] ? \mchip.top.bobby.uart_requests.queue [31] : \mchip.top.bobby.uart_requests.queue [23]);
	assign _1659_[7] = (\mchip.top.bobby.uart_requests.get_ptr [1] ? _0633_ : _0632_);
	assign _0634_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [8] : \mchip.top.bobby.uart_replies.queue [0]);
	assign _0635_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [24] : \mchip.top.bobby.uart_replies.queue [16]);
	assign _1658_[0] = (\mchip.top.bobby.uart_replies.get_ptr [1] ? _0635_ : _0634_);
	assign _0636_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [9] : \mchip.top.bobby.uart_replies.queue [1]);
	assign _0637_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [25] : \mchip.top.bobby.uart_replies.queue [17]);
	assign _1658_[1] = (\mchip.top.bobby.uart_replies.get_ptr [1] ? _0637_ : _0636_);
	assign _0638_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [10] : \mchip.top.bobby.uart_replies.queue [2]);
	assign _0639_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [26] : \mchip.top.bobby.uart_replies.queue [18]);
	assign _1658_[2] = (\mchip.top.bobby.uart_replies.get_ptr [1] ? _0639_ : _0638_);
	assign _0640_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [11] : \mchip.top.bobby.uart_replies.queue [3]);
	assign _0641_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [27] : \mchip.top.bobby.uart_replies.queue [19]);
	assign _1658_[3] = (\mchip.top.bobby.uart_replies.get_ptr [1] ? _0641_ : _0640_);
	assign _0642_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [12] : \mchip.top.bobby.uart_replies.queue [4]);
	assign _0643_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [28] : \mchip.top.bobby.uart_replies.queue [20]);
	assign _1658_[4] = (\mchip.top.bobby.uart_replies.get_ptr [1] ? _0643_ : _0642_);
	assign _0644_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [13] : \mchip.top.bobby.uart_replies.queue [5]);
	assign _0645_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [29] : \mchip.top.bobby.uart_replies.queue [21]);
	assign _1658_[5] = (\mchip.top.bobby.uart_replies.get_ptr [1] ? _0645_ : _0644_);
	assign _0646_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [14] : \mchip.top.bobby.uart_replies.queue [6]);
	assign _0647_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [30] : \mchip.top.bobby.uart_replies.queue [22]);
	assign _1658_[6] = (\mchip.top.bobby.uart_replies.get_ptr [1] ? _0647_ : _0646_);
	assign _0648_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [15] : \mchip.top.bobby.uart_replies.queue [7]);
	assign _0649_ = (\mchip.top.bobby.uart_replies.get_ptr [0] ? \mchip.top.bobby.uart_replies.queue [31] : \mchip.top.bobby.uart_replies.queue [23]);
	assign _1658_[7] = (\mchip.top.bobby.uart_replies.get_ptr [1] ? _0649_ : _0648_);
	assign _1635_[0] = ~\mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _1630_[0] = ~\mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _1628_[0] = ~\mchip.top.bobby.landing_fifo.get_ptr [0];
	assign _1640_[0] = ~\mchip.top.bobby.uart_replies.put_ptr [0];
	assign _1645_[0] = ~\mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1638_[0] = ~\mchip.top.bobby.uart_replies.get_ptr [0];
	assign _0650_ = _1510_ ^ \mchip.top.bobby.takeoff_fifo.count [1];
	assign _1637_[1] = _0650_ ^ \mchip.top.bobby.takeoff_fifo.count [0];
	assign _0651_ = ~(_1510_ & \mchip.top.bobby.takeoff_fifo.count [1]);
	assign _0652_ = ~(_0650_ & \mchip.top.bobby.takeoff_fifo.count [0]);
	assign _0653_ = ~(_0652_ & _0651_);
	assign _0654_ = _1510_ ^ \mchip.top.bobby.takeoff_fifo.count [2];
	assign _1637_[2] = _0654_ ^ _0653_;
	assign _0655_ = ~(_1510_ & \mchip.top.bobby.takeoff_fifo.count [2]);
	assign _0656_ = ~(_0654_ & _0653_);
	assign _0657_ = ~(_0656_ & _0655_);
	assign _0658_ = _1510_ ^ \mchip.top.bobby.takeoff_fifo.count [3];
	assign _1637_[3] = _0658_ ^ _0657_;
	assign _0659_ = ~(\mchip.top.bobby.takeoff_fifo.put_ptr [1] | \mchip.top.bobby.takeoff_fifo.put_ptr [0]);
	assign _0660_ = \mchip.top.bobby.takeoff_fifo.put_ptr [1] & \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _1636_[1] = ~(_0660_ | _0659_);
	assign _1636_[2] = _0660_ ^ \mchip.top.bobby.takeoff_fifo.put_ptr [2];
	assign _1634_[1] = \mchip.top.bobby.takeoff_fifo.get_ptr [1] ^ \mchip.top.bobby.takeoff_fifo.get_ptr [0];
	assign _0661_ = \mchip.top.bobby.takeoff_fifo.get_ptr [1] & \mchip.top.bobby.takeoff_fifo.get_ptr [0];
	assign _1634_[2] = _0661_ ^ \mchip.top.bobby.takeoff_fifo.get_ptr [2];
	assign _0662_ = _1576_ ^ \mchip.top.bobby.landing_fifo.count [1];
	assign _1632_[1] = _0662_ ^ \mchip.top.bobby.landing_fifo.count [0];
	assign _0663_ = ~(_1576_ & \mchip.top.bobby.landing_fifo.count [1]);
	assign _0664_ = ~(_0662_ & \mchip.top.bobby.landing_fifo.count [0]);
	assign _0665_ = ~(_0664_ & _0663_);
	assign _0666_ = _1576_ ^ \mchip.top.bobby.landing_fifo.count [2];
	assign _1632_[2] = _0666_ ^ _0665_;
	assign _0667_ = ~(_1576_ & \mchip.top.bobby.landing_fifo.count [2]);
	assign _0668_ = ~(_0666_ & _0665_);
	assign _0669_ = ~(_0668_ & _0667_);
	assign _0670_ = _1576_ ^ \mchip.top.bobby.landing_fifo.count [3];
	assign _1632_[3] = _0670_ ^ _0669_;
	assign _0671_ = ~(\mchip.top.bobby.landing_fifo.put_ptr [1] | \mchip.top.bobby.landing_fifo.put_ptr [0]);
	assign _0672_ = \mchip.top.bobby.landing_fifo.put_ptr [1] & \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _1631_[1] = ~(_0672_ | _0671_);
	assign _1631_[2] = _0672_ ^ \mchip.top.bobby.landing_fifo.put_ptr [2];
	assign _1653_[1] = \mchip.top.transmitter.data_counter [1] ^ \mchip.top.transmitter.data_counter [0];
	assign _0673_ = \mchip.top.transmitter.data_counter [1] & \mchip.top.transmitter.data_counter [0];
	assign _1653_[2] = _0673_ ^ \mchip.top.transmitter.data_counter [2];
	assign _0674_ = _0673_ & \mchip.top.transmitter.data_counter [2];
	assign _1653_[3] = _0674_ ^ \mchip.top.transmitter.data_counter [3];
	assign _1651_[1] = \mchip.top.receiver.conductor.clockCount [1] ^ \mchip.top.receiver.conductor.clockCount [0];
	assign _1651_[4] = _0360_ ^ \mchip.top.receiver.conductor.clockCount [4];
	assign _0675_ = _0364_ & \mchip.top.receiver.conductor.clockCount [6];
	assign _1651_[7] = _0675_ ^ \mchip.top.receiver.conductor.clockCount [7];
	assign _0676_ = _0363_ | _1393_;
	assign _0677_ = _0360_ & ~_0676_;
	assign _1651_[8] = _0677_ ^ \mchip.top.receiver.conductor.clockCount [8];
	assign _0678_ = _0677_ & \mchip.top.receiver.conductor.clockCount [8];
	assign _1651_[9] = _0678_ ^ \mchip.top.receiver.conductor.clockCount [9];
	assign _1629_[1] = \mchip.top.bobby.landing_fifo.get_ptr [1] ^ \mchip.top.bobby.landing_fifo.get_ptr [0];
	assign _0679_ = \mchip.top.bobby.landing_fifo.get_ptr [1] & \mchip.top.bobby.landing_fifo.get_ptr [0];
	assign _1629_[2] = _0679_ ^ \mchip.top.bobby.landing_fifo.get_ptr [2];
	assign _1644_[1] = \mchip.top.bobby.uart_requests.get_ptr [1] ^ \mchip.top.bobby.uart_requests.get_ptr [0];
	assign _0680_ = _1490_ ^ \mchip.top.bobby.uart_replies.count [1];
	assign _1642_[1] = _0680_ ^ \mchip.top.bobby.uart_replies.count [0];
	assign _0681_ = ~(_1490_ & \mchip.top.bobby.uart_replies.count [1]);
	assign _0682_ = ~(_0680_ & \mchip.top.bobby.uart_replies.count [0]);
	assign _0683_ = ~(_0682_ & _0681_);
	assign _0684_ = _1490_ ^ \mchip.top.bobby.uart_replies.count [2];
	assign _1642_[2] = _0684_ ^ _0683_;
	assign _0685_ = ~(\mchip.top.bobby.uart_replies.put_ptr [1] | \mchip.top.bobby.uart_replies.put_ptr [0]);
	assign _0686_ = \mchip.top.bobby.uart_replies.put_ptr [1] & \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _1641_[1] = ~(_0686_ | _0685_);
	assign _0687_ = \mchip.top.bobby.fsm.state [1] | \mchip.top.bobby.fsm.state [3];
	assign _0688_ = _1325_ & ~_0687_;
	assign _0001_ = _1333_ & ~_0688_;
	assign _0689_ = ~(_1331_ & _1333_);
	assign _0000_ = \mchip.top.bobby.fsm.state [0] & ~_0689_;
	assign _0690_ = ~_0685_;
	assign _0691_ = ~_1641_[1];
	assign _0692_ = ~(_0685_ & \mchip.top.bobby.reply_to_send [0]);
	assign _0693_ = _0692_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0694_ = _0691_ & ~_0693_;
	assign _0132_ = (_0685_ ? _0694_ : \mchip.top.bobby.uart_replies.queue [0]);
	assign _0695_ = ~(_0685_ & \mchip.top.bobby.reply_to_send [1]);
	assign _0696_ = _0695_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0697_ = _0691_ & ~_0696_;
	assign _0143_ = (_0685_ ? _0697_ : \mchip.top.bobby.uart_replies.queue [1]);
	assign _0698_ = ~(_0685_ & \mchip.top.bobby.reply_to_send [2]);
	assign _0699_ = _0698_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0700_ = _0691_ & ~_0699_;
	assign _0154_ = (_0685_ ? _0700_ : \mchip.top.bobby.uart_replies.queue [2]);
	assign _0701_ = ~(_0685_ & \mchip.top.bobby.reply_to_send [3]);
	assign _0702_ = _0701_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0703_ = _0691_ & ~_0702_;
	assign _0157_ = (_0685_ ? _0703_ : \mchip.top.bobby.uart_replies.queue [3]);
	assign _0704_ = ~(_0685_ & \mchip.top.bobby.reply_to_send [4]);
	assign _0705_ = _0704_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0706_ = _0691_ & ~_0705_;
	assign _0158_ = (_0685_ ? _0706_ : \mchip.top.bobby.uart_replies.queue [4]);
	assign _0707_ = ~(_0685_ & \mchip.top.bobby.reply_to_send [5]);
	assign _0708_ = _0707_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0709_ = _0691_ & ~_0708_;
	assign _0159_ = (_0685_ ? _0709_ : \mchip.top.bobby.uart_replies.queue [5]);
	assign _0710_ = ~(_0685_ & \mchip.top.bobby.reply_to_send [6]);
	assign _0711_ = _0710_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0712_ = _0691_ & ~_0711_;
	assign _0160_ = (_0685_ ? _0712_ : \mchip.top.bobby.uart_replies.queue [6]);
	assign _0713_ = ~(_0685_ & \mchip.top.bobby.reply_to_send [7]);
	assign _0714_ = _0713_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0715_ = _0691_ & ~_0714_;
	assign _0161_ = (_0685_ ? _0715_ : \mchip.top.bobby.uart_replies.queue [7]);
	assign _0716_ = ~(\mchip.top.bobby.reply_to_send [0] & \mchip.top.bobby.uart_replies.put_ptr [0]);
	assign _0717_ = _0716_ | ~_1641_[1];
	assign _0718_ = _0690_ & ~_0717_;
	assign _0719_ = \mchip.top.bobby.uart_replies.put_ptr [0] & ~\mchip.top.bobby.uart_replies.put_ptr [1];
	assign _0720_ = \mchip.top.bobby.uart_replies.queue [8] & ~_0719_;
	assign _0162_ = _0720_ | _0718_;
	assign _0721_ = ~(\mchip.top.bobby.reply_to_send [1] & \mchip.top.bobby.uart_replies.put_ptr [0]);
	assign _0722_ = _0721_ | ~_1641_[1];
	assign _0723_ = _0690_ & ~_0722_;
	assign _0724_ = \mchip.top.bobby.uart_replies.queue [9] & ~_0719_;
	assign _0163_ = _0724_ | _0723_;
	assign _0725_ = ~(\mchip.top.bobby.reply_to_send [2] & \mchip.top.bobby.uart_replies.put_ptr [0]);
	assign _0726_ = _0725_ | ~_1641_[1];
	assign _0727_ = _0690_ & ~_0726_;
	assign _0728_ = \mchip.top.bobby.uart_replies.queue [10] & ~_0719_;
	assign _0133_ = _0728_ | _0727_;
	assign _0729_ = ~(\mchip.top.bobby.reply_to_send [3] & \mchip.top.bobby.uart_replies.put_ptr [0]);
	assign _0730_ = _0729_ | ~_1641_[1];
	assign _0731_ = _0690_ & ~_0730_;
	assign _0732_ = \mchip.top.bobby.uart_replies.queue [11] & ~_0719_;
	assign _0134_ = _0732_ | _0731_;
	assign _0733_ = ~(\mchip.top.bobby.reply_to_send [4] & \mchip.top.bobby.uart_replies.put_ptr [0]);
	assign _0734_ = _0733_ | ~_1641_[1];
	assign _0735_ = _0690_ & ~_0734_;
	assign _0736_ = \mchip.top.bobby.uart_replies.queue [12] & ~_0719_;
	assign _0135_ = _0736_ | _0735_;
	assign _0737_ = ~(\mchip.top.bobby.reply_to_send [5] & \mchip.top.bobby.uart_replies.put_ptr [0]);
	assign _0738_ = _0737_ | ~_1641_[1];
	assign _0739_ = _0690_ & ~_0738_;
	assign _0740_ = \mchip.top.bobby.uart_replies.queue [13] & ~_0719_;
	assign _0136_ = _0740_ | _0739_;
	assign _0741_ = ~(\mchip.top.bobby.reply_to_send [6] & \mchip.top.bobby.uart_replies.put_ptr [0]);
	assign _0742_ = _0741_ | ~_1641_[1];
	assign _0743_ = _0690_ & ~_0742_;
	assign _0744_ = \mchip.top.bobby.uart_replies.queue [14] & ~_0719_;
	assign _0137_ = _0744_ | _0743_;
	assign _0745_ = ~(\mchip.top.bobby.reply_to_send [7] & \mchip.top.bobby.uart_replies.put_ptr [0]);
	assign _0746_ = _0745_ | ~_1641_[1];
	assign _0747_ = _0690_ & ~_0746_;
	assign _0748_ = \mchip.top.bobby.uart_replies.queue [15] & ~_0719_;
	assign _0138_ = _0748_ | _0747_;
	assign _0749_ = _0685_ | ~\mchip.top.bobby.reply_to_send [0];
	assign _0750_ = _0749_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0751_ = _0750_ | _0691_;
	assign _0752_ = _0690_ & ~_0751_;
	assign _0753_ = \mchip.top.bobby.uart_replies.put_ptr [1] & ~\mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0754_ = \mchip.top.bobby.uart_replies.queue [16] & ~_0753_;
	assign _0139_ = _0754_ | _0752_;
	assign _0755_ = _0685_ | ~\mchip.top.bobby.reply_to_send [1];
	assign _0756_ = _0755_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0757_ = _0756_ | _0691_;
	assign _0758_ = _0690_ & ~_0757_;
	assign _0759_ = \mchip.top.bobby.uart_replies.queue [17] & ~_0753_;
	assign _0140_ = _0759_ | _0758_;
	assign _0760_ = _0685_ | ~\mchip.top.bobby.reply_to_send [2];
	assign _0761_ = _0760_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0762_ = _0761_ | _0691_;
	assign _0763_ = _0690_ & ~_0762_;
	assign _0764_ = \mchip.top.bobby.uart_replies.queue [18] & ~_0753_;
	assign _0141_ = _0764_ | _0763_;
	assign _0765_ = _0685_ | ~\mchip.top.bobby.reply_to_send [3];
	assign _0766_ = _0765_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0767_ = _0766_ | _0691_;
	assign _0768_ = _0690_ & ~_0767_;
	assign _0769_ = \mchip.top.bobby.uart_replies.queue [19] & ~_0753_;
	assign _0142_ = _0769_ | _0768_;
	assign _0770_ = _0685_ | ~\mchip.top.bobby.reply_to_send [4];
	assign _0771_ = _0770_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0772_ = _0771_ | _0691_;
	assign _0773_ = _0690_ & ~_0772_;
	assign _0774_ = \mchip.top.bobby.uart_replies.queue [20] & ~_0753_;
	assign _0144_ = _0774_ | _0773_;
	assign _0775_ = _0685_ | ~\mchip.top.bobby.reply_to_send [5];
	assign _0776_ = _0775_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0777_ = _0776_ | _0691_;
	assign _0778_ = _0690_ & ~_0777_;
	assign _0779_ = \mchip.top.bobby.uart_replies.queue [21] & ~_0753_;
	assign _0145_ = _0779_ | _0778_;
	assign _0780_ = _0685_ | ~\mchip.top.bobby.reply_to_send [6];
	assign _0781_ = _0780_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0782_ = _0781_ | _0691_;
	assign _0783_ = _0690_ & ~_0782_;
	assign _0784_ = \mchip.top.bobby.uart_replies.queue [22] & ~_0753_;
	assign _0146_ = _0784_ | _0783_;
	assign _0785_ = _0685_ | ~\mchip.top.bobby.reply_to_send [7];
	assign _0786_ = _0785_ | \mchip.top.bobby.uart_replies.put_ptr [0];
	assign _0787_ = _0786_ | _0691_;
	assign _0788_ = _0690_ & ~_0787_;
	assign _0789_ = \mchip.top.bobby.uart_replies.queue [23] & ~_0753_;
	assign _0147_ = _0789_ | _0788_;
	assign _0790_ = _0716_ | _1641_[1];
	assign _0791_ = _0690_ & ~_0790_;
	assign _0792_ = \mchip.top.bobby.uart_replies.queue [24] & ~_0686_;
	assign _0148_ = _0792_ | _0791_;
	assign _0793_ = _0721_ | _1641_[1];
	assign _0794_ = _0690_ & ~_0793_;
	assign _0795_ = \mchip.top.bobby.uart_replies.queue [25] & ~_0686_;
	assign _0149_ = _0795_ | _0794_;
	assign _0796_ = _0725_ | _1641_[1];
	assign _0797_ = _0690_ & ~_0796_;
	assign _0798_ = \mchip.top.bobby.uart_replies.queue [26] & ~_0686_;
	assign _0150_ = _0798_ | _0797_;
	assign _0799_ = _0729_ | _1641_[1];
	assign _0800_ = _0690_ & ~_0799_;
	assign _0801_ = \mchip.top.bobby.uart_replies.queue [27] & ~_0686_;
	assign _0151_ = _0801_ | _0800_;
	assign _0802_ = _0733_ | _1641_[1];
	assign _0803_ = _0690_ & ~_0802_;
	assign _0804_ = \mchip.top.bobby.uart_replies.queue [28] & ~_0686_;
	assign _0152_ = _0804_ | _0803_;
	assign _0805_ = _0737_ | _1641_[1];
	assign _0806_ = _0690_ & ~_0805_;
	assign _0807_ = \mchip.top.bobby.uart_replies.queue [29] & ~_0686_;
	assign _0153_ = _0807_ | _0806_;
	assign _0808_ = _0741_ | _1641_[1];
	assign _0809_ = _0690_ & ~_0808_;
	assign _0810_ = \mchip.top.bobby.uart_replies.queue [30] & ~_0686_;
	assign _0155_ = _0810_ | _0809_;
	assign _0811_ = _0745_ | _1641_[1];
	assign _0812_ = _0690_ & ~_0811_;
	assign _0813_ = \mchip.top.bobby.uart_replies.queue [31] & ~_0686_;
	assign _0156_ = _0813_ | _0812_;
	assign _0814_ = _0671_ & ~\mchip.top.bobby.landing_fifo.put_ptr [2];
	assign _0815_ = ~(_0814_ & \mchip.top.bobby.uart_requests.data_out [4]);
	assign _0816_ = _0815_ | \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0817_ = _0816_ | _1631_[1];
	assign _0818_ = \mchip.top.bobby.landing_fifo.put_ptr [2] & ~_0671_;
	assign _0819_ = _0814_ & ~_0817_;
	assign _0820_ = ~(_0818_ | _0814_);
	assign _0821_ = ~(_0814_ & _1630_[0]);
	assign _0822_ = _0821_ | _1631_[1];
	assign _0823_ = _0822_ | _0820_;
	assign _0824_ = _0814_ & ~_0823_;
	assign _0825_ = \mchip.top.bobby.landing_fifo.queue [0] & ~_0824_;
	assign _0068_ = _0825_ | _0819_;
	assign _0826_ = ~(_0814_ & \mchip.top.bobby.uart_requests.data_out [5]);
	assign _0827_ = _0826_ | \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0828_ = _0827_ | _1631_[1];
	assign _0829_ = _0828_ | _0820_;
	assign _0830_ = _0814_ & ~_0829_;
	assign _0831_ = \mchip.top.bobby.landing_fifo.queue [1] & ~_0824_;
	assign _0079_ = _0831_ | _0830_;
	assign _0832_ = ~(_0814_ & \mchip.top.bobby.uart_requests.data_out [6]);
	assign _0833_ = _0832_ | \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0834_ = _0833_ | _1631_[1];
	assign _0835_ = _0834_ | _0820_;
	assign _0836_ = _0814_ & ~_0835_;
	assign _0837_ = \mchip.top.bobby.landing_fifo.queue [2] & ~_0824_;
	assign _0090_ = _0837_ | _0836_;
	assign _0838_ = ~(_0814_ & \mchip.top.bobby.uart_requests.data_out [7]);
	assign _0839_ = _0838_ | \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0840_ = _0839_ | _1631_[1];
	assign _0841_ = _0840_ | _0820_;
	assign _0842_ = _0814_ & ~_0841_;
	assign _0843_ = \mchip.top.bobby.landing_fifo.queue [3] & ~_0824_;
	assign _0093_ = _0843_ | _0842_;
	assign _0844_ = ~_0814_;
	assign _0845_ = ~(\mchip.top.bobby.landing_fifo.put_ptr [0] & \mchip.top.bobby.uart_requests.data_out [4]);
	assign _0846_ = _0845_ | ~_1631_[1];
	assign _0847_ = _0846_ | ~_0820_;
	assign _0848_ = _0844_ & ~_0847_;
	assign _0849_ = \mchip.top.bobby.landing_fifo.put_ptr [1] | ~\mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0850_ = _0849_ | ~_0820_;
	assign _0851_ = _0844_ & ~_0850_;
	assign _0852_ = \mchip.top.bobby.landing_fifo.queue [4] & ~_0851_;
	assign _0094_ = _0852_ | _0848_;
	assign _0853_ = ~(\mchip.top.bobby.landing_fifo.put_ptr [0] & \mchip.top.bobby.uart_requests.data_out [5]);
	assign _0854_ = _0853_ | ~_1631_[1];
	assign _0855_ = _0854_ | ~_0820_;
	assign _0856_ = _0844_ & ~_0855_;
	assign _0857_ = \mchip.top.bobby.landing_fifo.queue [5] & ~_0851_;
	assign _0095_ = _0857_ | _0856_;
	assign _0858_ = ~(\mchip.top.bobby.landing_fifo.put_ptr [0] & \mchip.top.bobby.uart_requests.data_out [6]);
	assign _0859_ = _0858_ | ~_1631_[1];
	assign _0860_ = _0859_ | ~_0820_;
	assign _0861_ = _0844_ & ~_0860_;
	assign _0862_ = \mchip.top.bobby.landing_fifo.queue [6] & ~_0851_;
	assign _0096_ = _0862_ | _0861_;
	assign _0863_ = ~(\mchip.top.bobby.landing_fifo.put_ptr [0] & \mchip.top.bobby.uart_requests.data_out [7]);
	assign _0864_ = _0863_ | ~_1631_[1];
	assign _0865_ = _0864_ | ~_0820_;
	assign _0866_ = _0844_ & ~_0865_;
	assign _0867_ = \mchip.top.bobby.landing_fifo.queue [7] & ~_0851_;
	assign _0097_ = _0867_ | _0866_;
	assign _0868_ = ~_0820_;
	assign _0869_ = ~_1631_[1];
	assign _0870_ = ~\mchip.top.bobby.uart_requests.data_out [4];
	assign _0871_ = _0814_ | _0870_;
	assign _0872_ = _0871_ | \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0873_ = _0872_ | _0869_;
	assign _0874_ = _0873_ | _0868_;
	assign _0875_ = _0844_ & ~_0874_;
	assign _0876_ = \mchip.top.bobby.landing_fifo.put_ptr [0] | ~\mchip.top.bobby.landing_fifo.put_ptr [1];
	assign _0877_ = _0876_ | ~_0820_;
	assign _0878_ = _0844_ & ~_0877_;
	assign _0879_ = \mchip.top.bobby.landing_fifo.queue [8] & ~_0878_;
	assign _0098_ = _0879_ | _0875_;
	assign _0880_ = _0814_ | _1294_;
	assign _0881_ = _0880_ | \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0882_ = _0881_ | _0869_;
	assign _0883_ = _0882_ | _0868_;
	assign _0884_ = _0844_ & ~_0883_;
	assign _0885_ = \mchip.top.bobby.landing_fifo.queue [9] & ~_0878_;
	assign _0099_ = _0885_ | _0884_;
	assign _0886_ = _0814_ | _1293_;
	assign _0887_ = _0886_ | \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0888_ = _0887_ | _0869_;
	assign _0889_ = _0888_ | _0868_;
	assign _0890_ = _0844_ & ~_0889_;
	assign _0891_ = \mchip.top.bobby.landing_fifo.queue [10] & ~_0878_;
	assign _0069_ = _0891_ | _0890_;
	assign _0892_ = _0814_ | _1292_;
	assign _0893_ = _0892_ | \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0894_ = _0893_ | _0869_;
	assign _0895_ = _0894_ | _0868_;
	assign _0896_ = _0844_ & ~_0895_;
	assign _0897_ = \mchip.top.bobby.landing_fifo.queue [11] & ~_0878_;
	assign _0070_ = _0897_ | _0896_;
	assign _0898_ = _0845_ | _1631_[1];
	assign _0899_ = _0898_ | ~_0820_;
	assign _0900_ = _0844_ & ~_0899_;
	assign _0901_ = ~(_0820_ & _0672_);
	assign _0902_ = _0844_ & ~_0901_;
	assign _0903_ = \mchip.top.bobby.landing_fifo.queue [12] & ~_0902_;
	assign _0071_ = _0903_ | _0900_;
	assign _0904_ = _0853_ | _1631_[1];
	assign _0905_ = _0904_ | ~_0820_;
	assign _0906_ = _0844_ & ~_0905_;
	assign _0907_ = \mchip.top.bobby.landing_fifo.queue [13] & ~_0902_;
	assign _0072_ = _0907_ | _0906_;
	assign _0908_ = _0858_ | _1631_[1];
	assign _0909_ = _0908_ | ~_0820_;
	assign _0910_ = _0844_ & ~_0909_;
	assign _0911_ = \mchip.top.bobby.landing_fifo.queue [14] & ~_0902_;
	assign _0073_ = _0911_ | _0910_;
	assign _0912_ = _0863_ | _1631_[1];
	assign _0913_ = _0912_ | ~_0820_;
	assign _0914_ = _0844_ & ~_0913_;
	assign _0915_ = \mchip.top.bobby.landing_fifo.queue [15] & ~_0902_;
	assign _0074_ = _0915_ | _0914_;
	assign _0916_ = _0872_ | _1631_[1];
	assign _0917_ = _0916_ | _0868_;
	assign _0918_ = _0844_ & ~_0917_;
	assign _0919_ = _0814_ | \mchip.top.bobby.landing_fifo.put_ptr [0];
	assign _0920_ = _0919_ | _1631_[1];
	assign _0921_ = _0920_ | _0868_;
	assign _0922_ = _0844_ & ~_0921_;
	assign _0923_ = \mchip.top.bobby.landing_fifo.queue [16] & ~_0922_;
	assign _0075_ = _0923_ | _0918_;
	assign _0924_ = _0881_ | _1631_[1];
	assign _0925_ = _0924_ | _0868_;
	assign _0926_ = _0844_ & ~_0925_;
	assign _0927_ = \mchip.top.bobby.landing_fifo.queue [17] & ~_0922_;
	assign _0076_ = _0927_ | _0926_;
	assign _0928_ = _0887_ | _1631_[1];
	assign _0929_ = _0928_ | _0868_;
	assign _0930_ = _0844_ & ~_0929_;
	assign _0931_ = \mchip.top.bobby.landing_fifo.queue [18] & ~_0922_;
	assign _0077_ = _0931_ | _0930_;
	assign _0932_ = _0893_ | _1631_[1];
	assign _0933_ = _0932_ | _0868_;
	assign _0934_ = _0844_ & ~_0933_;
	assign _0935_ = \mchip.top.bobby.landing_fifo.queue [19] & ~_0922_;
	assign _0078_ = _0935_ | _0934_;
	assign _0936_ = _0846_ | _0820_;
	assign _0937_ = _0844_ & ~_0936_;
	assign _0938_ = _0849_ | _0820_;
	assign _0939_ = _0844_ & ~_0938_;
	assign _0940_ = \mchip.top.bobby.landing_fifo.queue [20] & ~_0939_;
	assign _0080_ = _0940_ | _0937_;
	assign _0941_ = _0854_ | _0820_;
	assign _0942_ = _0844_ & ~_0941_;
	assign _0943_ = \mchip.top.bobby.landing_fifo.queue [21] & ~_0939_;
	assign _0081_ = _0943_ | _0942_;
	assign _0944_ = _0859_ | _0820_;
	assign _0945_ = _0844_ & ~_0944_;
	assign _0946_ = \mchip.top.bobby.landing_fifo.queue [22] & ~_0939_;
	assign _0082_ = _0946_ | _0945_;
	assign _0947_ = _0864_ | _0820_;
	assign _0948_ = _0844_ & ~_0947_;
	assign _0949_ = \mchip.top.bobby.landing_fifo.queue [23] & ~_0939_;
	assign _0083_ = _0949_ | _0948_;
	assign _0950_ = _0873_ | _0820_;
	assign _0951_ = _0844_ & ~_0950_;
	assign _0952_ = _0876_ | _0820_;
	assign _0953_ = _0844_ & ~_0952_;
	assign _0954_ = \mchip.top.bobby.landing_fifo.queue [24] & ~_0953_;
	assign _0084_ = _0954_ | _0951_;
	assign _0955_ = _0882_ | _0820_;
	assign _0956_ = _0844_ & ~_0955_;
	assign _0957_ = \mchip.top.bobby.landing_fifo.queue [25] & ~_0953_;
	assign _0085_ = _0957_ | _0956_;
	assign _0958_ = _0888_ | _0820_;
	assign _0959_ = _0844_ & ~_0958_;
	assign _0960_ = \mchip.top.bobby.landing_fifo.queue [26] & ~_0953_;
	assign _0086_ = _0960_ | _0959_;
	assign _0961_ = _0894_ | _0820_;
	assign _0962_ = _0844_ & ~_0961_;
	assign _0963_ = \mchip.top.bobby.landing_fifo.queue [27] & ~_0953_;
	assign _0087_ = _0963_ | _0962_;
	assign _0964_ = _0898_ | _0820_;
	assign _0965_ = _0844_ & ~_0964_;
	assign _0966_ = _0820_ | ~_0672_;
	assign _0967_ = _0844_ & ~_0966_;
	assign _0968_ = \mchip.top.bobby.landing_fifo.queue [28] & ~_0967_;
	assign _0088_ = _0968_ | _0965_;
	assign _0969_ = _0904_ | _0820_;
	assign _0970_ = _0844_ & ~_0969_;
	assign _0971_ = \mchip.top.bobby.landing_fifo.queue [29] & ~_0967_;
	assign _0089_ = _0971_ | _0970_;
	assign _0972_ = _0908_ | _0820_;
	assign _0973_ = _0844_ & ~_0972_;
	assign _0974_ = \mchip.top.bobby.landing_fifo.queue [30] & ~_0967_;
	assign _0091_ = _0974_ | _0973_;
	assign _0975_ = _0912_ | _0820_;
	assign _0976_ = _0844_ & ~_0975_;
	assign _0977_ = \mchip.top.bobby.landing_fifo.queue [31] & ~_0967_;
	assign _0092_ = _0977_ | _0976_;
	assign _0978_ = _0659_ & ~\mchip.top.bobby.takeoff_fifo.put_ptr [2];
	assign _0979_ = ~(_0978_ & \mchip.top.bobby.uart_requests.data_out [4]);
	assign _0980_ = _0979_ | \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _0981_ = _0980_ | _1636_[1];
	assign _0982_ = \mchip.top.bobby.takeoff_fifo.put_ptr [2] & ~_0659_;
	assign _0983_ = _0978_ & ~_0981_;
	assign _0984_ = ~(_0982_ | _0978_);
	assign _0985_ = ~(_0978_ & _1635_[0]);
	assign _0986_ = _0985_ | _1636_[1];
	assign _0987_ = _0986_ | _0984_;
	assign _0988_ = _0978_ & ~_0987_;
	assign _0989_ = \mchip.top.bobby.takeoff_fifo.queue [0] & ~_0988_;
	assign _0100_ = _0989_ | _0983_;
	assign _0990_ = ~(_0978_ & \mchip.top.bobby.uart_requests.data_out [5]);
	assign _0991_ = _0990_ | \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _0992_ = _0991_ | _1636_[1];
	assign _0993_ = _0992_ | _0984_;
	assign _0994_ = _0978_ & ~_0993_;
	assign _0995_ = \mchip.top.bobby.takeoff_fifo.queue [1] & ~_0988_;
	assign _0111_ = _0995_ | _0994_;
	assign _0996_ = ~(_0978_ & \mchip.top.bobby.uart_requests.data_out [6]);
	assign _0997_ = _0996_ | \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _0998_ = _0997_ | _1636_[1];
	assign _0999_ = _0998_ | _0984_;
	assign _1000_ = _0978_ & ~_0999_;
	assign _1001_ = \mchip.top.bobby.takeoff_fifo.queue [2] & ~_0988_;
	assign _0122_ = _1001_ | _1000_;
	assign _1002_ = ~(_0978_ & \mchip.top.bobby.uart_requests.data_out [7]);
	assign _1003_ = _1002_ | \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _1004_ = _1003_ | _1636_[1];
	assign _1005_ = _1004_ | _0984_;
	assign _1006_ = _0978_ & ~_1005_;
	assign _1007_ = \mchip.top.bobby.takeoff_fifo.queue [3] & ~_0988_;
	assign _0125_ = _1007_ | _1006_;
	assign _1008_ = ~_0978_;
	assign _1009_ = ~(\mchip.top.bobby.takeoff_fifo.put_ptr [0] & \mchip.top.bobby.uart_requests.data_out [4]);
	assign _1010_ = _1009_ | ~_1636_[1];
	assign _1011_ = _1010_ | ~_0984_;
	assign _1012_ = _1008_ & ~_1011_;
	assign _1013_ = \mchip.top.bobby.takeoff_fifo.put_ptr [1] | ~\mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _1014_ = _1013_ | ~_0984_;
	assign _1015_ = _1008_ & ~_1014_;
	assign _1016_ = \mchip.top.bobby.takeoff_fifo.queue [4] & ~_1015_;
	assign _0126_ = _1016_ | _1012_;
	assign _1017_ = ~(\mchip.top.bobby.takeoff_fifo.put_ptr [0] & \mchip.top.bobby.uart_requests.data_out [5]);
	assign _1018_ = _1017_ | ~_1636_[1];
	assign _1019_ = _1018_ | ~_0984_;
	assign _1020_ = _1008_ & ~_1019_;
	assign _1021_ = \mchip.top.bobby.takeoff_fifo.queue [5] & ~_1015_;
	assign _0127_ = _1021_ | _1020_;
	assign _1022_ = ~(\mchip.top.bobby.takeoff_fifo.put_ptr [0] & \mchip.top.bobby.uart_requests.data_out [6]);
	assign _1023_ = _1022_ | ~_1636_[1];
	assign _1024_ = _1023_ | ~_0984_;
	assign _1025_ = _1008_ & ~_1024_;
	assign _1026_ = \mchip.top.bobby.takeoff_fifo.queue [6] & ~_1015_;
	assign _0128_ = _1026_ | _1025_;
	assign _1027_ = ~(\mchip.top.bobby.takeoff_fifo.put_ptr [0] & \mchip.top.bobby.uart_requests.data_out [7]);
	assign _1028_ = _1027_ | ~_1636_[1];
	assign _1029_ = _1028_ | ~_0984_;
	assign _1030_ = _1008_ & ~_1029_;
	assign _1031_ = \mchip.top.bobby.takeoff_fifo.queue [7] & ~_1015_;
	assign _0129_ = _1031_ | _1030_;
	assign _1032_ = ~_0984_;
	assign _1033_ = ~_1636_[1];
	assign _1034_ = _0978_ | _0870_;
	assign _1035_ = _1034_ | \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _1036_ = _1035_ | _1033_;
	assign _1037_ = _1036_ | _1032_;
	assign _1038_ = _1008_ & ~_1037_;
	assign _1039_ = \mchip.top.bobby.takeoff_fifo.put_ptr [0] | ~\mchip.top.bobby.takeoff_fifo.put_ptr [1];
	assign _1040_ = _1039_ | ~_0984_;
	assign _1041_ = _1008_ & ~_1040_;
	assign _1042_ = \mchip.top.bobby.takeoff_fifo.queue [8] & ~_1041_;
	assign _0130_ = _1042_ | _1038_;
	assign _1043_ = _0978_ | _1294_;
	assign _1044_ = _1043_ | \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _1045_ = _1044_ | _1033_;
	assign _1046_ = _1045_ | _1032_;
	assign _1047_ = _1008_ & ~_1046_;
	assign _1048_ = \mchip.top.bobby.takeoff_fifo.queue [9] & ~_1041_;
	assign _0131_ = _1048_ | _1047_;
	assign _1049_ = _0978_ | _1293_;
	assign _1050_ = _1049_ | \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _1051_ = _1050_ | _1033_;
	assign _1052_ = _1051_ | _1032_;
	assign _1053_ = _1008_ & ~_1052_;
	assign _1054_ = \mchip.top.bobby.takeoff_fifo.queue [10] & ~_1041_;
	assign _0101_ = _1054_ | _1053_;
	assign _1055_ = _0978_ | _1292_;
	assign _1056_ = _1055_ | \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _1057_ = _1056_ | _1033_;
	assign _1058_ = _1057_ | _1032_;
	assign _1059_ = _1008_ & ~_1058_;
	assign _1060_ = \mchip.top.bobby.takeoff_fifo.queue [11] & ~_1041_;
	assign _0102_ = _1060_ | _1059_;
	assign _1061_ = _1009_ | _1636_[1];
	assign _1062_ = _1061_ | ~_0984_;
	assign _1063_ = _1008_ & ~_1062_;
	assign _1064_ = ~(_0984_ & _0660_);
	assign _1065_ = _1008_ & ~_1064_;
	assign _1066_ = \mchip.top.bobby.takeoff_fifo.queue [12] & ~_1065_;
	assign _0103_ = _1066_ | _1063_;
	assign _1067_ = _1017_ | _1636_[1];
	assign _1068_ = _1067_ | ~_0984_;
	assign _1069_ = _1008_ & ~_1068_;
	assign _1070_ = \mchip.top.bobby.takeoff_fifo.queue [13] & ~_1065_;
	assign _0104_ = _1070_ | _1069_;
	assign _1071_ = _1022_ | _1636_[1];
	assign _1072_ = _1071_ | ~_0984_;
	assign _1073_ = _1008_ & ~_1072_;
	assign _1074_ = \mchip.top.bobby.takeoff_fifo.queue [14] & ~_1065_;
	assign _0105_ = _1074_ | _1073_;
	assign _1075_ = _1027_ | _1636_[1];
	assign _1076_ = _1075_ | ~_0984_;
	assign _1077_ = _1008_ & ~_1076_;
	assign _1078_ = \mchip.top.bobby.takeoff_fifo.queue [15] & ~_1065_;
	assign _0106_ = _1078_ | _1077_;
	assign _1079_ = _1035_ | _1636_[1];
	assign _1080_ = _1079_ | _1032_;
	assign _1081_ = _1008_ & ~_1080_;
	assign _1082_ = _0978_ | \mchip.top.bobby.takeoff_fifo.put_ptr [0];
	assign _1083_ = _1082_ | _1636_[1];
	assign _1084_ = _1083_ | _1032_;
	assign _1085_ = _1008_ & ~_1084_;
	assign _1086_ = \mchip.top.bobby.takeoff_fifo.queue [16] & ~_1085_;
	assign _0107_ = _1086_ | _1081_;
	assign _1087_ = _1044_ | _1636_[1];
	assign _1088_ = _1087_ | _1032_;
	assign _1089_ = _1008_ & ~_1088_;
	assign _1090_ = \mchip.top.bobby.takeoff_fifo.queue [17] & ~_1085_;
	assign _0108_ = _1090_ | _1089_;
	assign _1091_ = _1050_ | _1636_[1];
	assign _1092_ = _1091_ | _1032_;
	assign _1093_ = _1008_ & ~_1092_;
	assign _1094_ = \mchip.top.bobby.takeoff_fifo.queue [18] & ~_1085_;
	assign _0109_ = _1094_ | _1093_;
	assign _1095_ = _1056_ | _1636_[1];
	assign _1096_ = _1095_ | _1032_;
	assign _1097_ = _1008_ & ~_1096_;
	assign _1098_ = \mchip.top.bobby.takeoff_fifo.queue [19] & ~_1085_;
	assign _0110_ = _1098_ | _1097_;
	assign _1099_ = _1010_ | _0984_;
	assign _1100_ = _1008_ & ~_1099_;
	assign _1101_ = _1013_ | _0984_;
	assign _1102_ = _1008_ & ~_1101_;
	assign _1103_ = \mchip.top.bobby.takeoff_fifo.queue [20] & ~_1102_;
	assign _0112_ = _1103_ | _1100_;
	assign _1104_ = _1018_ | _0984_;
	assign _1105_ = _1008_ & ~_1104_;
	assign _1106_ = \mchip.top.bobby.takeoff_fifo.queue [21] & ~_1102_;
	assign _0113_ = _1106_ | _1105_;
	assign _1107_ = _1023_ | _0984_;
	assign _1108_ = _1008_ & ~_1107_;
	assign _1109_ = \mchip.top.bobby.takeoff_fifo.queue [22] & ~_1102_;
	assign _0114_ = _1109_ | _1108_;
	assign _1110_ = _1028_ | _0984_;
	assign _1111_ = _1008_ & ~_1110_;
	assign _1112_ = \mchip.top.bobby.takeoff_fifo.queue [23] & ~_1102_;
	assign _0115_ = _1112_ | _1111_;
	assign _1113_ = _1036_ | _0984_;
	assign _1114_ = _1008_ & ~_1113_;
	assign _1115_ = _1039_ | _0984_;
	assign _1116_ = _1008_ & ~_1115_;
	assign _1117_ = \mchip.top.bobby.takeoff_fifo.queue [24] & ~_1116_;
	assign _0116_ = _1117_ | _1114_;
	assign _1118_ = _1045_ | _0984_;
	assign _1119_ = _1008_ & ~_1118_;
	assign _1120_ = \mchip.top.bobby.takeoff_fifo.queue [25] & ~_1116_;
	assign _0117_ = _1120_ | _1119_;
	assign _1121_ = _1051_ | _0984_;
	assign _1122_ = _1008_ & ~_1121_;
	assign _1123_ = \mchip.top.bobby.takeoff_fifo.queue [26] & ~_1116_;
	assign _0118_ = _1123_ | _1122_;
	assign _1124_ = _1057_ | _0984_;
	assign _1125_ = _1008_ & ~_1124_;
	assign _1126_ = \mchip.top.bobby.takeoff_fifo.queue [27] & ~_1116_;
	assign _0119_ = _1126_ | _1125_;
	assign _1127_ = _1061_ | _0984_;
	assign _1128_ = _1008_ & ~_1127_;
	assign _1129_ = _0984_ | ~_0660_;
	assign _1130_ = _1008_ & ~_1129_;
	assign _1131_ = \mchip.top.bobby.takeoff_fifo.queue [28] & ~_1130_;
	assign _0120_ = _1131_ | _1128_;
	assign _1132_ = _1067_ | _0984_;
	assign _1133_ = _1008_ & ~_1132_;
	assign _1134_ = \mchip.top.bobby.takeoff_fifo.queue [29] & ~_1130_;
	assign _0121_ = _1134_ | _1133_;
	assign _1135_ = _1071_ | _0984_;
	assign _1136_ = _1008_ & ~_1135_;
	assign _1137_ = \mchip.top.bobby.takeoff_fifo.queue [30] & ~_1130_;
	assign _0123_ = _1137_ | _1136_;
	assign _1138_ = _1075_ | _0984_;
	assign _1139_ = _1008_ & ~_1138_;
	assign _1140_ = \mchip.top.bobby.takeoff_fifo.queue [31] & ~_1130_;
	assign _0124_ = _1140_ | _1139_;
	assign _1141_ = ~(\mchip.top.bobby.uart_requests.put_ptr [1] | \mchip.top.bobby.uart_requests.put_ptr [0]);
	assign _1142_ = \mchip.top.bobby.uart_requests.put_ptr [1] & \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1646_[1] = ~(_1142_ | _1141_);
	assign _1143_ = ~_1141_;
	assign _1144_ = ~_1646_[1];
	assign _1145_ = ~(_1141_ & \mchip.top.receiver.data [0]);
	assign _1146_ = _1145_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1147_ = _1144_ & ~_1146_;
	assign _0164_ = (_1141_ ? _1147_ : \mchip.top.bobby.uart_requests.queue [0]);
	assign _1148_ = ~(_1141_ & \mchip.top.receiver.data [1]);
	assign _1149_ = _1148_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1150_ = _1144_ & ~_1149_;
	assign _0175_ = (_1141_ ? _1150_ : \mchip.top.bobby.uart_requests.queue [1]);
	assign _1151_ = ~(_1141_ & \mchip.top.receiver.data [2]);
	assign _1152_ = _1151_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1153_ = _1144_ & ~_1152_;
	assign _0186_ = (_1141_ ? _1153_ : \mchip.top.bobby.uart_requests.queue [2]);
	assign _1154_ = ~(_1141_ & \mchip.top.receiver.data [3]);
	assign _1155_ = _1154_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1156_ = _1144_ & ~_1155_;
	assign _0189_ = (_1141_ ? _1156_ : \mchip.top.bobby.uart_requests.queue [3]);
	assign _1157_ = ~(_1141_ & \mchip.top.receiver.data [4]);
	assign _1158_ = _1157_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1159_ = _1144_ & ~_1158_;
	assign _0190_ = (_1141_ ? _1159_ : \mchip.top.bobby.uart_requests.queue [4]);
	assign _1160_ = ~(_1141_ & \mchip.top.receiver.data [5]);
	assign _1161_ = _1160_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1162_ = _1144_ & ~_1161_;
	assign _0191_ = (_1141_ ? _1162_ : \mchip.top.bobby.uart_requests.queue [5]);
	assign _1163_ = ~(_1141_ & \mchip.top.receiver.data [6]);
	assign _1164_ = _1163_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1165_ = _1144_ & ~_1164_;
	assign _0192_ = (_1141_ ? _1165_ : \mchip.top.bobby.uart_requests.queue [6]);
	assign _1166_ = ~(_1141_ & \mchip.top.receiver.data [7]);
	assign _1167_ = _1166_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1168_ = _1144_ & ~_1167_;
	assign _0193_ = (_1141_ ? _1168_ : \mchip.top.bobby.uart_requests.queue [7]);
	assign _1169_ = ~(\mchip.top.receiver.data [0] & \mchip.top.bobby.uart_requests.put_ptr [0]);
	assign _1170_ = _1169_ | ~_1646_[1];
	assign _1171_ = _1143_ & ~_1170_;
	assign _1172_ = \mchip.top.bobby.uart_requests.put_ptr [0] & ~\mchip.top.bobby.uart_requests.put_ptr [1];
	assign _1173_ = \mchip.top.bobby.uart_requests.queue [8] & ~_1172_;
	assign _0194_ = _1173_ | _1171_;
	assign _1174_ = ~(\mchip.top.receiver.data [1] & \mchip.top.bobby.uart_requests.put_ptr [0]);
	assign _1175_ = _1174_ | ~_1646_[1];
	assign _1176_ = _1143_ & ~_1175_;
	assign _1177_ = \mchip.top.bobby.uart_requests.queue [9] & ~_1172_;
	assign _0195_ = _1177_ | _1176_;
	assign _1178_ = ~(\mchip.top.receiver.data [2] & \mchip.top.bobby.uart_requests.put_ptr [0]);
	assign _1179_ = _1178_ | ~_1646_[1];
	assign _1180_ = _1143_ & ~_1179_;
	assign _1181_ = \mchip.top.bobby.uart_requests.queue [10] & ~_1172_;
	assign _0165_ = _1181_ | _1180_;
	assign _1182_ = ~(\mchip.top.receiver.data [3] & \mchip.top.bobby.uart_requests.put_ptr [0]);
	assign _1183_ = _1182_ | ~_1646_[1];
	assign _1184_ = _1143_ & ~_1183_;
	assign _1185_ = \mchip.top.bobby.uart_requests.queue [11] & ~_1172_;
	assign _0166_ = _1185_ | _1184_;
	assign _1186_ = ~(\mchip.top.receiver.data [4] & \mchip.top.bobby.uart_requests.put_ptr [0]);
	assign _1187_ = _1186_ | ~_1646_[1];
	assign _1188_ = _1143_ & ~_1187_;
	assign _1189_ = \mchip.top.bobby.uart_requests.queue [12] & ~_1172_;
	assign _0167_ = _1189_ | _1188_;
	assign _1190_ = ~(\mchip.top.receiver.data [5] & \mchip.top.bobby.uart_requests.put_ptr [0]);
	assign _1191_ = _1190_ | ~_1646_[1];
	assign _1192_ = _1143_ & ~_1191_;
	assign _1193_ = \mchip.top.bobby.uart_requests.queue [13] & ~_1172_;
	assign _0168_ = _1193_ | _1192_;
	assign _1194_ = ~(\mchip.top.receiver.data [6] & \mchip.top.bobby.uart_requests.put_ptr [0]);
	assign _1195_ = _1194_ | ~_1646_[1];
	assign _1196_ = _1143_ & ~_1195_;
	assign _1197_ = \mchip.top.bobby.uart_requests.queue [14] & ~_1172_;
	assign _0169_ = _1197_ | _1196_;
	assign _1198_ = ~(\mchip.top.receiver.data [7] & \mchip.top.bobby.uart_requests.put_ptr [0]);
	assign _1199_ = _1198_ | ~_1646_[1];
	assign _1200_ = _1143_ & ~_1199_;
	assign _1201_ = \mchip.top.bobby.uart_requests.queue [15] & ~_1172_;
	assign _0170_ = _1201_ | _1200_;
	assign _1202_ = _1141_ | ~\mchip.top.receiver.data [0];
	assign _1203_ = _1202_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1204_ = _1203_ | _1144_;
	assign _1205_ = _1143_ & ~_1204_;
	assign _1206_ = \mchip.top.bobby.uart_requests.put_ptr [1] & ~\mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1207_ = \mchip.top.bobby.uart_requests.queue [16] & ~_1206_;
	assign _0171_ = _1207_ | _1205_;
	assign _1208_ = _1141_ | ~\mchip.top.receiver.data [1];
	assign _1209_ = _1208_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1210_ = _1209_ | _1144_;
	assign _1211_ = _1143_ & ~_1210_;
	assign _1212_ = \mchip.top.bobby.uart_requests.queue [17] & ~_1206_;
	assign _0172_ = _1212_ | _1211_;
	assign _1213_ = _1141_ | ~\mchip.top.receiver.data [2];
	assign _1214_ = _1213_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1215_ = _1214_ | _1144_;
	assign _1216_ = _1143_ & ~_1215_;
	assign _1217_ = \mchip.top.bobby.uart_requests.queue [18] & ~_1206_;
	assign _0173_ = _1217_ | _1216_;
	assign _1218_ = _1141_ | ~\mchip.top.receiver.data [3];
	assign _1219_ = _1218_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1220_ = _1219_ | _1144_;
	assign _1221_ = _1143_ & ~_1220_;
	assign _1222_ = \mchip.top.bobby.uart_requests.queue [19] & ~_1206_;
	assign _0174_ = _1222_ | _1221_;
	assign _1223_ = _1141_ | ~\mchip.top.receiver.data [4];
	assign _1224_ = _1223_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1225_ = _1224_ | _1144_;
	assign _1226_ = _1143_ & ~_1225_;
	assign _1227_ = \mchip.top.bobby.uart_requests.queue [20] & ~_1206_;
	assign _0176_ = _1227_ | _1226_;
	assign _1228_ = _1141_ | ~\mchip.top.receiver.data [5];
	assign _1229_ = _1228_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1230_ = _1229_ | _1144_;
	assign _1231_ = _1143_ & ~_1230_;
	assign _1232_ = \mchip.top.bobby.uart_requests.queue [21] & ~_1206_;
	assign _0177_ = _1232_ | _1231_;
	assign _1233_ = _1141_ | ~\mchip.top.receiver.data [6];
	assign _1234_ = _1233_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1235_ = _1234_ | _1144_;
	assign _1236_ = _1143_ & ~_1235_;
	assign _1237_ = \mchip.top.bobby.uart_requests.queue [22] & ~_1206_;
	assign _0178_ = _1237_ | _1236_;
	assign _1238_ = _1141_ | ~\mchip.top.receiver.data [7];
	assign _1239_ = _1238_ | \mchip.top.bobby.uart_requests.put_ptr [0];
	assign _1240_ = _1239_ | _1144_;
	assign _1241_ = _1143_ & ~_1240_;
	assign _1242_ = \mchip.top.bobby.uart_requests.queue [23] & ~_1206_;
	assign _0179_ = _1242_ | _1241_;
	assign _1243_ = _1169_ | _1646_[1];
	assign _1244_ = _1143_ & ~_1243_;
	assign _1245_ = \mchip.top.bobby.uart_requests.queue [24] & ~_1142_;
	assign _0180_ = _1245_ | _1244_;
	assign _1246_ = _1174_ | _1646_[1];
	assign _1247_ = _1143_ & ~_1246_;
	assign _1248_ = \mchip.top.bobby.uart_requests.queue [25] & ~_1142_;
	assign _0181_ = _1248_ | _1247_;
	assign _1249_ = _1178_ | _1646_[1];
	assign _1250_ = _1143_ & ~_1249_;
	assign _1251_ = \mchip.top.bobby.uart_requests.queue [26] & ~_1142_;
	assign _0182_ = _1251_ | _1250_;
	assign _1252_ = _1182_ | _1646_[1];
	assign _1253_ = _1143_ & ~_1252_;
	assign _1254_ = \mchip.top.bobby.uart_requests.queue [27] & ~_1142_;
	assign _0183_ = _1254_ | _1253_;
	assign _1255_ = _1186_ | _1646_[1];
	assign _1256_ = _1143_ & ~_1255_;
	assign _1257_ = \mchip.top.bobby.uart_requests.queue [28] & ~_1142_;
	assign _0184_ = _1257_ | _1256_;
	assign _1258_ = _1190_ | _1646_[1];
	assign _1259_ = _1143_ & ~_1258_;
	assign _1260_ = \mchip.top.bobby.uart_requests.queue [29] & ~_1142_;
	assign _0185_ = _1260_ | _1259_;
	assign _1261_ = _1194_ | _1646_[1];
	assign _1262_ = _1143_ & ~_1261_;
	assign _1263_ = \mchip.top.bobby.uart_requests.queue [30] & ~_1142_;
	assign _0187_ = _1263_ | _1262_;
	assign _1264_ = _1198_ | _1646_[1];
	assign _1265_ = _1143_ & ~_1264_;
	assign _1266_ = \mchip.top.bobby.uart_requests.queue [31] & ~_1142_;
	assign _0188_ = _1266_ | _1265_;
	assign _1649_[1] = \mchip.top.receiver.data_counter [1] ^ \mchip.top.receiver.data_counter [0];
	assign _1267_ = \mchip.top.receiver.data_counter [1] & \mchip.top.receiver.data_counter [0];
	assign _1649_[2] = _1267_ ^ \mchip.top.receiver.data_counter [2];
	assign _1268_ = _1267_ & \mchip.top.receiver.data_counter [2];
	assign _1649_[3] = _1268_ ^ \mchip.top.receiver.data_counter [3];
	assign _1269_ = _1476_ ^ \mchip.top.bobby.uart_requests.count [1];
	assign _1647_[1] = _1269_ ^ \mchip.top.bobby.uart_requests.count [0];
	assign _1270_ = ~(_1476_ & \mchip.top.bobby.uart_requests.count [1]);
	assign _1271_ = ~(_1269_ & \mchip.top.bobby.uart_requests.count [0]);
	assign _1272_ = ~(_1271_ & _1270_);
	assign _1273_ = _1476_ ^ \mchip.top.bobby.uart_requests.count [2];
	assign _1647_[2] = _1273_ ^ _1272_;
	assign _1655_[1] = \mchip.top.transmitter.conductor.clockCount [1] ^ \mchip.top.transmitter.conductor.clockCount [0];
	assign _1274_ = \mchip.top.transmitter.conductor.clockCount [1] & \mchip.top.transmitter.conductor.clockCount [0];
	assign _1655_[2] = _1274_ ^ \mchip.top.transmitter.conductor.clockCount [2];
	assign _1275_ = _1274_ & \mchip.top.transmitter.conductor.clockCount [2];
	assign _1655_[3] = _1275_ ^ \mchip.top.transmitter.conductor.clockCount [3];
	assign _1276_ = ~(\mchip.top.transmitter.conductor.clockCount [3] & \mchip.top.transmitter.conductor.clockCount [2]);
	assign _1277_ = _1274_ & ~_1276_;
	assign _1655_[4] = _1277_ ^ \mchip.top.transmitter.conductor.clockCount [4];
	assign _1278_ = _1277_ & \mchip.top.transmitter.conductor.clockCount [4];
	assign _1655_[5] = _1278_ ^ \mchip.top.transmitter.conductor.clockCount [5];
	assign _1279_ = ~(\mchip.top.transmitter.conductor.clockCount [4] & \mchip.top.transmitter.conductor.clockCount [5]);
	assign _1280_ = _1277_ & ~_1279_;
	assign _1655_[6] = _1280_ ^ \mchip.top.transmitter.conductor.clockCount [6];
	assign _1281_ = _1280_ & \mchip.top.transmitter.conductor.clockCount [6];
	assign _1655_[7] = _1281_ ^ \mchip.top.transmitter.conductor.clockCount [7];
	assign _1282_ = _1279_ | _1425_;
	assign _1283_ = _1277_ & ~_1282_;
	assign _1655_[8] = _1283_ ^ \mchip.top.transmitter.conductor.clockCount [8];
	assign _1284_ = _1283_ & \mchip.top.transmitter.conductor.clockCount [8];
	assign _1655_[9] = _1284_ ^ \mchip.top.transmitter.conductor.clockCount [9];
	assign _1639_[1] = \mchip.top.bobby.uart_replies.get_ptr [1] ^ \mchip.top.bobby.uart_replies.get_ptr [0];
	always @(posedge io_in[12]) \mchip.top.receiver.fsm.state [0] <= _0008_;
	always @(posedge io_in[12]) \mchip.top.receiver.fsm.state [1] <= _0009_;
	always @(posedge io_in[12]) \mchip.top.receiver.fsm.state [2] <= _0010_;
	always @(posedge io_in[12]) \mchip.top.receiver.fsm.state [3] <= _0011_;
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [0] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [0] <= _1654_[0];
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [1] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [1] <= _1655_[1];
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [2] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [2] <= _1655_[2];
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [3] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [3] <= _1655_[3];
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [4] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [4] <= _1655_[4];
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [5] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [5] <= _1655_[5];
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [6] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [6] <= _1655_[6];
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [7] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [7] <= _1655_[7];
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [8] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [8] <= _1655_[8];
	always @(posedge io_in[12])
		if (_0036_)
			\mchip.top.transmitter.conductor.clockCount [9] <= 1'h0;
		else
			\mchip.top.transmitter.conductor.clockCount [9] <= _1655_[9];
	always @(posedge io_in[12]) \mchip.top.bobby.fsm.state [0] <= _0002_;
	always @(posedge io_in[12]) \mchip.top.bobby.fsm.state [1] <= _0003_;
	always @(posedge io_in[12]) \mchip.top.bobby.fsm.state [2] <= _0004_;
	always @(posedge io_in[12]) \mchip.top.bobby.fsm.state [3] <= _0005_;
	always @(posedge io_in[12]) \mchip.top.bobby.fsm.state [4] <= _0000_;
	always @(posedge io_in[12]) \mchip.top.bobby.fsm.state [5] <= _0006_;
	always @(posedge io_in[12]) \mchip.top.bobby.fsm.state [6] <= _0007_;
	always @(posedge io_in[12]) \mchip.top.bobby.fsm.state [7] <= _0001_;
	always @(posedge io_in[12]) \mchip.top.transmitter.fsm.state [0] <= _0012_;
	always @(posedge io_in[12]) \mchip.top.transmitter.fsm.state [1] <= _0013_;
	always @(posedge io_in[12]) \mchip.top.transmitter.fsm.state [2] <= _0014_;
	always @(posedge io_in[12]) \mchip.top.transmitter.fsm.state [3] <= _0015_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [6] <= 1'h0;
		else if (_0029_)
			\mchip.top.bobby.runway_manager.runway [6] <= \mchip.top.bobby.runway_manager.plane_id_lock [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [7] <= 1'h0;
		else if (_0029_)
			\mchip.top.bobby.runway_manager.runway [7] <= \mchip.top.bobby.runway_manager.plane_id_lock [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [8] <= 1'h0;
		else if (_0029_)
			\mchip.top.bobby.runway_manager.runway [8] <= \mchip.top.bobby.runway_manager.plane_id_lock [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [9] <= 1'h0;
		else if (_0029_)
			\mchip.top.bobby.runway_manager.runway [9] <= \mchip.top.bobby.runway_manager.plane_id_lock [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [5] <= 1'h0;
		else if (_0030_)
			\mchip.top.bobby.runway_manager.runway [5] <= _0040_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [0] <= 1'h0;
		else if (_0031_)
			\mchip.top.bobby.runway_manager.runway [0] <= _0040_;
	always @(posedge io_in[12]) \mchip.top.ro_temp [0] <= io_in[1];
	always @(posedge io_in[12]) \mchip.top.ro_temp [1] <= io_in[2];
	always @(posedge io_in[12]) \mchip.top.ro_sync [0] <= \mchip.top.ro_temp [0];
	always @(posedge io_in[12]) \mchip.top.ro_sync [1] <= \mchip.top.ro_temp [1];
	always @(posedge io_in[12]) \mchip.top.eo_temp  <= io_in[3];
	always @(posedge io_in[12]) \mchip.top.eo_sync  <= \mchip.top.eo_temp ;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [0] <= _0164_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [1] <= _0175_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [2] <= _0186_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [3] <= _0189_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [4] <= _0190_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [5] <= _0191_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [6] <= _0192_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [7] <= _0193_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [8] <= _0194_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [9] <= _0195_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [10] <= _0165_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [11] <= _0166_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [12] <= _0167_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [13] <= _0168_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [14] <= _0169_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [15] <= _0170_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [16] <= _0171_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [17] <= _0172_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [18] <= _0173_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [19] <= _0174_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [20] <= _0176_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [21] <= _0177_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [22] <= _0178_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [23] <= _0179_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [24] <= _0180_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [25] <= _0181_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [26] <= _0182_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [27] <= _0183_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [28] <= _0184_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [29] <= _0185_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [30] <= _0187_;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.top.bobby.uart_requests.queue [31] <= _0188_;
	always @(posedge io_in[12])
		if (_0197_)
			\mchip.top.receiver.data_counter [0] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data_counter [0] <= _1648_[0];
	always @(posedge io_in[12])
		if (_0197_)
			\mchip.top.receiver.data_counter [1] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data_counter [1] <= _1649_[1];
	always @(posedge io_in[12])
		if (_0197_)
			\mchip.top.receiver.data_counter [2] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data_counter [2] <= _1649_[2];
	always @(posedge io_in[12])
		if (_0197_)
			\mchip.top.receiver.data_counter [3] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data_counter [3] <= _1649_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.receiver.data [0] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data [0] <= \mchip.top.receiver.data [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.receiver.data [1] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data [1] <= \mchip.top.receiver.data [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.receiver.data [2] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data [2] <= \mchip.top.receiver.data [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.receiver.data [3] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data [3] <= \mchip.top.receiver.data [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.receiver.data [4] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data [4] <= \mchip.top.receiver.data [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.receiver.data [5] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data [5] <= \mchip.top.receiver.data [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.receiver.data [6] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data [6] <= \mchip.top.receiver.data [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.receiver.data [7] <= 1'h0;
		else if (_0196_)
			\mchip.top.receiver.data [7] <= io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.transmitter.tx  <= 1'h1;
		else
			\mchip.top.transmitter.tx  <= _0202_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.transmitter.saved_data [0] <= 1'h0;
		else if (_0016_)
			\mchip.top.transmitter.saved_data [0] <= _0203_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.transmitter.saved_data [1] <= 1'h0;
		else if (_0016_)
			\mchip.top.transmitter.saved_data [1] <= _0204_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.transmitter.saved_data [2] <= 1'h0;
		else if (_0016_)
			\mchip.top.transmitter.saved_data [2] <= _0205_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.transmitter.saved_data [3] <= 1'h0;
		else if (_0016_)
			\mchip.top.transmitter.saved_data [3] <= _0206_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.transmitter.saved_data [4] <= 1'h0;
		else if (_0016_)
			\mchip.top.transmitter.saved_data [4] <= _0207_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.transmitter.saved_data [5] <= 1'h0;
		else if (_0016_)
			\mchip.top.transmitter.saved_data [5] <= _0208_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.transmitter.saved_data [6] <= 1'h0;
		else if (_0016_)
			\mchip.top.transmitter.saved_data [6] <= _0209_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.transmitter.saved_data [7] <= 1'h0;
		else if (_0016_)
			\mchip.top.transmitter.saved_data [7] <= _0210_;
	always @(posedge io_in[12])
		if (_0201_)
			\mchip.top.transmitter.data_bit  <= 1'h0;
		else if (_0199_)
			\mchip.top.transmitter.data_bit  <= \mchip.top.transmitter.saved_data [0];
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.top.receiver.conductor.clockCount [0] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [0] <= _1650_[0];
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.top.receiver.conductor.clockCount [1] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [1] <= _1651_[1];
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.top.receiver.conductor.clockCount [4] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [4] <= _1651_[4];
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.top.receiver.conductor.clockCount [7] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [7] <= _1651_[7];
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.top.receiver.conductor.clockCount [8] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [8] <= _1651_[8];
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.top.receiver.conductor.clockCount [9] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [9] <= _1651_[9];
	always @(posedge io_in[12])
		if (_0200_)
			\mchip.top.transmitter.data_counter [0] <= 1'h0;
		else if (_0199_)
			\mchip.top.transmitter.data_counter [0] <= _1652_[0];
	always @(posedge io_in[12])
		if (_0200_)
			\mchip.top.transmitter.data_counter [1] <= 1'h0;
		else if (_0199_)
			\mchip.top.transmitter.data_counter [1] <= _1653_[1];
	always @(posedge io_in[12])
		if (_0200_)
			\mchip.top.transmitter.data_counter [2] <= 1'h0;
		else if (_0199_)
			\mchip.top.transmitter.data_counter [2] <= _1653_[2];
	always @(posedge io_in[12])
		if (_0200_)
			\mchip.top.transmitter.data_counter [3] <= 1'h0;
		else if (_0199_)
			\mchip.top.transmitter.data_counter [3] <= _1653_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [1] <= 1'h0;
		else if (_0028_)
			\mchip.top.bobby.runway_manager.runway [1] <= \mchip.top.bobby.runway_manager.plane_id_lock [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [2] <= 1'h0;
		else if (_0028_)
			\mchip.top.bobby.runway_manager.runway [2] <= \mchip.top.bobby.runway_manager.plane_id_lock [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [3] <= 1'h0;
		else if (_0028_)
			\mchip.top.bobby.runway_manager.runway [3] <= \mchip.top.bobby.runway_manager.plane_id_lock [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.runway_manager.runway [4] <= 1'h0;
		else if (_0028_)
			\mchip.top.bobby.runway_manager.runway [4] <= \mchip.top.bobby.runway_manager.plane_id_lock [3];
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [0] <= _0068_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [1] <= _0079_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [2] <= _0090_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [3] <= _0093_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [4] <= _0094_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [5] <= _0095_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [6] <= _0096_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [7] <= _0097_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [8] <= _0098_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [9] <= _0099_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [10] <= _0069_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [11] <= _0070_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [12] <= _0071_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [13] <= _0072_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [14] <= _0073_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [15] <= _0074_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [16] <= _0075_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [17] <= _0076_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [18] <= _0077_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [19] <= _0078_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [20] <= _0080_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [21] <= _0081_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [22] <= _0082_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [23] <= _0083_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [24] <= _0084_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [25] <= _0085_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [26] <= _0086_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [27] <= _0087_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [28] <= _0088_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [29] <= _0089_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [30] <= _0091_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.top.bobby.landing_fifo.queue [31] <= _0092_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.data_out [0] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.data_out [0] <= _1658_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.data_out [1] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.data_out [1] <= _1658_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.data_out [2] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.data_out [2] <= _1658_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.data_out [3] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.data_out [3] <= _1658_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.data_out [4] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.data_out [4] <= _1658_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.data_out [5] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.data_out [5] <= _1658_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.data_out [6] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.data_out [6] <= _1658_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.data_out [7] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.data_out [7] <= _1658_[7];
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [0] <= _0100_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [1] <= _0111_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [2] <= _0122_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [3] <= _0125_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [4] <= _0126_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [5] <= _0127_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [6] <= _0128_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [7] <= _0129_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [8] <= _0130_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [9] <= _0131_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [10] <= _0101_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [11] <= _0102_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [12] <= _0103_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [13] <= _0104_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [14] <= _0105_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [15] <= _0106_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [16] <= _0107_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [17] <= _0108_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [18] <= _0109_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [19] <= _0110_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [20] <= _0112_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [21] <= _0113_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [22] <= _0114_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [23] <= _0115_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [24] <= _0116_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [25] <= _0117_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [26] <= _0118_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [27] <= _0119_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [28] <= _0120_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [29] <= _0121_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [30] <= _0123_;
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.top.bobby.takeoff_fifo.queue [31] <= _0124_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.count [0] <= 1'h0;
		else if (_0023_)
			\mchip.top.bobby.uart_replies.count [0] <= _1642_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.count [1] <= 1'h0;
		else if (_0023_)
			\mchip.top.bobby.uart_replies.count [1] <= _1642_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.count [2] <= 1'h0;
		else if (_0023_)
			\mchip.top.bobby.uart_replies.count [2] <= _1642_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.put_ptr [0] <= 1'h0;
		else if (_0022_)
			\mchip.top.bobby.uart_replies.put_ptr [0] <= _1640_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.put_ptr [1] <= 1'h0;
		else if (_0022_)
			\mchip.top.bobby.uart_replies.put_ptr [1] <= _1641_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.get_ptr [0] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.get_ptr [0] <= _1638_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_replies.get_ptr [1] <= 1'h0;
		else if (_1490_)
			\mchip.top.bobby.uart_replies.get_ptr [1] <= _1639_[1];
	always @(posedge io_in[12])
		if (_0198_)
			\mchip.top.receiver.conductor.clockCount [2] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [2] <= _0041_;
	always @(posedge io_in[12])
		if (_0198_)
			\mchip.top.receiver.conductor.clockCount [3] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [3] <= _0042_;
	always @(posedge io_in[12])
		if (_0198_)
			\mchip.top.receiver.conductor.clockCount [5] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [5] <= _0043_;
	always @(posedge io_in[12])
		if (_0198_)
			\mchip.top.receiver.conductor.clockCount [6] <= 1'h0;
		else
			\mchip.top.receiver.conductor.clockCount [6] <= _0044_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.fsm.takeoff_first  <= 1'h0;
		else if (\mchip.top.bobby.fsm.reverse_takeoff_first )
			\mchip.top.bobby.fsm.takeoff_first  <= _0038_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [0] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [0] <= _0052_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [1] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [1] <= _0059_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [2] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [2] <= _0060_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [3] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [3] <= _0061_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [4] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [4] <= _0062_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [5] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [5] <= _0063_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [6] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [6] <= _0064_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [7] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [7] <= _0065_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [8] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [8] <= _0066_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [9] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [9] <= _0067_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [10] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [10] <= _0053_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [11] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [11] <= _0054_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [12] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [12] <= _0055_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [13] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [13] <= _0056_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [14] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [14] <= _0057_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.id_manager.taken_id [15] <= 1'h0;
		else if (_0017_)
			\mchip.top.bobby.id_manager.taken_id [15] <= _0058_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.data_out [0] <= 1'h0;
		else if (_1576_)
			\mchip.top.bobby.landing_fifo.data_out [0] <= _1656_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.data_out [1] <= 1'h0;
		else if (_1576_)
			\mchip.top.bobby.landing_fifo.data_out [1] <= _1656_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.data_out [2] <= 1'h0;
		else if (_1576_)
			\mchip.top.bobby.landing_fifo.data_out [2] <= _1656_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.data_out [3] <= 1'h0;
		else if (_1576_)
			\mchip.top.bobby.landing_fifo.data_out [3] <= _1656_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.count [0] <= 1'h0;
		else if (_0033_)
			\mchip.top.bobby.landing_fifo.count [0] <= _1632_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.count [1] <= 1'h0;
		else if (_0033_)
			\mchip.top.bobby.landing_fifo.count [1] <= _1632_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.count [2] <= 1'h0;
		else if (_0033_)
			\mchip.top.bobby.landing_fifo.count [2] <= _1632_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.count [3] <= 1'h0;
		else if (_0033_)
			\mchip.top.bobby.landing_fifo.count [3] <= _1632_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.put_ptr [0] <= 1'h0;
		else if (_0032_)
			\mchip.top.bobby.landing_fifo.put_ptr [0] <= _1630_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.put_ptr [1] <= 1'h0;
		else if (_0032_)
			\mchip.top.bobby.landing_fifo.put_ptr [1] <= _1631_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.put_ptr [2] <= 1'h0;
		else if (_0032_)
			\mchip.top.bobby.landing_fifo.put_ptr [2] <= _1631_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.get_ptr [0] <= 1'h0;
		else if (_1576_)
			\mchip.top.bobby.landing_fifo.get_ptr [0] <= _1628_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.get_ptr [1] <= 1'h0;
		else if (_1576_)
			\mchip.top.bobby.landing_fifo.get_ptr [1] <= _1629_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.landing_fifo.get_ptr [2] <= 1'h0;
		else if (_1576_)
			\mchip.top.bobby.landing_fifo.get_ptr [2] <= _1629_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.data_out [0] <= 1'h0;
		else if (_1510_)
			\mchip.top.bobby.takeoff_fifo.data_out [0] <= _1657_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.data_out [1] <= 1'h0;
		else if (_1510_)
			\mchip.top.bobby.takeoff_fifo.data_out [1] <= _1657_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.data_out [2] <= 1'h0;
		else if (_1510_)
			\mchip.top.bobby.takeoff_fifo.data_out [2] <= _1657_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.data_out [3] <= 1'h0;
		else if (_1510_)
			\mchip.top.bobby.takeoff_fifo.data_out [3] <= _1657_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.reply_fsm.state  <= 1'h0;
		else
			\mchip.top.bobby.reply_fsm.state  <= \mchip.top.bobby.reply_fsm.next_state ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.count [0] <= 1'h0;
		else if (_0026_)
			\mchip.top.bobby.takeoff_fifo.count [0] <= _1637_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.count [1] <= 1'h0;
		else if (_0026_)
			\mchip.top.bobby.takeoff_fifo.count [1] <= _1637_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.count [2] <= 1'h0;
		else if (_0026_)
			\mchip.top.bobby.takeoff_fifo.count [2] <= _1637_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.count [3] <= 1'h0;
		else if (_0026_)
			\mchip.top.bobby.takeoff_fifo.count [3] <= _1637_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.put_ptr [0] <= 1'h0;
		else if (_0025_)
			\mchip.top.bobby.takeoff_fifo.put_ptr [0] <= _1635_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.put_ptr [1] <= 1'h0;
		else if (_0025_)
			\mchip.top.bobby.takeoff_fifo.put_ptr [1] <= _1636_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.put_ptr [2] <= 1'h0;
		else if (_0025_)
			\mchip.top.bobby.takeoff_fifo.put_ptr [2] <= _1636_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.get_ptr [0] <= 1'h0;
		else if (_1510_)
			\mchip.top.bobby.takeoff_fifo.get_ptr [0] <= _1633_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.get_ptr [1] <= 1'h0;
		else if (_1510_)
			\mchip.top.bobby.takeoff_fifo.get_ptr [1] <= _1634_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.takeoff_fifo.get_ptr [2] <= 1'h0;
		else if (_1510_)
			\mchip.top.bobby.takeoff_fifo.get_ptr [2] <= _1634_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.data_out [0] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.data_out [0] <= _1659_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.data_out [1] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.data_out [1] <= _1659_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.data_out [2] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.data_out [2] <= _1659_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.data_out [3] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.data_out [3] <= _1659_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.data_out [4] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.data_out [4] <= _1659_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.data_out [5] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.data_out [5] <= _1659_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.data_out [6] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.data_out [6] <= _1659_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.data_out [7] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.data_out [7] <= _1659_[7];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [0] <= _0132_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [1] <= _0143_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [2] <= _0154_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [3] <= _0157_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [4] <= _0158_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [5] <= _0159_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [6] <= _0160_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [7] <= _0161_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [8] <= _0162_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [9] <= _0163_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [10] <= _0133_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [11] <= _0134_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [12] <= _0135_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [13] <= _0136_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [14] <= _0137_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [15] <= _0138_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [16] <= _0139_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [17] <= _0140_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [18] <= _0141_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [19] <= _0142_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [20] <= _0144_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [21] <= _0145_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [22] <= _0146_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [23] <= _0147_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [24] <= _0148_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [25] <= _0149_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [26] <= _0150_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [27] <= _0151_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [28] <= _0152_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [29] <= _0153_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [30] <= _0155_;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.top.bobby.uart_replies.queue [31] <= _0156_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.count [0] <= 1'h0;
		else if (_0020_)
			\mchip.top.bobby.uart_requests.count [0] <= _1647_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.count [1] <= 1'h0;
		else if (_0020_)
			\mchip.top.bobby.uart_requests.count [1] <= _1647_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.count [2] <= 1'h0;
		else if (_0020_)
			\mchip.top.bobby.uart_requests.count [2] <= _1647_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.put_ptr [0] <= 1'h0;
		else if (_0019_)
			\mchip.top.bobby.uart_requests.put_ptr [0] <= _1645_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.put_ptr [1] <= 1'h0;
		else if (_0019_)
			\mchip.top.bobby.uart_requests.put_ptr [1] <= _1646_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.get_ptr [0] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.get_ptr [0] <= _1643_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.uart_requests.get_ptr [1] <= 1'h0;
		else if (_1476_)
			\mchip.top.bobby.uart_requests.get_ptr [1] <= _1644_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.reply_to_send [0] <= 1'h0;
		else if (_0035_)
			\mchip.top.bobby.reply_to_send [0] <= _0047_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.reply_to_send [1] <= 1'h0;
		else if (_0035_)
			\mchip.top.bobby.reply_to_send [1] <= _0045_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.reply_to_send [2] <= 1'h0;
		else if (_0035_)
			\mchip.top.bobby.reply_to_send [2] <= _0046_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.reply_to_send [3] <= 1'h0;
		else if (_0035_)
			\mchip.top.bobby.reply_to_send [3] <= _0039_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.reply_to_send [4] <= 1'h0;
		else if (_0035_)
			\mchip.top.bobby.reply_to_send [4] <= _0048_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.reply_to_send [5] <= 1'h0;
		else if (_0035_)
			\mchip.top.bobby.reply_to_send [5] <= _0049_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.reply_to_send [6] <= 1'h0;
		else if (_0035_)
			\mchip.top.bobby.reply_to_send [6] <= _0050_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.reply_to_send [7] <= 1'h0;
		else if (_0035_)
			\mchip.top.bobby.reply_to_send [7] <= _0051_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.emergency_id [0] <= 1'h0;
		else if (\mchip.top.bobby.fsm.set_emergency )
			\mchip.top.bobby.emergency_id [0] <= \mchip.top.bobby.uart_requests.data_out [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.emergency_id [1] <= 1'h0;
		else if (\mchip.top.bobby.fsm.set_emergency )
			\mchip.top.bobby.emergency_id [1] <= \mchip.top.bobby.uart_requests.data_out [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.emergency_id [2] <= 1'h0;
		else if (\mchip.top.bobby.fsm.set_emergency )
			\mchip.top.bobby.emergency_id [2] <= \mchip.top.bobby.uart_requests.data_out [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.emergency_id [3] <= 1'h0;
		else if (\mchip.top.bobby.fsm.set_emergency )
			\mchip.top.bobby.emergency_id [3] <= \mchip.top.bobby.uart_requests.data_out [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.bobby.emergency  <= 1'h0;
		else if (_0018_)
			\mchip.top.bobby.emergency  <= \mchip.top.bobby.fsm.set_emergency ;
	assign _1628_[2:1] = \mchip.top.bobby.landing_fifo.get_ptr [2:1];
	assign _1629_[0] = _1628_[0];
	assign _1630_[2:1] = \mchip.top.bobby.landing_fifo.put_ptr [2:1];
	assign _1631_[0] = _1630_[0];
	assign _1633_[2:1] = \mchip.top.bobby.takeoff_fifo.get_ptr [2:1];
	assign _1634_[0] = _1633_[0];
	assign _1635_[2:1] = \mchip.top.bobby.takeoff_fifo.put_ptr [2:1];
	assign _1636_[0] = _1635_[0];
	assign _1638_[1] = \mchip.top.bobby.uart_replies.get_ptr [1];
	assign _1639_[0] = _1638_[0];
	assign _1640_[1] = \mchip.top.bobby.uart_replies.put_ptr [1];
	assign _1641_[0] = _1640_[0];
	assign _1643_[1] = \mchip.top.bobby.uart_requests.get_ptr [1];
	assign _1644_[0] = _1643_[0];
	assign _1645_[1] = \mchip.top.bobby.uart_requests.put_ptr [1];
	assign _1646_[0] = _1645_[0];
	assign _1648_[3:1] = \mchip.top.receiver.data_counter [3:1];
	assign _1649_[0] = _1648_[0];
	assign _1650_[9:1] = \mchip.top.receiver.conductor.clockCount [9:1];
	assign {_1651_[6:5], _1651_[3:2], _1651_[0]} = {4'h0, _1650_[0]};
	assign _1652_[3:1] = \mchip.top.transmitter.data_counter [3:1];
	assign _1653_[0] = _1652_[0];
	assign _1654_[9:1] = \mchip.top.transmitter.conductor.clockCount [9:1];
	assign _1655_[0] = _1654_[0];
	assign {io_out[13:4], io_out[1:0]} = {7'h00, \mchip.top.sending , \mchip.top.receiver.fsm.receiving , \mchip.top.bobby.emergency_out , \mchip.top.framing_error , \mchip.top.transmitter.tx };
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {5'h00, \mchip.top.sending , \mchip.top.receiver.fsm.receiving , \mchip.top.bobby.emergency_out , io_out[3:2], \mchip.top.framing_error , \mchip.top.transmitter.tx };
	assign \mchip.reset  = io_in[13];
	assign \mchip.top.bobby.all_id  = \mchip.top.bobby.id_manager.taken_id ;
	assign \mchip.top.bobby.cleared_id_to_lock  = \mchip.top.bobby.runway_manager.plane_id_lock ;
	assign \mchip.top.bobby.cleared_landing_id  = \mchip.top.bobby.landing_fifo.data_out ;
	assign \mchip.top.bobby.cleared_takeoff_id  = \mchip.top.bobby.takeoff_fifo.data_out ;
	assign \mchip.top.bobby.clock  = io_in[12];
	assign \mchip.top.bobby.emergency_override  = \mchip.top.eo_sync ;
	assign \mchip.top.bobby.fsm.all_id  = \mchip.top.bobby.id_manager.taken_id ;
	assign \mchip.top.bobby.fsm.clock  = io_in[12];
	assign \mchip.top.bobby.fsm.emergency  = \mchip.top.bobby.emergency_out ;
	assign \mchip.top.bobby.fsm.emergency_id  = \mchip.top.bobby.emergency_id ;
	assign \mchip.top.bobby.fsm.msg_action  = {1'h0, \mchip.top.bobby.uart_requests.data_out [0]};
	assign \mchip.top.bobby.fsm.msg_type  = \mchip.top.bobby.uart_requests.data_out [3:1];
	assign \mchip.top.bobby.fsm.plane_id  = \mchip.top.bobby.uart_requests.data_out [7:4];
	assign \mchip.top.bobby.fsm.reset  = io_in[13];
	assign \mchip.top.bobby.fsm.runway  = \mchip.top.bobby.runway_manager.runway ;
	assign \mchip.top.bobby.fsm.runway_active  = io_out[3:2];
	assign \mchip.top.bobby.fsm.uart_request  = \mchip.top.bobby.uart_requests.data_out ;
	assign \mchip.top.bobby.id_manager.all_id  = \mchip.top.bobby.id_manager.taken_id ;
	assign \mchip.top.bobby.id_manager.clock  = io_in[12];
	assign \mchip.top.bobby.id_manager.reset  = io_in[13];
	assign \mchip.top.bobby.landing_fifo.clock  = io_in[12];
	assign \mchip.top.bobby.landing_fifo.data_in  = \mchip.top.bobby.uart_requests.data_out [7:4];
	assign \mchip.top.bobby.landing_fifo.reset  = io_in[13];
	assign \mchip.top.bobby.reply_fsm.clock  = io_in[12];
	assign \mchip.top.bobby.reply_fsm.reset  = io_in[13];
	assign \mchip.top.bobby.reply_fsm.send_reply  = \mchip.top.bobby.reply_fsm.next_state ;
	assign \mchip.top.bobby.reply_fsm.uart_tx_send  = \mchip.top.bobby.reply_fsm.state ;
	assign \mchip.top.bobby.reset  = io_in[13];
	assign \mchip.top.bobby.runway  = \mchip.top.bobby.runway_manager.runway ;
	assign \mchip.top.bobby.runway_active  = io_out[3:2];
	assign \mchip.top.bobby.runway_manager.clock  = io_in[12];
	assign \mchip.top.bobby.runway_manager.plane_id_unlock  = \mchip.top.bobby.uart_requests.data_out [7:4];
	assign \mchip.top.bobby.runway_manager.reset  = io_in[13];
	assign \mchip.top.bobby.runway_manager.runway_active  = io_out[3:2];
	assign \mchip.top.bobby.runway_manager.runway_override  = \mchip.top.ro_sync ;
	assign \mchip.top.bobby.runway_override  = \mchip.top.ro_sync ;
	assign \mchip.top.bobby.send_reply  = \mchip.top.bobby.reply_fsm.next_state ;
	assign \mchip.top.bobby.set_emergency  = \mchip.top.bobby.fsm.set_emergency ;
	assign \mchip.top.bobby.takeoff_fifo.clock  = io_in[12];
	assign \mchip.top.bobby.takeoff_fifo.data_in  = \mchip.top.bobby.uart_requests.data_out [7:4];
	assign \mchip.top.bobby.takeoff_fifo.reset  = io_in[13];
	assign \mchip.top.bobby.uart_replies.clock  = io_in[12];
	assign \mchip.top.bobby.uart_replies.data_in  = \mchip.top.bobby.reply_to_send ;
	assign \mchip.top.bobby.uart_replies.re  = \mchip.top.bobby.reply_fsm.next_state ;
	assign \mchip.top.bobby.uart_replies.reset  = io_in[13];
	assign \mchip.top.bobby.uart_request  = \mchip.top.bobby.uart_requests.data_out ;
	assign \mchip.top.bobby.uart_requests.clock  = io_in[12];
	assign \mchip.top.bobby.uart_requests.data_in  = \mchip.top.receiver.data ;
	assign \mchip.top.bobby.uart_requests.reset  = io_in[13];
	assign \mchip.top.bobby.uart_rx_data  = \mchip.top.receiver.data ;
	assign \mchip.top.bobby.uart_tx_data  = \mchip.top.bobby.uart_replies.data_out ;
	assign \mchip.top.bobby.uart_tx_send  = \mchip.top.bobby.reply_fsm.state ;
	assign \mchip.top.clock  = io_in[12];
	assign \mchip.top.emergency  = \mchip.top.bobby.emergency_out ;
	assign \mchip.top.emergency_override  = io_in[3];
	assign \mchip.top.receiver.clock  = io_in[12];
	assign \mchip.top.receiver.conductor.clock  = io_in[12];
	assign \mchip.top.receiver.conductor.reset  = io_in[13];
	assign \mchip.top.receiver.conductor.start_tx  = 1'h0;
	assign \mchip.top.receiver.framing_error  = \mchip.top.framing_error ;
	assign \mchip.top.receiver.fsm.clock  = io_in[12];
	assign \mchip.top.receiver.fsm.framing_error  = \mchip.top.framing_error ;
	assign \mchip.top.receiver.fsm.reset  = io_in[13];
	assign \mchip.top.receiver.fsm.rx  = io_in[0];
	assign \mchip.top.receiver.receiving  = \mchip.top.receiver.fsm.receiving ;
	assign \mchip.top.receiver.reset  = io_in[13];
	assign \mchip.top.receiver.rx  = io_in[0];
	assign \mchip.top.receiving  = \mchip.top.receiver.fsm.receiving ;
	assign \mchip.top.reset  = io_in[13];
	assign \mchip.top.runway_active  = io_out[3:2];
	assign \mchip.top.runway_override  = io_in[2:1];
	assign \mchip.top.rx  = io_in[0];
	assign \mchip.top.transmitter.clock  = io_in[12];
	assign \mchip.top.transmitter.conductor.clock  = io_in[12];
	assign \mchip.top.transmitter.conductor.reset  = io_in[13];
	assign \mchip.top.transmitter.conductor.start_rx  = 1'h0;
	assign \mchip.top.transmitter.data  = \mchip.top.bobby.uart_replies.data_out ;
	assign \mchip.top.transmitter.fsm.clock  = io_in[12];
	assign \mchip.top.transmitter.fsm.reset  = io_in[13];
	assign \mchip.top.transmitter.fsm.send  = \mchip.top.bobby.reply_fsm.state ;
	assign \mchip.top.transmitter.fsm.sending  = \mchip.top.sending ;
	assign \mchip.top.transmitter.reset  = io_in[13];
	assign \mchip.top.transmitter.send  = \mchip.top.bobby.reply_fsm.state ;
	assign \mchip.top.transmitter.sending  = \mchip.top.sending ;
	assign \mchip.top.tx  = \mchip.top.transmitter.tx ;
	assign \mchip.top.uart_rx_data  = \mchip.top.receiver.data ;
	assign \mchip.top.uart_tx_data  = \mchip.top.bobby.uart_replies.data_out ;
	assign \mchip.top.uart_tx_send  = \mchip.top.bobby.reply_fsm.state ;
endmodule
module d17_cporco_clockbox (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire [18:0] _1321_;
	wire [18:0] _1322_;
	wire [29:0] _1323_;
	wire [23:0] _1324_;
	wire [23:0] _1325_;
	wire [3:0] _1326_;
	wire [3:0] _1327_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.blink_drive ;
	reg [18:0] \mchip.button_count ;
	reg [23:0] \mchip.chrono_count ;
	reg [3:0] \mchip.chrono_time0 ;
	reg [3:0] \mchip.chrono_time1 ;
	reg [3:0] \mchip.chrono_time2 ;
	reg [3:0] \mchip.chrono_time3 ;
	wire \mchip.clock ;
	reg [29:0] \mchip.clock_count ;
	reg [1:0] \mchip.clock_digit_sel ;
	reg [3:0] \mchip.clock_time0 ;
	reg [3:0] \mchip.clock_time1 ;
	reg [3:0] \mchip.clock_time2 ;
	reg [3:0] \mchip.clock_time3 ;
	reg [2:0] \mchip.cur_state ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.leddrive0.blink ;
	wire [1:0] \mchip.leddrive0.blink_sel ;
	wire [4:0] \mchip.leddrive0.cd0.col0 ;
	wire [4:0] \mchip.leddrive0.cd0.col1 ;
	wire [4:0] \mchip.leddrive0.cd0.col2 ;
	wire [4:0] \mchip.leddrive0.cd1.col0 ;
	wire [4:0] \mchip.leddrive0.cd1.col1 ;
	wire [4:0] \mchip.leddrive0.cd1.col2 ;
	wire [4:0] \mchip.leddrive0.cd2.col0 ;
	wire [4:0] \mchip.leddrive0.cd2.col1 ;
	wire [4:0] \mchip.leddrive0.cd2.col2 ;
	wire [4:0] \mchip.leddrive0.cd3.col0 ;
	wire [4:0] \mchip.leddrive0.cd3.col1 ;
	wire [4:0] \mchip.leddrive0.cd3.col2 ;
	wire \mchip.leddrive0.clock ;
	reg [3:0] \mchip.leddrive0.col_sel ;
	wire [10:0] \mchip.leddrive0.colcount0.D ;
	reg [10:0] \mchip.leddrive0.colcount0.Q ;
	wire \mchip.leddrive0.colcount0.clock ;
	wire \mchip.leddrive0.colcount0.en ;
	wire \mchip.leddrive0.colcount0.reset ;
	wire [4:0] \mchip.leddrive0.dig0col0 ;
	wire [4:0] \mchip.leddrive0.dig0col1 ;
	wire [4:0] \mchip.leddrive0.dig0col2 ;
	wire [4:0] \mchip.leddrive0.dig1col0 ;
	wire [4:0] \mchip.leddrive0.dig1col1 ;
	wire [4:0] \mchip.leddrive0.dig1col2 ;
	wire [4:0] \mchip.leddrive0.dig2col0 ;
	wire [4:0] \mchip.leddrive0.dig2col1 ;
	wire [4:0] \mchip.leddrive0.dig2col2 ;
	wire [4:0] \mchip.leddrive0.dig3col0 ;
	wire [4:0] \mchip.leddrive0.dig3col1 ;
	wire [4:0] \mchip.leddrive0.dig3col2 ;
	wire [10:0] \mchip.leddrive0.in_colcount ;
	reg [23:0] \mchip.leddrive0.out_clockcount ;
	wire [10:0] \mchip.leddrive0.out_colcount ;
	reg [5:0] \mchip.leddrive0.power_mode ;
	wire \mchip.leddrive0.reset ;
	wire \mchip.leddrive0.reset_colcount ;
	wire [4:0] \mchip.leddrive0.row_L ;
	reg \mchip.mode_bounce ;
	reg \mchip.mode_buf ;
	reg \mchip.mode_tmp0 ;
	reg \mchip.mode_tmp1 ;
	wire \mchip.modehold0.button ;
	reg \mchip.modehold0.button_latched ;
	reg [2:0] \mchip.modehold0.button_state ;
	wire [24:0] \mchip.modehold0.buttoncount.D ;
	reg [24:0] \mchip.modehold0.buttoncount.Q ;
	wire \mchip.modehold0.buttoncount.clock ;
	wire \mchip.modehold0.buttoncount.en ;
	wire \mchip.modehold0.buttoncount.reset ;
	wire \mchip.modehold0.clear_buttoncount ;
	wire \mchip.modehold0.clock ;
	wire \mchip.modehold0.en_buttoncount ;
	wire \mchip.modehold0.en_buttonlatch ;
	wire [24:0] \mchip.modehold0.in_buttoncount ;
	wire [24:0] \mchip.modehold0.out_buttoncount ;
	wire \mchip.modehold0.reset ;
	wire \mchip.modehold0.reset_buttoncount ;
	reg \mchip.pm ;
	reg \mchip.power_bounce ;
	reg \mchip.power_buf ;
	reg \mchip.power_state ;
	wire \mchip.power_state_next ;
	reg \mchip.power_tmp0 ;
	reg \mchip.power_tmp1 ;
	wire \mchip.reset ;
	reg \mchip.run_chrono ;
	reg \mchip.start_bounce ;
	reg \mchip.start_buf ;
	reg \mchip.start_state ;
	wire \mchip.start_state_next ;
	reg \mchip.start_tmp0 ;
	reg \mchip.start_tmp1 ;
	reg \mchip.stop_bounce ;
	reg \mchip.stop_buf ;
	reg \mchip.stop_tmp0 ;
	reg \mchip.stop_tmp1 ;
	wire \mchip.stophold0.button ;
	reg \mchip.stophold0.button_latched ;
	reg [2:0] \mchip.stophold0.button_state ;
	wire [24:0] \mchip.stophold0.buttoncount.D ;
	reg [24:0] \mchip.stophold0.buttoncount.Q ;
	wire \mchip.stophold0.buttoncount.clock ;
	wire \mchip.stophold0.buttoncount.en ;
	wire \mchip.stophold0.buttoncount.reset ;
	wire \mchip.stophold0.clear_buttoncount ;
	wire \mchip.stophold0.clock ;
	wire \mchip.stophold0.en_buttoncount ;
	wire \mchip.stophold0.en_buttonlatch ;
	wire [24:0] \mchip.stophold0.in_buttoncount ;
	wire [24:0] \mchip.stophold0.out_buttoncount ;
	wire \mchip.stophold0.reset ;
	wire \mchip.stophold0.reset_buttoncount ;
	assign _0922_ = _0921_ | _0920_;
	assign _0923_ = _0922_ | _0919_;
	assign _0924_ = \mchip.chrono_count [14] | ~\mchip.chrono_count [15];
	assign _0925_ = \mchip.chrono_count [13] | ~\mchip.chrono_count [12];
	assign _0926_ = _0925_ | _0924_;
	assign _0927_ = \mchip.chrono_count [11] | ~\mchip.chrono_count [10];
	assign _0928_ = \mchip.chrono_count [8] | ~\mchip.chrono_count [9];
	assign _0929_ = _0928_ | _0927_;
	assign _0930_ = _0929_ | _0926_;
	assign _0931_ = \mchip.chrono_count [6] | ~\mchip.chrono_count [7];
	assign _0932_ = \mchip.chrono_count [4] | \mchip.chrono_count [5];
	assign _0933_ = _0932_ | _0931_;
	assign _0934_ = \mchip.chrono_count [2] | \mchip.chrono_count [3];
	assign _0935_ = \mchip.chrono_count [0] | \mchip.chrono_count [1];
	assign _0936_ = _0935_ | _0934_;
	assign _0937_ = _0936_ | _0933_;
	assign _0938_ = _0937_ | _0930_;
	assign _0939_ = _0938_ | _0923_;
	assign _0940_ = \mchip.run_chrono  & ~_0939_;
	assign _0941_ = \mchip.chrono_time0 [3] & ~\mchip.chrono_time0 [2];
	assign _0942_ = \mchip.chrono_time0 [0] & ~\mchip.chrono_time0 [1];
	assign _0943_ = _0942_ & _0941_;
	assign _0944_ = \mchip.chrono_time1 [2] & ~\mchip.chrono_time1 [3];
	assign _0945_ = \mchip.chrono_time1 [0] & ~\mchip.chrono_time1 [1];
	assign _0946_ = _0945_ & _0944_;
	assign _0947_ = ~(_0946_ & _0943_);
	assign _0948_ = \mchip.chrono_time2 [3] & ~\mchip.chrono_time2 [2];
	assign _0949_ = \mchip.chrono_time2 [0] & ~\mchip.chrono_time2 [1];
	assign _0950_ = _0949_ & _0948_;
	assign _0951_ = ~_0950_;
	assign _0952_ = _0951_ | _0031_;
	assign _0953_ = _0952_ | _0947_;
	assign _0019_ = _0940_ & ~_0953_;
	assign _0954_ = ~_0943_;
	assign _0955_ = _0954_ | _0939_;
	assign _0956_ = ~_0946_;
	assign _0957_ = _0956_ | _0031_;
	assign _0958_ = _0957_ | _0955_;
	assign _0020_ = \mchip.run_chrono  & ~_0958_;
	assign _0959_ = ~(\mchip.stophold0.buttoncount.Q [22] | \mchip.stophold0.buttoncount.Q [23]);
	assign _0960_ = ~(\mchip.stophold0.buttoncount.Q [20] & \mchip.stophold0.buttoncount.Q [21]);
	assign _0961_ = _0959_ & ~_0960_;
	assign _0962_ = \mchip.stophold0.buttoncount.Q [18] | \mchip.stophold0.buttoncount.Q [19];
	assign _0963_ = ~(_0962_ | \mchip.stophold0.buttoncount.Q [17]);
	assign _0964_ = _0961_ & ~_0963_;
	assign _0965_ = _0959_ & ~_0964_;
	assign _0966_ = \mchip.stophold0.buttoncount.Q [17] | ~\mchip.stophold0.buttoncount.Q [16];
	assign _0967_ = _0966_ | _0962_;
	assign _0968_ = _0961_ & ~_0967_;
	assign _0969_ = ~(\mchip.stophold0.buttoncount.Q [14] | \mchip.stophold0.buttoncount.Q [15]);
	assign _0970_ = \mchip.stophold0.buttoncount.Q [13] & \mchip.stophold0.buttoncount.Q [12];
	assign _0971_ = _0969_ & ~_0970_;
	assign _0972_ = \mchip.stophold0.buttoncount.Q [12] | ~\mchip.stophold0.buttoncount.Q [13];
	assign _0973_ = _0969_ & ~_0972_;
	assign _0974_ = ~(\mchip.stophold0.buttoncount.Q [8] | \mchip.stophold0.buttoncount.Q [9]);
	assign _0975_ = ~(\mchip.stophold0.buttoncount.Q [10] & \mchip.stophold0.buttoncount.Q [11]);
	assign _0976_ = _0975_ | _0974_;
	assign _0977_ = _0973_ & ~_0976_;
	assign _0978_ = _0971_ & ~_0977_;
	assign _0979_ = _0968_ & ~_0978_;
	assign _0980_ = _0965_ & ~_0979_;
	assign _0981_ = \mchip.stophold0.buttoncount.Q [24] & ~_0980_;
	assign _0982_ = ~(\mchip.stophold0.buttoncount.Q [1] | \mchip.stophold0.buttoncount.Q [0]);
	assign _0983_ = \mchip.stophold0.buttoncount.Q [2] | \mchip.stophold0.buttoncount.Q [3];
	assign _0984_ = _0982_ & ~_0983_;
	assign _0985_ = \mchip.stophold0.buttoncount.Q [6] | \mchip.stophold0.buttoncount.Q [7];
	assign _0986_ = \mchip.stophold0.buttoncount.Q [4] | \mchip.stophold0.buttoncount.Q [5];
	assign _0987_ = _0986_ | _0985_;
	assign _0988_ = _0984_ & ~_0987_;
	assign _0989_ = \mchip.stophold0.buttoncount.Q [9] | ~\mchip.stophold0.buttoncount.Q [8];
	assign _0990_ = ~(_0989_ | _0975_);
	assign _0991_ = ~(_0990_ & _0973_);
	assign _0992_ = _0988_ & ~_0991_;
	assign _0993_ = ~(_0968_ & \mchip.stophold0.buttoncount.Q [24]);
	assign _0994_ = _0992_ & ~_0993_;
	assign \mchip.stophold0.en_buttonlatch  = _0994_ | _0981_;
	assign _0995_ = _0954_ | _0031_;
	assign _0021_ = _0940_ & ~_0995_;
	assign \mchip.modehold0.buttoncount.D [0] = ~\mchip.modehold0.buttoncount.Q [0];
	assign _0996_ = _0939_ | _0031_;
	assign _0022_ = \mchip.run_chrono  & ~_0996_;
	assign _0023_ = \mchip.run_chrono  & ~_0031_;
	assign _0997_ = \mchip.power_state  & ~\mchip.power_buf ;
	assign _0998_ = _0997_ | io_in[13];
	assign _0999_ = \mchip.leddrive0.power_mode [5] & ~_0998_;
	assign _1000_ = io_in[13] | ~_0997_;
	assign _1001_ = \mchip.leddrive0.power_mode [3] & ~_1000_;
	assign _0008_ = _1001_ | _0999_;
	assign _1002_ = ~_0915_;
	assign _1003_ = _0909_ | _0906_;
	assign _1004_ = \mchip.clock_digit_sel [0] & ~\mchip.clock_digit_sel [1];
	assign _1005_ = _1004_ | _0905_;
	assign _1006_ = _1005_ | _1003_;
	assign _1007_ = _0868_ & ~_1006_;
	assign _1008_ = _1007_ | _0912_;
	assign _0016_ = _1002_ & ~_1008_;
	assign _1009_ = ~\mchip.stop_buf ;
	assign _1010_ = \mchip.stophold0.button_latched  | io_in[13];
	assign _1011_ = _1010_ | _1009_;
	assign _1012_ = \mchip.stophold0.button_state [2] & ~_1011_;
	assign _1013_ = io_in[13] | ~\mchip.stop_buf ;
	assign _1014_ = \mchip.stophold0.button_state [0] & ~_1013_;
	assign _0014_ = _1014_ | _1012_;
	assign _1015_ = io_in[13] | ~\mchip.stophold0.button_latched ;
	assign _1016_ = \mchip.stophold0.button_state [2] & ~_1015_;
	assign _1017_ = \mchip.stophold0.button_state [1] & ~_1013_;
	assign _0013_ = _1017_ | _1016_;
	assign _1018_ = _1009_ & ~_1010_;
	assign _1019_ = ~(\mchip.stop_buf  | io_in[13]);
	assign _1020_ = ~(\mchip.stophold0.button_state [1] | \mchip.stophold0.button_state [0]);
	assign _1021_ = _1019_ & ~_1020_;
	assign _1022_ = _1021_ | io_in[13];
	assign _0012_ = _1022_ | _1018_;
	assign _1023_ = ~\mchip.mode_buf ;
	assign _1024_ = io_in[13] | \mchip.modehold0.button_latched ;
	assign _1025_ = _1024_ | _1023_;
	assign _1026_ = \mchip.modehold0.button_state [2] & ~_1025_;
	assign _1027_ = io_in[13] | ~\mchip.mode_buf ;
	assign _1028_ = \mchip.modehold0.button_state [0] & ~_1027_;
	assign _0011_ = _1028_ | _1026_;
	assign _1029_ = io_in[13] | ~\mchip.modehold0.button_latched ;
	assign _1030_ = \mchip.modehold0.button_state [2] & ~_1029_;
	assign _1031_ = \mchip.modehold0.button_state [1] & ~_1027_;
	assign _0010_ = _1031_ | _1030_;
	assign _1032_ = _1023_ & ~_1024_;
	assign _1033_ = ~(\mchip.mode_buf  | io_in[13]);
	assign _1034_ = ~(\mchip.modehold0.button_state [1] | \mchip.modehold0.button_state [0]);
	assign _1035_ = _1033_ & ~_1034_;
	assign _1036_ = _1035_ | io_in[13];
	assign _0009_ = _1036_ | _1032_;
	assign _1037_ = \mchip.cur_state [2] & ~_0833_;
	assign _1038_ = ~(\mchip.cur_state [2] | \mchip.cur_state [1]);
	assign _1039_ = _0835_ & ~_1038_;
	assign _1040_ = _1039_ | _1037_;
	assign _1041_ = \mchip.cur_state [0] & ~_0831_;
	assign _1042_ = _1041_ | io_in[13];
	assign _0000_ = _1042_ | _1040_;
	assign _1043_ = \mchip.leddrive0.power_mode [2] & ~_1000_;
	assign _1044_ = \mchip.leddrive0.power_mode [0] & ~_0998_;
	assign _1045_ = _1044_ | io_in[13];
	assign _0003_ = _1045_ | _1043_;
	assign _1046_ = \mchip.leddrive0.power_mode [4] & ~_0998_;
	assign _1047_ = \mchip.leddrive0.power_mode [1] & ~_1000_;
	assign _0007_ = _1047_ | _1046_;
	assign _1048_ = ~(\mchip.button_count [0] | \mchip.button_count [1]);
	assign _1049_ = \mchip.button_count [2] | \mchip.button_count [3];
	assign _1050_ = _1048_ & ~_1049_;
	assign _1051_ = \mchip.button_count [6] | \mchip.button_count [7];
	assign _1052_ = \mchip.button_count [4] | ~\mchip.button_count [5];
	assign _1053_ = _1052_ | _1051_;
	assign _1054_ = _1050_ & ~_1053_;
	assign _1055_ = \mchip.button_count [14] | ~\mchip.button_count [15];
	assign _1056_ = \mchip.button_count [12] | ~\mchip.button_count [13];
	assign _1057_ = _1056_ | _1055_;
	assign _1058_ = \mchip.button_count [10] | \mchip.button_count [11];
	assign _1059_ = \mchip.button_count [9] | ~\mchip.button_count [8];
	assign _1060_ = _1059_ | _1058_;
	assign _1061_ = _1060_ | _1057_;
	assign _1062_ = _1054_ & ~_1061_;
	assign _1063_ = \mchip.button_count [16] & \mchip.button_count [17];
	assign _1064_ = ~(_1063_ & \mchip.button_count [18]);
	assign _0094_ = _1062_ & ~_1064_;
	assign _0024_ = _0094_ | io_in[13];
	assign _1065_ = ~(\mchip.leddrive0.colcount0.Q [0] | \mchip.leddrive0.colcount0.Q [1]);
	assign _1066_ = \mchip.leddrive0.colcount0.Q [2] & \mchip.leddrive0.colcount0.Q [3];
	assign _1067_ = _1066_ & _1065_;
	assign _1068_ = ~(\mchip.leddrive0.colcount0.Q [6] & \mchip.leddrive0.colcount0.Q [7]);
	assign _1069_ = ~(\mchip.leddrive0.colcount0.Q [4] & \mchip.leddrive0.colcount0.Q [5]);
	assign _1070_ = _1069_ | _1068_;
	assign _1071_ = _1067_ & ~_1070_;
	assign _1072_ = \mchip.leddrive0.colcount0.Q [8] & \mchip.leddrive0.colcount0.Q [9];
	assign _1073_ = ~(_1072_ & \mchip.leddrive0.colcount0.Q [10]);
	assign _0095_ = _1071_ & ~_1073_;
	assign _1326_[0] = ~\mchip.leddrive0.col_sel [0];
	assign _1074_ = \mchip.leddrive0.power_mode [3] & ~_0998_;
	assign _1075_ = \mchip.leddrive0.power_mode [4] & ~_1000_;
	assign _0006_ = _1075_ | _1074_;
	assign _0088_ = \mchip.clock_digit_sel [1] & ~\mchip.clock_digit_sel [0];
	assign _1076_ = ~(_0088_ | _1004_);
	assign _1077_ = _0907_ | ~_1076_;
	assign _1078_ = _0910_ & ~_1077_;
	assign _1079_ = _1078_ | _0912_;
	assign _0015_ = _1002_ & ~_1079_;
	assign _1080_ = \mchip.leddrive0.power_mode [2] & ~_0998_;
	assign _1081_ = \mchip.leddrive0.power_mode [5] & ~_1000_;
	assign _0005_ = _1081_ | _1080_;
	assign _1082_ = \mchip.leddrive0.power_mode [1] & ~_0998_;
	assign _1083_ = \mchip.leddrive0.power_mode [0] & ~_1000_;
	assign _0004_ = _1083_ | _1082_;
	assign _1084_ = \mchip.cur_state [0] & ~_0833_;
	assign _1085_ = \mchip.cur_state [2] & ~_0831_;
	assign _0002_ = _1085_ | _1084_;
	assign _1086_ = ~(\mchip.leddrive0.out_clockcount [0] | \mchip.leddrive0.out_clockcount [1]);
	assign _1087_ = \mchip.leddrive0.out_clockcount [2] | \mchip.leddrive0.out_clockcount [3];
	assign _1088_ = _1086_ & ~_1087_;
	assign _1089_ = \mchip.leddrive0.out_clockcount [6] | ~\mchip.leddrive0.out_clockcount [7];
	assign _1090_ = \mchip.leddrive0.out_clockcount [4] | \mchip.leddrive0.out_clockcount [5];
	assign _1091_ = _1090_ | _1089_;
	assign _1092_ = _1088_ & ~_1091_;
	assign _1093_ = \mchip.leddrive0.out_clockcount [14] | ~\mchip.leddrive0.out_clockcount [15];
	assign _1094_ = \mchip.leddrive0.out_clockcount [13] | ~\mchip.leddrive0.out_clockcount [12];
	assign _1095_ = _1094_ | _1093_;
	assign _1096_ = \mchip.leddrive0.out_clockcount [11] | ~\mchip.leddrive0.out_clockcount [10];
	assign _1097_ = \mchip.leddrive0.out_clockcount [8] | ~\mchip.leddrive0.out_clockcount [9];
	assign _1098_ = _1097_ | _1096_;
	assign _1099_ = _1098_ | _1095_;
	assign _1100_ = _1092_ & ~_1099_;
	assign _1101_ = \mchip.leddrive0.out_clockcount [22] | ~\mchip.leddrive0.out_clockcount [23];
	assign _1102_ = \mchip.leddrive0.out_clockcount [21] | ~\mchip.leddrive0.out_clockcount [20];
	assign _1103_ = _1102_ | _1101_;
	assign _1104_ = \mchip.leddrive0.out_clockcount [18] | ~\mchip.leddrive0.out_clockcount [19];
	assign _1105_ = \mchip.leddrive0.out_clockcount [16] | \mchip.leddrive0.out_clockcount [17];
	assign _1106_ = _1105_ | _1104_;
	assign _1107_ = _1106_ | _1103_;
	assign _1108_ = _1100_ & ~_1107_;
	assign _0090_ = _1108_ | io_in[13];
	assign _1109_ = ~(\mchip.leddrive0.col_sel [3] & \mchip.leddrive0.col_sel [2]);
	assign _1110_ = ~(\mchip.leddrive0.col_sel [1] | \mchip.leddrive0.col_sel [0]);
	assign _1111_ = _1110_ & ~_1109_;
	assign _1112_ = _1111_ & _0095_;
	assign _0091_ = _1112_ | io_in[13];
	assign _1113_ = ~(\mchip.stophold0.button_state [2] & \mchip.stophold0.button_latched );
	assign _1114_ = \mchip.cur_state [1] & ~_1113_;
	assign _0033_ = _1114_ | io_in[13];
	assign _1115_ = ~(\mchip.leddrive0.col_sel [3] | \mchip.leddrive0.col_sel [2]);
	assign _1116_ = \mchip.leddrive0.col_sel [0] & ~\mchip.leddrive0.col_sel [1];
	assign _1117_ = _1116_ & _1115_;
	assign _1118_ = \mchip.leddrive0.col_sel [1] & ~\mchip.leddrive0.col_sel [0];
	assign _1119_ = _1118_ & _1115_;
	assign _1120_ = _1119_ | _1117_;
	assign _1121_ = \mchip.leddrive0.col_sel [1] & \mchip.leddrive0.col_sel [0];
	assign _1122_ = _1121_ & _1115_;
	assign _1123_ = \mchip.leddrive0.col_sel [3] | ~\mchip.leddrive0.col_sel [2];
	assign _1124_ = _1110_ & ~_1123_;
	assign _1125_ = _1124_ | _1122_;
	assign _1126_ = _1125_ | _1120_;
	assign _1127_ = _1115_ & _1110_;
	assign _1128_ = _1127_ | _1126_;
	assign _1129_ = _1116_ & ~_1123_;
	assign _1130_ = _1118_ & ~_1123_;
	assign _1131_ = _1130_ | _1129_;
	assign _1132_ = _1121_ & ~_1123_;
	assign _1133_ = \mchip.leddrive0.col_sel [2] | ~\mchip.leddrive0.col_sel [3];
	assign _1134_ = _1110_ & ~_1133_;
	assign _1135_ = _1134_ | _1132_;
	assign _1136_ = _1135_ | _1131_;
	assign _1137_ = _1116_ & ~_1133_;
	assign _1138_ = _1118_ & ~_1133_;
	assign _1139_ = _1138_ | _1137_;
	assign _1140_ = _1121_ & ~_1133_;
	assign _1141_ = _1140_ | _1111_;
	assign _1142_ = _1141_ | _1139_;
	assign _1143_ = _1142_ | _1136_;
	assign _1144_ = _1143_ | _1128_;
	assign _1145_ = (\mchip.cur_state [1] ? \mchip.chrono_time3 [3] : \mchip.clock_time3 [3]);
	assign _1146_ = ~_1145_;
	assign _1147_ = (\mchip.cur_state [1] ? \mchip.chrono_time3 [0] : \mchip.clock_time3 [0]);
	assign _1148_ = (\mchip.cur_state [1] ? \mchip.chrono_time3 [1] : \mchip.clock_time3 [1]);
	assign _1149_ = _1147_ | ~_1148_;
	assign _1150_ = _1148_ | ~_1147_;
	assign _1151_ = ~(_1150_ & _1149_);
	assign _1152_ = (\mchip.cur_state [1] ? \mchip.chrono_time3 [2] : \mchip.clock_time3 [2]);
	assign _1153_ = _1151_ | ~_1152_;
	assign _1154_ = _1153_ | ~_1146_;
	assign _1155_ = \mchip.leddrive0.out_clockcount [22] & \mchip.leddrive0.out_clockcount [21];
	assign _1156_ = ~\mchip.leddrive0.out_clockcount [20];
	assign _1157_ = \mchip.leddrive0.out_clockcount [20] & ~\mchip.leddrive0.out_clockcount [19];
	assign _1158_ = \mchip.leddrive0.out_clockcount [18] | \mchip.leddrive0.out_clockcount [17];
	assign _1159_ = _1157_ & ~_1158_;
	assign _1160_ = _1159_ | _1156_;
	assign _1161_ = \mchip.leddrive0.out_clockcount [18] | ~\mchip.leddrive0.out_clockcount [17];
	assign _1162_ = _1157_ & ~_1161_;
	assign _1163_ = ~(\mchip.leddrive0.out_clockcount [14] & \mchip.leddrive0.out_clockcount [13]);
	assign _1164_ = \mchip.leddrive0.out_clockcount [16] | \mchip.leddrive0.out_clockcount [15];
	assign _1165_ = _1164_ | ~_1163_;
	assign _1166_ = _1162_ & ~_1165_;
	assign _1167_ = _1166_ | _1160_;
	assign _1168_ = _1164_ | _1163_;
	assign _1169_ = _1162_ & ~_1168_;
	assign _1170_ = \mchip.leddrive0.out_clockcount [12] & ~\mchip.leddrive0.out_clockcount [11];
	assign _1171_ = \mchip.leddrive0.out_clockcount [10] | \mchip.leddrive0.out_clockcount [9];
	assign _1172_ = _1170_ & ~_1171_;
	assign _1173_ = \mchip.leddrive0.out_clockcount [8] | \mchip.leddrive0.out_clockcount [7];
	assign _1174_ = \mchip.leddrive0.out_clockcount [7] & ~\mchip.leddrive0.out_clockcount [8];
	assign _1175_ = \mchip.leddrive0.out_clockcount [6] & \mchip.leddrive0.out_clockcount [5];
	assign _1176_ = _1174_ & ~_1175_;
	assign _1177_ = _1173_ & ~_1176_;
	assign _1178_ = _1172_ & ~_1177_;
	assign _1179_ = \mchip.leddrive0.out_clockcount [12] & ~_1178_;
	assign _1180_ = _1169_ & ~_1179_;
	assign _1181_ = _1180_ | _1167_;
	assign _1182_ = _1181_ | ~_1155_;
	assign _1183_ = _1182_ & ~\mchip.leddrive0.out_clockcount [23];
	assign _1184_ = \mchip.leddrive0.out_clockcount [0] & \mchip.leddrive0.out_clockcount [1];
	assign _1185_ = ~(\mchip.leddrive0.out_clockcount [2] & \mchip.leddrive0.out_clockcount [3]);
	assign _1186_ = _1184_ & ~_1185_;
	assign _1187_ = ~(\mchip.leddrive0.out_clockcount [7] & \mchip.leddrive0.out_clockcount [6]);
	assign _1188_ = \mchip.leddrive0.out_clockcount [5] | ~\mchip.leddrive0.out_clockcount [4];
	assign _1189_ = _1188_ | _1187_;
	assign _1190_ = _1186_ & ~_1189_;
	assign _1191_ = \mchip.leddrive0.out_clockcount [15] | ~\mchip.leddrive0.out_clockcount [14];
	assign _1192_ = ~(\mchip.leddrive0.out_clockcount [12] & \mchip.leddrive0.out_clockcount [13]);
	assign _1193_ = _1192_ | _1191_;
	assign _1194_ = \mchip.leddrive0.out_clockcount [10] | \mchip.leddrive0.out_clockcount [11];
	assign _1195_ = \mchip.leddrive0.out_clockcount [9] | \mchip.leddrive0.out_clockcount [8];
	assign _1196_ = _1195_ | _1194_;
	assign _1197_ = _1196_ | _1193_;
	assign _1198_ = _1190_ & ~_1197_;
	assign _1199_ = ~(\mchip.leddrive0.out_clockcount [20] & \mchip.leddrive0.out_clockcount [21]);
	assign _1200_ = \mchip.leddrive0.out_clockcount [22] & ~\mchip.leddrive0.out_clockcount [23];
	assign _1201_ = _1199_ | ~_1200_;
	assign _1202_ = \mchip.leddrive0.out_clockcount [19] | \mchip.leddrive0.out_clockcount [18];
	assign _1203_ = \mchip.leddrive0.out_clockcount [16] | ~\mchip.leddrive0.out_clockcount [17];
	assign _1204_ = _1203_ | _1202_;
	assign _1205_ = _1204_ | _1201_;
	assign _1206_ = _1198_ & ~_1205_;
	assign _1207_ = _1183_ & ~_1206_;
	assign _1208_ = \mchip.leddrive0.out_clockcount [19] & \mchip.leddrive0.out_clockcount [18];
	assign _1209_ = \mchip.leddrive0.out_clockcount [20] | \mchip.leddrive0.out_clockcount [21];
	assign _1210_ = _1209_ | _1208_;
	assign _1211_ = _1208_ & ~_1209_;
	assign _1212_ = \mchip.leddrive0.out_clockcount [15] | \mchip.leddrive0.out_clockcount [14];
	assign _1213_ = _1212_ | _1105_;
	assign _1214_ = _1211_ & ~_1213_;
	assign _1215_ = _1210_ & ~_1214_;
	assign _1216_ = _1191_ | _1105_;
	assign _1217_ = _1211_ & ~_1216_;
	assign _1218_ = \mchip.leddrive0.out_clockcount [12] | \mchip.leddrive0.out_clockcount [13];
	assign _1219_ = _1218_ | \mchip.leddrive0.out_clockcount [11];
	assign _1220_ = \mchip.leddrive0.out_clockcount [10] | ~\mchip.leddrive0.out_clockcount [11];
	assign _1221_ = ~(_1220_ | _1218_);
	assign _1222_ = ~(\mchip.leddrive0.out_clockcount [9] & \mchip.leddrive0.out_clockcount [8]);
	assign _1223_ = \mchip.leddrive0.out_clockcount [7] | \mchip.leddrive0.out_clockcount [6];
	assign _1224_ = _1223_ & ~_1222_;
	assign _1225_ = _1221_ & ~_1224_;
	assign _1226_ = _1219_ & ~_1225_;
	assign _1227_ = _1217_ & ~_1226_;
	assign _1228_ = _1215_ & ~_1227_;
	assign _1229_ = _1200_ & ~_1228_;
	assign _1230_ = ~(\mchip.leddrive0.out_clockcount [23] | \mchip.leddrive0.out_clockcount [22]);
	assign _1231_ = _1230_ | _1229_;
	assign _1232_ = ~(\mchip.leddrive0.out_clockcount [4] & \mchip.leddrive0.out_clockcount [5]);
	assign _1233_ = _1232_ | _1223_;
	assign _1234_ = _1186_ & ~_1233_;
	assign _1235_ = _1218_ | _1191_;
	assign _1236_ = _1222_ | _1220_;
	assign _1237_ = _1236_ | _1235_;
	assign _1238_ = _1234_ & ~_1237_;
	assign _1239_ = _1209_ | ~_1200_;
	assign _1240_ = _1105_ | ~_1208_;
	assign _1241_ = _1240_ | _1239_;
	assign _1242_ = _1238_ & ~_1241_;
	assign _1243_ = _1231_ & ~_1242_;
	assign _1244_ = \mchip.leddrive0.out_clockcount [21] & ~\mchip.leddrive0.out_clockcount [20];
	assign _1245_ = ~(_1244_ & _1230_);
	assign _1246_ = \mchip.leddrive0.out_clockcount [19] | ~\mchip.leddrive0.out_clockcount [18];
	assign _1247_ = _1246_ | _1203_;
	assign _1248_ = _1247_ | _1245_;
	assign _1249_ = \mchip.leddrive0.out_clockcount [12] | ~\mchip.leddrive0.out_clockcount [13];
	assign _1250_ = _1249_ | _1212_;
	assign _1251_ = \mchip.leddrive0.out_clockcount [9] | ~\mchip.leddrive0.out_clockcount [8];
	assign _1252_ = _1251_ | _1096_;
	assign _1253_ = _1252_ | _1250_;
	assign _1254_ = ~(_1188_ | _1089_);
	assign _1255_ = ~(_1254_ & _1186_);
	assign _1256_ = _1255_ | _1253_;
	assign _1257_ = _1256_ | _1248_;
	assign _1258_ = \mchip.leddrive0.out_clockcount [22] | \mchip.leddrive0.out_clockcount [21];
	assign _1259_ = \mchip.leddrive0.out_clockcount [21] & ~\mchip.leddrive0.out_clockcount [22];
	assign _1260_ = \mchip.leddrive0.out_clockcount [18] & \mchip.leddrive0.out_clockcount [17];
	assign _1261_ = \mchip.leddrive0.out_clockcount [20] | \mchip.leddrive0.out_clockcount [19];
	assign _1262_ = _1261_ | _1260_;
	assign _1263_ = _1260_ & ~_1261_;
	assign _1264_ = \mchip.leddrive0.out_clockcount [14] | \mchip.leddrive0.out_clockcount [13];
	assign _1265_ = _1264_ | _1164_;
	assign _1266_ = _1263_ & ~_1265_;
	assign _1267_ = _1262_ & ~_1266_;
	assign _1268_ = \mchip.leddrive0.out_clockcount [14] | ~\mchip.leddrive0.out_clockcount [13];
	assign _1269_ = _1268_ | _1164_;
	assign _1270_ = _1263_ & ~_1269_;
	assign _1271_ = ~(\mchip.leddrive0.out_clockcount [12] | \mchip.leddrive0.out_clockcount [11]);
	assign _1272_ = \mchip.leddrive0.out_clockcount [10] | ~_1271_;
	assign _1273_ = \mchip.leddrive0.out_clockcount [9] | ~\mchip.leddrive0.out_clockcount [10];
	assign _1274_ = _1271_ & ~_1273_;
	assign _1275_ = \mchip.leddrive0.out_clockcount [8] & \mchip.leddrive0.out_clockcount [7];
	assign _1276_ = ~(\mchip.leddrive0.out_clockcount [6] | \mchip.leddrive0.out_clockcount [5]);
	assign _1277_ = _1275_ & ~_1276_;
	assign _1278_ = _1274_ & ~_1277_;
	assign _1279_ = _1272_ & ~_1278_;
	assign _1280_ = _1270_ & ~_1279_;
	assign _1281_ = _1267_ & ~_1280_;
	assign _1282_ = _1259_ & ~_1281_;
	assign _1283_ = _1258_ & ~_1282_;
	assign _1284_ = _1283_ | \mchip.leddrive0.out_clockcount [23];
	assign _1285_ = _1257_ & ~_1284_;
	assign _1286_ = _1243_ & ~_1285_;
	assign _1287_ = _1207_ & ~_1286_;
	assign _1288_ = _1287_ | _0905_;
	assign _1289_ = _1288_ | ~_0088_;
	assign _1290_ = \mchip.cur_state [2] | \mchip.cur_state [0];
	assign _1291_ = _1290_ | \mchip.cur_state [1];
	assign _1292_ = ~(\mchip.clock_time3 [2] | \mchip.clock_time3 [3]);
	assign _1293_ = \mchip.clock_time3 [0] | \mchip.clock_time3 [1];
	assign _1294_ = _1292_ & ~_1293_;
	assign _1295_ = _1290_ & ~_1294_;
	assign _1296_ = _1295_ | \mchip.cur_state [1];
	assign _1297_ = ~(_1296_ & _1291_);
	assign _1298_ = _1289_ & ~_1297_;
	assign _1299_ = _1298_ & _1154_;
	assign _1300_ = _1299_ | ~_1127_;
	assign _1301_ = _1117_ & ~_1299_;
	assign _1302_ = _1119_ & ~_1298_;
	assign _1303_ = _1302_ | _1301_;
	assign _1304_ = (\mchip.cur_state [1] ? \mchip.chrono_time2 [3] : \mchip.clock_time2 [3]);
	assign _1305_ = ~_1304_;
	assign _1306_ = (\mchip.cur_state [1] ? \mchip.chrono_time2 [0] : \mchip.clock_time2 [0]);
	assign _1307_ = (\mchip.cur_state [1] ? \mchip.chrono_time2 [1] : \mchip.clock_time2 [1]);
	assign _1308_ = _1306_ | ~_1307_;
	assign _1309_ = _1307_ | ~_1306_;
	assign _1310_ = ~(_1309_ & _1308_);
	assign _1311_ = (\mchip.cur_state [1] ? \mchip.chrono_time2 [2] : \mchip.clock_time2 [2]);
	assign _1312_ = _1310_ | ~_1311_;
	assign _1313_ = _1305_ & ~_1312_;
	assign _1314_ = _1289_ & ~_1313_;
	assign _1315_ = _1122_ & ~_1314_;
	assign _1316_ = _1124_ & ~_1314_;
	assign _1317_ = _1316_ | _1315_;
	assign _1318_ = _1317_ | _1303_;
	assign _1319_ = _1300_ & ~_1318_;
	assign _1320_ = _1129_ & ~_1289_;
	assign _0096_ = _1320_ | _1130_;
	assign _0097_ = (\mchip.cur_state [1] ? \mchip.chrono_time1 [3] : \mchip.clock_time1 [3]);
	assign _0098_ = ~_0097_;
	assign _0099_ = (\mchip.cur_state [1] ? \mchip.chrono_time1 [0] : \mchip.clock_time1 [0]);
	assign _0100_ = (\mchip.cur_state [1] ? \mchip.chrono_time1 [1] : \mchip.clock_time1 [1]);
	assign _0101_ = _0099_ | ~_0100_;
	assign _0102_ = _0100_ | ~_0099_;
	assign _0103_ = ~(_0102_ & _0101_);
	assign _0104_ = (\mchip.cur_state [1] ? \mchip.chrono_time1 [2] : \mchip.clock_time1 [2]);
	assign _0105_ = _0103_ | ~_0104_;
	assign _0106_ = _0105_ | ~_0098_;
	assign _0107_ = _1288_ | ~_1004_;
	assign _0108_ = _0107_ & _0106_;
	assign _0109_ = _1132_ & ~_0108_;
	assign _0110_ = _1134_ & ~_0108_;
	assign _0111_ = _0110_ | _0109_;
	assign _0112_ = _0111_ | _0096_;
	assign _0113_ = _1137_ & ~_0107_;
	assign _0114_ = (\mchip.cur_state [1] ? \mchip.chrono_time0 [3] : \mchip.clock_time0 [3]);
	assign _0115_ = ~_0114_;
	assign _0116_ = (\mchip.cur_state [1] ? \mchip.chrono_time0 [0] : \mchip.clock_time0 [0]);
	assign _0117_ = (\mchip.cur_state [1] ? \mchip.chrono_time0 [1] : \mchip.clock_time0 [1]);
	assign _0118_ = _0116_ | ~_0117_;
	assign _0119_ = _0117_ | ~_0116_;
	assign _0120_ = ~(_0119_ & _0118_);
	assign _0121_ = (\mchip.cur_state [1] ? \mchip.chrono_time0 [2] : \mchip.clock_time0 [2]);
	assign _0122_ = _0120_ | ~_0121_;
	assign _0123_ = _0122_ | ~_0115_;
	assign _0124_ = _1288_ | ~_0906_;
	assign _0125_ = _0124_ & _0123_;
	assign _0126_ = _1138_ & ~_0125_;
	assign _0127_ = _0126_ | _0113_;
	assign _0128_ = _1140_ & ~_0125_;
	assign _0129_ = _1111_ & ~_0124_;
	assign _0130_ = _0129_ | _0128_;
	assign _0131_ = _0130_ | _0127_;
	assign _0132_ = _0131_ | _0112_;
	assign _0133_ = _1319_ & ~_0132_;
	assign _0134_ = _1144_ & ~_0133_;
	assign _0135_ = \mchip.leddrive0.power_mode [4] | \mchip.leddrive0.power_mode [3];
	assign _0136_ = \mchip.leddrive0.power_mode [2] | \mchip.leddrive0.power_mode [5];
	assign _0137_ = _0136_ | _0135_;
	assign _0138_ = _0137_ | \mchip.leddrive0.power_mode [1];
	assign _0139_ = \mchip.leddrive0.colcount0.Q [8] | \mchip.leddrive0.colcount0.Q [9];
	assign _0140_ = \mchip.leddrive0.colcount0.Q [8] & ~\mchip.leddrive0.colcount0.Q [9];
	assign _0141_ = ~(\mchip.leddrive0.colcount0.Q [4] | \mchip.leddrive0.colcount0.Q [5]);
	assign _0142_ = \mchip.leddrive0.colcount0.Q [7] & ~\mchip.leddrive0.colcount0.Q [6];
	assign _0143_ = _0142_ & _0141_;
	assign _0144_ = \mchip.leddrive0.colcount0.Q [7] & ~_0143_;
	assign _0145_ = \mchip.leddrive0.colcount0.Q [5] | ~\mchip.leddrive0.colcount0.Q [4];
	assign _0146_ = _0142_ & ~_0145_;
	assign _0147_ = \mchip.leddrive0.colcount0.Q [2] | ~\mchip.leddrive0.colcount0.Q [3];
	assign _0148_ = _1065_ & ~_0147_;
	assign _0149_ = \mchip.leddrive0.colcount0.Q [3] & ~_0148_;
	assign _0150_ = _0146_ & ~_0149_;
	assign _0151_ = _0144_ & ~_0150_;
	assign _0152_ = _0140_ & ~_0151_;
	assign _0153_ = _0139_ & ~_0152_;
	assign _0154_ = _0153_ | \mchip.leddrive0.colcount0.Q [10];
	assign _0155_ = _0148_ & _0146_;
	assign _0156_ = ~\mchip.leddrive0.colcount0.Q [10];
	assign _0157_ = ~(_0140_ & _0156_);
	assign _0158_ = _0155_ & ~_0157_;
	assign _0159_ = _0158_ | _0154_;
	assign _0160_ = \mchip.leddrive0.power_mode [4] & ~_0159_;
	assign _0161_ = \mchip.leddrive0.colcount0.Q [2] | \mchip.leddrive0.colcount0.Q [3];
	assign _0162_ = _1065_ & ~_0161_;
	assign _0163_ = \mchip.leddrive0.colcount0.Q [6] | \mchip.leddrive0.colcount0.Q [7];
	assign _0164_ = _0163_ | _1069_;
	assign _0165_ = _0162_ & ~_0164_;
	assign _0166_ = ~(_1072_ & _0156_);
	assign _0167_ = _0165_ & ~_0166_;
	assign _0168_ = _1069_ & ~_0163_;
	assign _0169_ = _0168_ | _0165_;
	assign _0170_ = _1072_ & ~_0169_;
	assign _0171_ = _0170_ | \mchip.leddrive0.colcount0.Q [10];
	assign _0172_ = _0171_ | _0167_;
	assign _0173_ = \mchip.leddrive0.power_mode [3] & ~_0172_;
	assign _0174_ = _0173_ | _0160_;
	assign _0175_ = \mchip.leddrive0.colcount0.Q [7] & ~\mchip.leddrive0.colcount0.Q [8];
	assign _0176_ = \mchip.leddrive0.colcount0.Q [9] | ~\mchip.leddrive0.colcount0.Q [10];
	assign _0177_ = _0175_ & ~_0176_;
	assign _0178_ = ~(\mchip.leddrive0.colcount0.Q [6] & \mchip.leddrive0.colcount0.Q [5]);
	assign _0179_ = \mchip.leddrive0.colcount0.Q [6] & ~\mchip.leddrive0.colcount0.Q [5];
	assign _0180_ = ~(\mchip.leddrive0.colcount0.Q [4] | \mchip.leddrive0.colcount0.Q [3]);
	assign _0181_ = _0179_ & ~_0180_;
	assign _0182_ = _0178_ & ~_0181_;
	assign _0183_ = _0177_ & ~_0182_;
	assign _0184_ = \mchip.leddrive0.colcount0.Q [8] & ~_0176_;
	assign _0185_ = \mchip.leddrive0.colcount0.Q [10] & \mchip.leddrive0.colcount0.Q [9];
	assign _0186_ = _0185_ | _0184_;
	assign _0187_ = _0186_ | _0183_;
	assign _0188_ = _1068_ | ~_0141_;
	assign _0189_ = _0148_ & ~_0188_;
	assign _0190_ = _0139_ | _0156_;
	assign _0191_ = _0189_ & ~_0190_;
	assign _0192_ = _0191_ | _0187_;
	assign _0193_ = \mchip.leddrive0.power_mode [5] & ~_0192_;
	assign _0194_ = \mchip.leddrive0.colcount0.Q [8] | \mchip.leddrive0.colcount0.Q [7];
	assign _0195_ = _0178_ & ~_0194_;
	assign _0196_ = _0185_ & ~_0195_;
	assign _0197_ = \mchip.leddrive0.colcount0.Q [7] | ~\mchip.leddrive0.colcount0.Q [6];
	assign _0198_ = \mchip.leddrive0.colcount0.Q [4] | ~\mchip.leddrive0.colcount0.Q [5];
	assign _0199_ = _0198_ | _0197_;
	assign _0200_ = _0162_ & ~_0199_;
	assign _0201_ = \mchip.leddrive0.colcount0.Q [8] | ~\mchip.leddrive0.colcount0.Q [9];
	assign _0202_ = _0201_ | _0156_;
	assign _0203_ = _0200_ & ~_0202_;
	assign _0204_ = _0203_ | _0196_;
	assign _0205_ = \mchip.leddrive0.power_mode [2] & ~_0204_;
	assign _0206_ = _0205_ | _0193_;
	assign _0207_ = _0206_ | _0174_;
	assign _0208_ = _0138_ & ~_0207_;
	assign io_out[4] = _0208_ | _0134_;
	assign _0209_ = _0121_ | _0117_;
	assign _0210_ = ~(_0121_ | _0119_);
	assign _0211_ = (_0114_ ? _0209_ : _0210_);
	assign _0212_ = _0211_ & _0124_;
	assign _0213_ = _0212_ | ~_1140_;
	assign _0214_ = ~(_0117_ & _0116_);
	assign _0215_ = ~(_0117_ | _0116_);
	assign _0216_ = _0215_ | ~_0214_;
	assign _0217_ = _0216_ | _0121_;
	assign _0218_ = _0115_ & ~_0217_;
	assign _0219_ = _0124_ & ~_0218_;
	assign _0220_ = _1111_ & ~_0219_;
	assign _0221_ = _0213_ & ~_0220_;
	assign _0222_ = ~(_0100_ & _0099_);
	assign _0223_ = ~(_0100_ | _0099_);
	assign _0224_ = _0223_ | ~_0222_;
	assign _0225_ = _0224_ | _0104_;
	assign _0226_ = _0098_ & ~_0225_;
	assign _0227_ = _0107_ & ~_0226_;
	assign _0228_ = _1137_ & ~_0227_;
	assign _0229_ = (_0121_ ? _0118_ : _0116_);
	assign _0230_ = (_0114_ ? _0210_ : _0229_);
	assign _0231_ = _0124_ & ~_0230_;
	assign _0232_ = _1138_ & ~_0231_;
	assign _0233_ = _0232_ | _0228_;
	assign _0234_ = _0221_ & ~_0233_;
	assign _0235_ = ~(_1307_ & _1306_);
	assign _0236_ = ~(_1307_ | _1306_);
	assign _0237_ = _0236_ | ~_0235_;
	assign _0238_ = _0237_ | _1311_;
	assign _0239_ = _1305_ & ~_0238_;
	assign _0240_ = _1289_ & ~_0239_;
	assign _0241_ = _1129_ & ~_0240_;
	assign _0242_ = ~(_0104_ | _0102_);
	assign _0243_ = (_0104_ ? _0101_ : _0099_);
	assign _0244_ = (_0097_ ? _0242_ : _0243_);
	assign _0245_ = _0107_ & ~_0244_;
	assign _0246_ = _1132_ & ~_0245_;
	assign _0247_ = _0104_ | _0100_;
	assign _0248_ = (_0097_ ? _0247_ : _0242_);
	assign _0249_ = _0248_ & _0107_;
	assign _0250_ = _1134_ & ~_0249_;
	assign _0251_ = _0250_ | _0246_;
	assign _0252_ = _0251_ | _0241_;
	assign _0253_ = _0234_ & ~_0252_;
	assign _0254_ = ~(_1152_ | _1150_);
	assign _0255_ = (_1152_ ? _1149_ : _1147_);
	assign _0256_ = (_1145_ ? _0254_ : _0255_);
	assign _0257_ = _1298_ & ~_0256_;
	assign _0258_ = _1127_ & ~_0257_;
	assign _0259_ = _1152_ | _1148_;
	assign _0260_ = (_1145_ ? _0259_ : _0254_);
	assign _0261_ = _0260_ & _1298_;
	assign _0262_ = _1117_ & ~_0261_;
	assign _0263_ = ~(_1148_ & _1147_);
	assign _0264_ = ~(_1148_ | _1147_);
	assign _0265_ = _0264_ | ~_0263_;
	assign _0266_ = _0265_ | _1152_;
	assign _0267_ = _1146_ & ~_0266_;
	assign _0268_ = _1298_ & ~_0267_;
	assign _0269_ = _1119_ & ~_0268_;
	assign _0270_ = _0269_ | _0262_;
	assign _0271_ = ~(_1311_ | _1309_);
	assign _0272_ = (_1311_ ? _1308_ : _1306_);
	assign _0273_ = (_1304_ ? _0271_ : _0272_);
	assign _0274_ = _1289_ & ~_0273_;
	assign _0275_ = _1122_ & ~_0274_;
	assign _0276_ = _1311_ | _1307_;
	assign _0277_ = (_1304_ ? _0276_ : _0271_);
	assign _0278_ = _0277_ & _1289_;
	assign _0279_ = _1124_ & ~_0278_;
	assign _0280_ = _0279_ | _0275_;
	assign _0281_ = _0280_ | _0270_;
	assign _0282_ = _0281_ | _0258_;
	assign _0283_ = _0253_ & ~_0282_;
	assign _0284_ = _1144_ & ~_0283_;
	assign io_out[5] = _0284_ | _0208_;
	assign _0285_ = _0210_ & ~_0114_;
	assign _0286_ = _0124_ & ~_0285_;
	assign _0287_ = _0286_ | ~_1111_;
	assign _0288_ = ~_0215_;
	assign _0289_ = (_0121_ ? _0214_ : _0288_);
	assign _0290_ = _0115_ & ~_0289_;
	assign _0291_ = _0124_ & ~_0290_;
	assign _0292_ = _1140_ & ~_0291_;
	assign _0293_ = _0287_ & ~_0292_;
	assign _0294_ = _0242_ & ~_0097_;
	assign _0295_ = _0107_ & ~_0294_;
	assign _0296_ = _1137_ & ~_0295_;
	assign _0297_ = (_0121_ ? _0214_ : _0119_);
	assign _0298_ = _0115_ & ~_0297_;
	assign _0299_ = _0124_ & ~_0298_;
	assign _0300_ = _1138_ & ~_0299_;
	assign _0301_ = _0300_ | _0296_;
	assign _0302_ = _0293_ & ~_0301_;
	assign _0303_ = _0271_ & ~_1304_;
	assign _0304_ = _1289_ & ~_0303_;
	assign _0305_ = _1129_ & ~_0304_;
	assign _0306_ = \mchip.pm  & \mchip.cur_state [2];
	assign _0307_ = _1130_ & ~_0306_;
	assign _0308_ = _0307_ | _0305_;
	assign _0309_ = (_0104_ ? _0222_ : _0102_);
	assign _0310_ = _0098_ & ~_0309_;
	assign _0311_ = _0107_ & ~_0310_;
	assign _0312_ = _1132_ & ~_0311_;
	assign _0313_ = ~_0223_;
	assign _0314_ = (_0104_ ? _0222_ : _0313_);
	assign _0315_ = _0098_ & ~_0314_;
	assign _0316_ = _0107_ & ~_0315_;
	assign _0317_ = _1134_ & ~_0316_;
	assign _0318_ = _0317_ | _0312_;
	assign _0319_ = _0318_ | _0308_;
	assign _0320_ = _0302_ & ~_0319_;
	assign _0321_ = (_1152_ ? _0263_ : _1150_);
	assign _0322_ = _1146_ & ~_0321_;
	assign _0323_ = _1298_ & ~_0322_;
	assign _0324_ = _1127_ & ~_0323_;
	assign _0325_ = ~_0264_;
	assign _0326_ = (_1152_ ? _0263_ : _0325_);
	assign _0327_ = _1146_ & ~_0326_;
	assign _0328_ = _1298_ & ~_0327_;
	assign _0329_ = _1117_ & ~_0328_;
	assign _0330_ = _0254_ & ~_1145_;
	assign _0331_ = _1298_ & ~_0330_;
	assign _0332_ = _1119_ & ~_0331_;
	assign _0333_ = _0332_ | _0329_;
	assign _0334_ = (_1311_ ? _0235_ : _1309_);
	assign _0335_ = _1305_ & ~_0334_;
	assign _0336_ = _1289_ & ~_0335_;
	assign _0337_ = _1122_ & ~_0336_;
	assign _0338_ = ~_0236_;
	assign _0339_ = (_1311_ ? _0235_ : _0338_);
	assign _0340_ = _1305_ & ~_0339_;
	assign _0341_ = _1289_ & ~_0340_;
	assign _0342_ = _1124_ & ~_0341_;
	assign _0343_ = _0342_ | _0337_;
	assign _0344_ = _0343_ | _0333_;
	assign _0345_ = _0344_ | _0324_;
	assign _0346_ = _0320_ & ~_0345_;
	assign _0347_ = _1144_ & ~_0346_;
	assign io_out[6] = _0347_ | _0208_;
	assign _0348_ = (_0121_ ? _0216_ : _0119_);
	assign _0349_ = _0115_ & ~_0348_;
	assign _0350_ = _0124_ & ~_0349_;
	assign _0351_ = _1111_ & ~_0350_;
	assign _0352_ = _0213_ & ~_0351_;
	assign _0353_ = (_0104_ ? _0224_ : _0102_);
	assign _0354_ = _0098_ & ~_0353_;
	assign _0355_ = _0107_ & ~_0354_;
	assign _0356_ = _1137_ & ~_0355_;
	assign _0357_ = (_0121_ ? _0214_ : _0215_);
	assign _0358_ = _0115_ & ~_0357_;
	assign _0359_ = _0124_ & ~_0358_;
	assign _0360_ = _1138_ & ~_0359_;
	assign _0361_ = _0360_ | _0356_;
	assign _0362_ = _0352_ & ~_0361_;
	assign _0363_ = (_1311_ ? _0237_ : _1309_);
	assign _0364_ = _1305_ & ~_0363_;
	assign _0365_ = _1289_ & ~_0364_;
	assign _0366_ = _1129_ & ~_0365_;
	assign _0367_ = (_0104_ ? _0222_ : _0223_);
	assign _0368_ = _0098_ & ~_0367_;
	assign _0369_ = _0107_ & ~_0368_;
	assign _0370_ = _1132_ & ~_0369_;
	assign _0371_ = _0370_ | _0250_;
	assign _0372_ = _0371_ | _0366_;
	assign _0373_ = _0362_ & ~_0372_;
	assign _0374_ = (_1152_ ? _0263_ : _0264_);
	assign _0375_ = _1146_ & ~_0374_;
	assign _0376_ = _1298_ & ~_0375_;
	assign _0377_ = _1127_ & ~_0376_;
	assign _0378_ = (_1152_ ? _0265_ : _1150_);
	assign _0379_ = _1146_ & ~_0378_;
	assign _0380_ = _1298_ & ~_0379_;
	assign _0381_ = _1119_ & ~_0380_;
	assign _0382_ = _0381_ | _0262_;
	assign _0383_ = (_1311_ ? _0235_ : _0236_);
	assign _0384_ = _1305_ & ~_0383_;
	assign _0385_ = _1289_ & ~_0384_;
	assign _0386_ = _1122_ & ~_0385_;
	assign _0387_ = _0386_ | _0279_;
	assign _0388_ = _0387_ | _0382_;
	assign _0389_ = _0388_ | _0377_;
	assign _0390_ = _0373_ & ~_0389_;
	assign _0391_ = _1144_ & ~_0390_;
	assign io_out[7] = _0391_ | _0208_;
	assign _0392_ = ~(_0215_ & _0121_);
	assign _0393_ = _0115_ & ~_0392_;
	assign _0394_ = _0124_ & ~_0393_;
	assign _0395_ = _1140_ & ~_0394_;
	assign _0396_ = _0287_ & ~_0395_;
	assign _0397_ = _1138_ & ~_0124_;
	assign _0398_ = _0397_ | _0296_;
	assign _0399_ = _0396_ & ~_0398_;
	assign _0400_ = _0305_ | _1130_;
	assign _0401_ = _1132_ & ~_0107_;
	assign _0402_ = ~(_0223_ & _0104_);
	assign _0403_ = _0098_ & ~_0402_;
	assign _0404_ = _0107_ & ~_0403_;
	assign _0405_ = _1134_ & ~_0404_;
	assign _0406_ = _0405_ | _0401_;
	assign _0407_ = _0406_ | _0400_;
	assign _0408_ = _0399_ & ~_0407_;
	assign _0409_ = _1127_ & ~_1298_;
	assign _0410_ = ~(_0264_ & _1152_);
	assign _0411_ = _1146_ & ~_0410_;
	assign _0412_ = _1298_ & ~_0411_;
	assign _0413_ = _1117_ & ~_0412_;
	assign _0414_ = _0413_ | _0332_;
	assign _0415_ = _1122_ & ~_1289_;
	assign _0416_ = ~(_0236_ & _1311_);
	assign _0417_ = _1305_ & ~_0416_;
	assign _0418_ = _1289_ & ~_0417_;
	assign _0419_ = _1124_ & ~_0418_;
	assign _0420_ = _0419_ | _0415_;
	assign _0421_ = _0420_ | _0414_;
	assign _0422_ = _0421_ | _0409_;
	assign _0423_ = _0408_ & ~_0422_;
	assign _0424_ = _1144_ & ~_0423_;
	assign io_out[8] = _0424_ | _0208_;
	assign _0425_ = \mchip.clock_time3 [1] | ~\mchip.clock_time3 [0];
	assign _0426_ = _1292_ & ~_0425_;
	assign _0427_ = \mchip.clock_time2 [2] | \mchip.clock_time2 [3];
	assign _0428_ = \mchip.clock_time2 [1] | ~\mchip.clock_time2 [0];
	assign _0429_ = _0428_ | _0427_;
	assign _0430_ = _0426_ & ~_0429_;
	assign _0431_ = _0430_ ^ \mchip.pm ;
	assign _0432_ = \mchip.clock_time2 [0] | ~\mchip.clock_time2 [1];
	assign _0433_ = _0432_ | _0427_;
	assign _0434_ = _0426_ & ~_0433_;
	assign _0435_ = (_0434_ ? \mchip.pm  : _0431_);
	assign _0436_ = \mchip.clock_time2 [2] | ~\mchip.clock_time2 [3];
	assign _0437_ = ~(_0436_ | _0428_);
	assign _0438_ = (_0437_ ? \mchip.pm  : _0435_);
	assign _0439_ = \mchip.clock_time1 [2] & ~\mchip.clock_time1 [3];
	assign _0440_ = \mchip.clock_time1 [0] & ~\mchip.clock_time1 [1];
	assign _0441_ = _0440_ & _0439_;
	assign _0442_ = ~_0441_;
	assign _0443_ = (_0441_ ? _0438_ : \mchip.pm );
	assign _0444_ = \mchip.clock_time0 [3] & ~\mchip.clock_time0 [2];
	assign _0445_ = \mchip.clock_time0 [0] & ~\mchip.clock_time0 [1];
	assign _0446_ = _0445_ & _0444_;
	assign _0447_ = ~_0446_;
	assign _0448_ = (_0446_ ? _0443_ : \mchip.pm );
	assign _0449_ = _0443_ & _1004_;
	assign _0450_ = _0438_ & _0088_;
	assign _0451_ = _0450_ | _0449_;
	assign _0452_ = (_1076_ ? _0448_ : _0451_);
	assign _0034_ = (\mchip.cur_state [2] ? _0452_ : _0448_);
	assign _0089_ = ~(\mchip.clock_digit_sel [0] ^ \mchip.clock_digit_sel [1]);
	assign _0084_ = ~(_0446_ | \mchip.clock_time0 [0]);
	assign _0453_ = ~_0444_;
	assign _0454_ = \mchip.clock_time0 [1] & ~\mchip.clock_time0 [0];
	assign _0085_ = (_0445_ ? _0453_ : _0454_);
	assign _0455_ = \mchip.clock_time0 [1] & \mchip.clock_time0 [0];
	assign _0456_ = _0455_ ^ \mchip.clock_time0 [2];
	assign _0086_ = _0456_ & ~_0446_;
	assign _0457_ = ~(_0455_ & \mchip.clock_time0 [2]);
	assign _0458_ = _0457_ ^ \mchip.clock_time0 [3];
	assign _0087_ = _0447_ & ~_0458_;
	assign _0459_ = ~(_0441_ | \mchip.clock_time1 [0]);
	assign _0460_ = (_0446_ ? _0459_ : \mchip.clock_time1 [0]);
	assign _0461_ = (_1004_ ? _0459_ : _0460_);
	assign _0080_ = (\mchip.cur_state [2] ? _0461_ : _0460_);
	assign _0462_ = ~_0439_;
	assign _0463_ = \mchip.clock_time1 [1] & ~\mchip.clock_time1 [0];
	assign _0464_ = (_0440_ ? _0462_ : _0463_);
	assign _0465_ = (_0446_ ? _0464_ : \mchip.clock_time1 [1]);
	assign _0466_ = (_1004_ ? _0464_ : _0465_);
	assign _0081_ = (\mchip.cur_state [2] ? _0466_ : _0465_);
	assign _0467_ = \mchip.clock_time1 [1] & \mchip.clock_time1 [0];
	assign _0468_ = _0467_ ^ \mchip.clock_time1 [2];
	assign _0469_ = _0468_ & ~_0441_;
	assign _0470_ = (_0446_ ? _0469_ : \mchip.clock_time1 [2]);
	assign _0471_ = (_1004_ ? _0469_ : _0470_);
	assign _0082_ = (\mchip.cur_state [2] ? _0471_ : _0470_);
	assign _0472_ = ~(_0467_ & \mchip.clock_time1 [2]);
	assign _0473_ = _0472_ ^ \mchip.clock_time1 [3];
	assign _0474_ = _0442_ & ~_0473_;
	assign _0475_ = (_0446_ ? _0474_ : \mchip.clock_time1 [3]);
	assign _0476_ = (_1004_ ? _0474_ : _0475_);
	assign _0083_ = (\mchip.cur_state [2] ? _0476_ : _0475_);
	assign _0477_ = \mchip.clock_time2 [0] & ~_0434_;
	assign _0478_ = ~(_0477_ | _0437_);
	assign _0479_ = (_0441_ ? _0478_ : \mchip.clock_time2 [0]);
	assign _0480_ = (_0446_ ? _0479_ : \mchip.clock_time2 [0]);
	assign _0481_ = _0479_ & _1004_;
	assign _0482_ = _0478_ & _0088_;
	assign _0483_ = _0482_ | _0481_;
	assign _0484_ = (_1076_ ? _0480_ : _0483_);
	assign _0076_ = (\mchip.cur_state [2] ? _0484_ : _0480_);
	assign _0485_ = _0432_ & _0428_;
	assign _0486_ = _0485_ | _0434_;
	assign _0487_ = ~(_0486_ | _0437_);
	assign _0488_ = (_0441_ ? _0487_ : \mchip.clock_time2 [1]);
	assign _0489_ = (_0446_ ? _0488_ : \mchip.clock_time2 [1]);
	assign _0490_ = _0488_ & _1004_;
	assign _0491_ = _0487_ & _0088_;
	assign _0492_ = _0491_ | _0490_;
	assign _0493_ = (_1076_ ? _0489_ : _0492_);
	assign _0077_ = (\mchip.cur_state [2] ? _0493_ : _0489_);
	assign _0494_ = ~\mchip.clock_time2 [2];
	assign _0495_ = \mchip.clock_time2 [1] & \mchip.clock_time2 [0];
	assign _0496_ = _0495_ ^ _0494_;
	assign _0497_ = _0496_ | _0434_;
	assign _0498_ = ~(_0497_ | _0437_);
	assign _0499_ = (_0441_ ? _0498_ : \mchip.clock_time2 [2]);
	assign _0500_ = (_0446_ ? _0499_ : \mchip.clock_time2 [2]);
	assign _0501_ = _0499_ & _1004_;
	assign _0502_ = _0498_ & _0088_;
	assign _0503_ = _0502_ | _0501_;
	assign _0504_ = (_1076_ ? _0500_ : _0503_);
	assign _0078_ = (\mchip.cur_state [2] ? _0504_ : _0500_);
	assign _0505_ = ~(_0495_ & \mchip.clock_time2 [2]);
	assign _0506_ = _0505_ ^ \mchip.clock_time2 [3];
	assign _0507_ = _0506_ | _0434_;
	assign _0508_ = ~(_0507_ | _0437_);
	assign _0509_ = (_0441_ ? _0508_ : \mchip.clock_time2 [3]);
	assign _0510_ = (_0446_ ? _0509_ : \mchip.clock_time2 [3]);
	assign _0511_ = _0509_ & _1004_;
	assign _0512_ = _0508_ & _0088_;
	assign _0513_ = _0512_ | _0511_;
	assign _0514_ = (_1076_ ? _0510_ : _0513_);
	assign _0079_ = (\mchip.cur_state [2] ? _0514_ : _0510_);
	assign _0515_ = \mchip.clock_time3 [0] & ~_0434_;
	assign _0516_ = ~(_0515_ | _0437_);
	assign _0517_ = ~_0516_;
	assign _0518_ = (_0441_ ? _0517_ : \mchip.clock_time3 [0]);
	assign _0519_ = (_0446_ ? _0518_ : \mchip.clock_time3 [0]);
	assign _0520_ = _0518_ & _1004_;
	assign _0521_ = _0088_ & ~_0516_;
	assign _0522_ = _0521_ | _0520_;
	assign _0523_ = (_1076_ ? _0519_ : _0522_);
	assign _0072_ = (\mchip.cur_state [2] ? _0523_ : _0519_);
	assign _0524_ = _0434_ | ~\mchip.clock_time3 [1];
	assign _0525_ = ~(_0524_ | _0437_);
	assign _0526_ = (_0441_ ? _0525_ : \mchip.clock_time3 [1]);
	assign _0527_ = (_0446_ ? _0526_ : \mchip.clock_time3 [1]);
	assign _0528_ = _0526_ & _1004_;
	assign _0529_ = _0525_ & _0088_;
	assign _0530_ = _0529_ | _0528_;
	assign _0531_ = (_1076_ ? _0527_ : _0530_);
	assign _0073_ = (\mchip.cur_state [2] ? _0531_ : _0527_);
	assign _0532_ = _0434_ | ~\mchip.clock_time3 [2];
	assign _0533_ = ~(_0532_ | _0437_);
	assign _0534_ = (_0441_ ? _0533_ : \mchip.clock_time3 [2]);
	assign _0535_ = (_0446_ ? _0534_ : \mchip.clock_time3 [2]);
	assign _0536_ = _0534_ & _1004_;
	assign _0537_ = _0533_ & _0088_;
	assign _0538_ = _0537_ | _0536_;
	assign _0539_ = (_1076_ ? _0535_ : _0538_);
	assign _0074_ = (\mchip.cur_state [2] ? _0539_ : _0535_);
	assign _0540_ = _0434_ | ~\mchip.clock_time3 [3];
	assign _0541_ = ~(_0540_ | _0437_);
	assign _0542_ = (_0441_ ? _0541_ : \mchip.clock_time3 [3]);
	assign _0543_ = (_0446_ ? _0542_ : \mchip.clock_time3 [3]);
	assign _0544_ = _0542_ & _1004_;
	assign _0545_ = _0541_ & _0088_;
	assign _0546_ = _0545_ | _0544_;
	assign _0547_ = (_1076_ ? _0543_ : _0546_);
	assign _0075_ = (\mchip.cur_state [2] ? _0547_ : _0543_);
	assign _0047_ = ~(_0939_ & \mchip.chrono_count [0]);
	assign _0548_ = \mchip.chrono_count [0] & \mchip.chrono_count [1];
	assign _0549_ = _0548_ | ~_0935_;
	assign _0058_ = _0939_ & ~_0549_;
	assign _0550_ = ~(_0548_ ^ \mchip.chrono_count [2]);
	assign _0063_ = _0939_ & ~_0550_;
	assign _0551_ = ~(_0548_ & \mchip.chrono_count [2]);
	assign _0552_ = _0551_ ^ \mchip.chrono_count [3];
	assign _0064_ = _0939_ & ~_0552_;
	assign _0553_ = ~(\mchip.chrono_count [2] & \mchip.chrono_count [3]);
	assign _0554_ = _0548_ & ~_0553_;
	assign _0555_ = ~(_0554_ ^ \mchip.chrono_count [4]);
	assign _0065_ = _0939_ & ~_0555_;
	assign _0556_ = ~(_0554_ & \mchip.chrono_count [4]);
	assign _0557_ = _0556_ ^ \mchip.chrono_count [5];
	assign _0066_ = _0939_ & ~_0557_;
	assign _0558_ = ~(\mchip.chrono_count [4] & \mchip.chrono_count [5]);
	assign _0559_ = _0554_ & ~_0558_;
	assign _0560_ = ~(_0559_ ^ \mchip.chrono_count [6]);
	assign _0067_ = _0939_ & ~_0560_;
	assign _0561_ = ~(_0559_ & \mchip.chrono_count [6]);
	assign _0562_ = _0561_ ^ \mchip.chrono_count [7];
	assign _0068_ = _0939_ & ~_0562_;
	assign _0563_ = ~(\mchip.chrono_count [7] & \mchip.chrono_count [6]);
	assign _0564_ = _0563_ | _0558_;
	assign _0565_ = _0554_ & ~_0564_;
	assign _0566_ = ~(_0565_ ^ \mchip.chrono_count [8]);
	assign _0069_ = _0939_ & ~_0566_;
	assign _0567_ = ~(_0565_ & \mchip.chrono_count [8]);
	assign _0568_ = _0567_ ^ \mchip.chrono_count [9];
	assign _0070_ = _0939_ & ~_0568_;
	assign _0569_ = ~(\mchip.chrono_count [9] & \mchip.chrono_count [8]);
	assign _0570_ = _0565_ & ~_0569_;
	assign _0571_ = ~(_0570_ ^ \mchip.chrono_count [10]);
	assign _0048_ = _0939_ & ~_0571_;
	assign _0572_ = ~(_0570_ & \mchip.chrono_count [10]);
	assign _0573_ = _0572_ ^ \mchip.chrono_count [11];
	assign _0049_ = _0939_ & ~_0573_;
	assign _0574_ = ~(\mchip.chrono_count [10] & \mchip.chrono_count [11]);
	assign _0575_ = _0574_ | _0569_;
	assign _0576_ = _0565_ & ~_0575_;
	assign _0577_ = ~(_0576_ ^ \mchip.chrono_count [12]);
	assign _0050_ = _0939_ & ~_0577_;
	assign _0578_ = ~(_0576_ & \mchip.chrono_count [12]);
	assign _0579_ = _0578_ ^ \mchip.chrono_count [13];
	assign _0051_ = _0939_ & ~_0579_;
	assign _0580_ = ~(\mchip.chrono_count [12] & \mchip.chrono_count [13]);
	assign _0581_ = _0576_ & ~_0580_;
	assign _0582_ = ~(_0581_ ^ \mchip.chrono_count [14]);
	assign _0052_ = _0939_ & ~_0582_;
	assign _0583_ = ~(_0581_ & \mchip.chrono_count [14]);
	assign _0584_ = _0583_ ^ \mchip.chrono_count [15];
	assign _0053_ = _0939_ & ~_0584_;
	assign _0585_ = ~(\mchip.chrono_count [15] & \mchip.chrono_count [14]);
	assign _0586_ = _0585_ | _0580_;
	assign _0587_ = _0586_ | _0575_;
	assign _0588_ = _0565_ & ~_0587_;
	assign _0589_ = ~(_0588_ ^ \mchip.chrono_count [16]);
	assign _0054_ = _0939_ & ~_0589_;
	assign _0590_ = ~(_0588_ & \mchip.chrono_count [16]);
	assign _0591_ = _0590_ ^ \mchip.chrono_count [17];
	assign _0055_ = _0939_ & ~_0591_;
	assign _0592_ = ~(\mchip.chrono_count [16] & \mchip.chrono_count [17]);
	assign _0593_ = _0588_ & ~_0592_;
	assign _0594_ = ~(_0593_ ^ \mchip.chrono_count [18]);
	assign _0056_ = _0939_ & ~_0594_;
	assign _0595_ = ~(_0593_ & \mchip.chrono_count [18]);
	assign _0596_ = _0595_ ^ \mchip.chrono_count [19];
	assign _0057_ = _0939_ & ~_0596_;
	assign _0597_ = ~(\mchip.chrono_count [19] & \mchip.chrono_count [18]);
	assign _0598_ = _0597_ | _0592_;
	assign _0599_ = _0588_ & ~_0598_;
	assign _0600_ = ~(_0599_ ^ \mchip.chrono_count [20]);
	assign _0059_ = _0939_ & ~_0600_;
	assign _0601_ = ~(_0599_ & \mchip.chrono_count [20]);
	assign _0602_ = _0601_ ^ \mchip.chrono_count [21];
	assign _0060_ = _0939_ & ~_0602_;
	assign _0603_ = ~(\mchip.chrono_count [20] & \mchip.chrono_count [21]);
	assign _0604_ = _0599_ & ~_0603_;
	assign _0605_ = ~(_0604_ ^ \mchip.chrono_count [22]);
	assign _0061_ = _0939_ & ~_0605_;
	assign _0606_ = ~(_0604_ & \mchip.chrono_count [22]);
	assign _0607_ = _0606_ ^ \mchip.chrono_count [23];
	assign _0062_ = _0939_ & ~_0607_;
	assign _0043_ = ~(_0943_ | \mchip.chrono_time0 [0]);
	assign _0608_ = ~_0941_;
	assign _0609_ = \mchip.chrono_time0 [1] & ~\mchip.chrono_time0 [0];
	assign _0044_ = (_0942_ ? _0608_ : _0609_);
	assign _0610_ = \mchip.chrono_time0 [1] & \mchip.chrono_time0 [0];
	assign _0611_ = _0610_ ^ \mchip.chrono_time0 [2];
	assign _0045_ = _0611_ & ~_0943_;
	assign _0612_ = ~(_0610_ & \mchip.chrono_time0 [2]);
	assign _0613_ = _0612_ ^ \mchip.chrono_time0 [3];
	assign _0046_ = _0954_ & ~_0613_;
	assign _0039_ = ~(_0946_ | \mchip.chrono_time1 [0]);
	assign _0614_ = ~_0944_;
	assign _0615_ = \mchip.chrono_time1 [1] & ~\mchip.chrono_time1 [0];
	assign _0040_ = (_0945_ ? _0614_ : _0615_);
	assign _0616_ = \mchip.chrono_time1 [1] & \mchip.chrono_time1 [0];
	assign _0617_ = _0616_ ^ \mchip.chrono_time1 [2];
	assign _0041_ = _0617_ & ~_0946_;
	assign _0618_ = ~(_0616_ & \mchip.chrono_time1 [2]);
	assign _0619_ = _0618_ ^ \mchip.chrono_time1 [3];
	assign _0042_ = _0956_ & ~_0619_;
	assign _0027_ = ~(_0950_ | \mchip.chrono_time2 [0]);
	assign _0620_ = ~_0948_;
	assign _0621_ = \mchip.chrono_time2 [1] & ~\mchip.chrono_time2 [0];
	assign _0028_ = (_0949_ ? _0620_ : _0621_);
	assign _0622_ = \mchip.chrono_time2 [1] & \mchip.chrono_time2 [0];
	assign _0623_ = _0622_ ^ \mchip.chrono_time2 [2];
	assign _0029_ = _0623_ & ~_0950_;
	assign _0624_ = ~(_0622_ & \mchip.chrono_time2 [2]);
	assign _0625_ = _0624_ ^ \mchip.chrono_time2 [3];
	assign _0030_ = _0951_ & ~_0625_;
	assign _0626_ = \mchip.chrono_time3 [3] & ~\mchip.chrono_time3 [2];
	assign _0627_ = \mchip.chrono_time3 [1] | \mchip.chrono_time3 [0];
	assign _0628_ = _0626_ & ~_0627_;
	assign _0035_ = ~(_0628_ | \mchip.chrono_time3 [0]);
	assign _0036_ = \mchip.chrono_time3 [1] ^ \mchip.chrono_time3 [0];
	assign _0629_ = \mchip.chrono_time3 [1] & \mchip.chrono_time3 [0];
	assign _0630_ = _0629_ ^ \mchip.chrono_time3 [2];
	assign _0037_ = _0630_ & ~_0628_;
	assign _0631_ = _0629_ & \mchip.chrono_time3 [2];
	assign _0632_ = _0631_ ^ \mchip.chrono_time3 [3];
	assign _0038_ = _0632_ & ~_0628_;
	assign _1321_[0] = ~\mchip.button_count [0];
	assign _1324_[0] = ~\mchip.leddrive0.out_clockcount [0];
	assign \mchip.leddrive0.colcount0.D [0] = ~\mchip.leddrive0.colcount0.Q [0];
	assign \mchip.leddrive0.colcount0.reset  = _0095_ | io_in[13];
	assign _0633_ = \mchip.modehold0.button_state [2] | ~_1034_;
	assign _0634_ = _1034_ & ~_0828_;
	assign _0635_ = _0633_ & ~_0634_;
	assign _0092_ = _0635_ | io_in[13];
	assign _0636_ = \mchip.stophold0.button_state [2] | ~_1020_;
	assign _0637_ = _1020_ & _0909_;
	assign _0638_ = _0636_ & ~_0637_;
	assign _0093_ = _0638_ | io_in[13];
	assign _0071_ = _0866_ | ~\mchip.clock_count [0];
	assign \mchip.modehold0.buttoncount.reset  = \mchip.modehold0.button_state [0] | io_in[13];
	assign \mchip.stophold0.buttoncount.reset  = \mchip.stophold0.button_state [0] | io_in[13];
	assign _1327_[1] = _1118_ | _1116_;
	assign _1327_[2] = _1121_ ^ \mchip.leddrive0.col_sel [2];
	assign _0639_ = _1121_ & \mchip.leddrive0.col_sel [2];
	assign _1327_[3] = _0639_ ^ \mchip.leddrive0.col_sel [3];
	assign \mchip.modehold0.buttoncount.D [1] = \mchip.modehold0.buttoncount.Q [0] ^ \mchip.modehold0.buttoncount.Q [1];
	assign _0640_ = \mchip.modehold0.buttoncount.Q [0] & \mchip.modehold0.buttoncount.Q [1];
	assign \mchip.modehold0.buttoncount.D [2] = _0640_ ^ \mchip.modehold0.buttoncount.Q [2];
	assign _0641_ = _0640_ & \mchip.modehold0.buttoncount.Q [2];
	assign \mchip.modehold0.buttoncount.D [3] = _0641_ ^ \mchip.modehold0.buttoncount.Q [3];
	assign _0642_ = ~(\mchip.modehold0.buttoncount.Q [2] & \mchip.modehold0.buttoncount.Q [3]);
	assign _0643_ = _0640_ & ~_0642_;
	assign \mchip.modehold0.buttoncount.D [4] = _0643_ ^ \mchip.modehold0.buttoncount.Q [4];
	assign _0644_ = _0643_ & \mchip.modehold0.buttoncount.Q [4];
	assign \mchip.modehold0.buttoncount.D [5] = _0644_ ^ \mchip.modehold0.buttoncount.Q [5];
	assign _0645_ = ~(\mchip.modehold0.buttoncount.Q [4] & \mchip.modehold0.buttoncount.Q [5]);
	assign _0646_ = _0643_ & ~_0645_;
	assign \mchip.modehold0.buttoncount.D [6] = _0646_ ^ \mchip.modehold0.buttoncount.Q [6];
	assign _0647_ = _0646_ & \mchip.modehold0.buttoncount.Q [6];
	assign \mchip.modehold0.buttoncount.D [7] = _0647_ ^ \mchip.modehold0.buttoncount.Q [7];
	assign _0648_ = ~(\mchip.modehold0.buttoncount.Q [6] & \mchip.modehold0.buttoncount.Q [7]);
	assign _0649_ = _0648_ | _0645_;
	assign _0650_ = _0643_ & ~_0649_;
	assign \mchip.modehold0.buttoncount.D [8] = _0650_ ^ \mchip.modehold0.buttoncount.Q [8];
	assign _0651_ = _0650_ & \mchip.modehold0.buttoncount.Q [8];
	assign \mchip.modehold0.buttoncount.D [9] = _0651_ ^ \mchip.modehold0.buttoncount.Q [9];
	assign _0652_ = ~(\mchip.modehold0.buttoncount.Q [8] & \mchip.modehold0.buttoncount.Q [9]);
	assign _0653_ = _0650_ & ~_0652_;
	assign \mchip.modehold0.buttoncount.D [10] = _0653_ ^ \mchip.modehold0.buttoncount.Q [10];
	assign _0654_ = _0653_ & \mchip.modehold0.buttoncount.Q [10];
	assign \mchip.modehold0.buttoncount.D [11] = _0654_ ^ \mchip.modehold0.buttoncount.Q [11];
	assign _0655_ = _0652_ | _0885_;
	assign _0656_ = _0655_ | ~_0650_;
	assign \mchip.modehold0.buttoncount.D [12] = ~(_0656_ ^ \mchip.modehold0.buttoncount.Q [12]);
	assign _0657_ = \mchip.modehold0.buttoncount.Q [12] & ~_0656_;
	assign \mchip.modehold0.buttoncount.D [13] = _0657_ ^ \mchip.modehold0.buttoncount.Q [13];
	assign _0658_ = _0880_ & ~_0656_;
	assign \mchip.modehold0.buttoncount.D [14] = _0658_ ^ \mchip.modehold0.buttoncount.Q [14];
	assign _0659_ = _0658_ & \mchip.modehold0.buttoncount.Q [14];
	assign \mchip.modehold0.buttoncount.D [15] = _0659_ ^ \mchip.modehold0.buttoncount.Q [15];
	assign _0660_ = \mchip.modehold0.buttoncount.Q [14] & \mchip.modehold0.buttoncount.Q [15];
	assign _0661_ = ~(_0660_ & _0880_);
	assign _0662_ = _0661_ | _0655_;
	assign _0663_ = _0650_ & ~_0662_;
	assign \mchip.modehold0.buttoncount.D [16] = _0663_ ^ \mchip.modehold0.buttoncount.Q [16];
	assign _0664_ = _0663_ & \mchip.modehold0.buttoncount.Q [16];
	assign \mchip.modehold0.buttoncount.D [17] = _0664_ ^ \mchip.modehold0.buttoncount.Q [17];
	assign _0665_ = ~(\mchip.modehold0.buttoncount.Q [16] & \mchip.modehold0.buttoncount.Q [17]);
	assign _0666_ = _0663_ & ~_0665_;
	assign \mchip.modehold0.buttoncount.D [18] = _0666_ ^ \mchip.modehold0.buttoncount.Q [18];
	assign _0667_ = _0666_ & \mchip.modehold0.buttoncount.Q [18];
	assign \mchip.modehold0.buttoncount.D [19] = _0667_ ^ \mchip.modehold0.buttoncount.Q [19];
	assign _0668_ = ~(\mchip.modehold0.buttoncount.Q [18] & \mchip.modehold0.buttoncount.Q [19]);
	assign _0669_ = _0668_ | _0665_;
	assign _0670_ = _0669_ | ~_0663_;
	assign \mchip.modehold0.buttoncount.D [20] = ~(_0670_ ^ \mchip.modehold0.buttoncount.Q [20]);
	assign _0671_ = \mchip.modehold0.buttoncount.Q [20] & ~_0670_;
	assign \mchip.modehold0.buttoncount.D [21] = _0671_ ^ \mchip.modehold0.buttoncount.Q [21];
	assign _0672_ = ~(_0670_ | _0870_);
	assign \mchip.modehold0.buttoncount.D [22] = _0672_ ^ \mchip.modehold0.buttoncount.Q [22];
	assign _0673_ = _0672_ & \mchip.modehold0.buttoncount.Q [22];
	assign \mchip.modehold0.buttoncount.D [23] = _0673_ ^ \mchip.modehold0.buttoncount.Q [23];
	assign _0674_ = ~(\mchip.modehold0.buttoncount.Q [22] & \mchip.modehold0.buttoncount.Q [23]);
	assign _0675_ = _0674_ | _0870_;
	assign _0676_ = _0675_ | _0669_;
	assign _0677_ = _0663_ & ~_0676_;
	assign \mchip.modehold0.buttoncount.D [24] = _0677_ ^ \mchip.modehold0.buttoncount.Q [24];
	assign \mchip.stophold0.buttoncount.D [1] = \mchip.stophold0.buttoncount.Q [1] ^ \mchip.stophold0.buttoncount.Q [0];
	assign _0678_ = \mchip.stophold0.buttoncount.Q [1] & \mchip.stophold0.buttoncount.Q [0];
	assign \mchip.stophold0.buttoncount.D [2] = _0678_ ^ \mchip.stophold0.buttoncount.Q [2];
	assign _0679_ = _0678_ & \mchip.stophold0.buttoncount.Q [2];
	assign \mchip.stophold0.buttoncount.D [3] = _0679_ ^ \mchip.stophold0.buttoncount.Q [3];
	assign _0680_ = ~(\mchip.stophold0.buttoncount.Q [2] & \mchip.stophold0.buttoncount.Q [3]);
	assign _0681_ = _0678_ & ~_0680_;
	assign \mchip.stophold0.buttoncount.D [4] = _0681_ ^ \mchip.stophold0.buttoncount.Q [4];
	assign _0682_ = _0681_ & \mchip.stophold0.buttoncount.Q [4];
	assign \mchip.stophold0.buttoncount.D [5] = _0682_ ^ \mchip.stophold0.buttoncount.Q [5];
	assign _0683_ = ~(\mchip.stophold0.buttoncount.Q [4] & \mchip.stophold0.buttoncount.Q [5]);
	assign _0684_ = _0681_ & ~_0683_;
	assign \mchip.stophold0.buttoncount.D [6] = _0684_ ^ \mchip.stophold0.buttoncount.Q [6];
	assign _0685_ = _0684_ & \mchip.stophold0.buttoncount.Q [6];
	assign \mchip.stophold0.buttoncount.D [7] = _0685_ ^ \mchip.stophold0.buttoncount.Q [7];
	assign _0686_ = ~(\mchip.stophold0.buttoncount.Q [6] & \mchip.stophold0.buttoncount.Q [7]);
	assign _0687_ = _0686_ | _0683_;
	assign _0688_ = _0681_ & ~_0687_;
	assign \mchip.stophold0.buttoncount.D [8] = _0688_ ^ \mchip.stophold0.buttoncount.Q [8];
	assign _0689_ = _0688_ & \mchip.stophold0.buttoncount.Q [8];
	assign \mchip.stophold0.buttoncount.D [9] = _0689_ ^ \mchip.stophold0.buttoncount.Q [9];
	assign _0690_ = ~(\mchip.stophold0.buttoncount.Q [8] & \mchip.stophold0.buttoncount.Q [9]);
	assign _0691_ = _0688_ & ~_0690_;
	assign \mchip.stophold0.buttoncount.D [10] = _0691_ ^ \mchip.stophold0.buttoncount.Q [10];
	assign _0692_ = _0691_ & \mchip.stophold0.buttoncount.Q [10];
	assign \mchip.stophold0.buttoncount.D [11] = _0692_ ^ \mchip.stophold0.buttoncount.Q [11];
	assign _0693_ = _0690_ | _0975_;
	assign _0694_ = _0693_ | ~_0688_;
	assign \mchip.stophold0.buttoncount.D [12] = ~(_0694_ ^ \mchip.stophold0.buttoncount.Q [12]);
	assign _0695_ = \mchip.stophold0.buttoncount.Q [12] & ~_0694_;
	assign \mchip.stophold0.buttoncount.D [13] = _0695_ ^ \mchip.stophold0.buttoncount.Q [13];
	assign _0696_ = _0970_ & ~_0694_;
	assign \mchip.stophold0.buttoncount.D [14] = _0696_ ^ \mchip.stophold0.buttoncount.Q [14];
	assign _0697_ = _0696_ & \mchip.stophold0.buttoncount.Q [14];
	assign \mchip.stophold0.buttoncount.D [15] = _0697_ ^ \mchip.stophold0.buttoncount.Q [15];
	assign _0698_ = \mchip.stophold0.buttoncount.Q [14] & \mchip.stophold0.buttoncount.Q [15];
	assign _0699_ = ~(_0698_ & _0970_);
	assign _0700_ = _0699_ | _0693_;
	assign _0701_ = _0688_ & ~_0700_;
	assign \mchip.stophold0.buttoncount.D [16] = _0701_ ^ \mchip.stophold0.buttoncount.Q [16];
	assign _0702_ = _0701_ & \mchip.stophold0.buttoncount.Q [16];
	assign \mchip.stophold0.buttoncount.D [17] = _0702_ ^ \mchip.stophold0.buttoncount.Q [17];
	assign _0703_ = ~(\mchip.stophold0.buttoncount.Q [16] & \mchip.stophold0.buttoncount.Q [17]);
	assign _0704_ = _0701_ & ~_0703_;
	assign \mchip.stophold0.buttoncount.D [18] = _0704_ ^ \mchip.stophold0.buttoncount.Q [18];
	assign _0705_ = _0704_ & \mchip.stophold0.buttoncount.Q [18];
	assign \mchip.stophold0.buttoncount.D [19] = _0705_ ^ \mchip.stophold0.buttoncount.Q [19];
	assign _0706_ = ~(\mchip.stophold0.buttoncount.Q [18] & \mchip.stophold0.buttoncount.Q [19]);
	assign _0707_ = _0706_ | _0703_;
	assign _0708_ = _0707_ | ~_0701_;
	assign \mchip.stophold0.buttoncount.D [20] = ~(_0708_ ^ \mchip.stophold0.buttoncount.Q [20]);
	assign _0709_ = \mchip.stophold0.buttoncount.Q [20] & ~_0708_;
	assign \mchip.stophold0.buttoncount.D [21] = _0709_ ^ \mchip.stophold0.buttoncount.Q [21];
	assign _0710_ = ~(_0708_ | _0960_);
	assign \mchip.stophold0.buttoncount.D [22] = _0710_ ^ \mchip.stophold0.buttoncount.Q [22];
	assign _0711_ = _0710_ & \mchip.stophold0.buttoncount.Q [22];
	assign \mchip.stophold0.buttoncount.D [23] = _0711_ ^ \mchip.stophold0.buttoncount.Q [23];
	assign _0712_ = ~(\mchip.stophold0.buttoncount.Q [22] & \mchip.stophold0.buttoncount.Q [23]);
	assign _0713_ = _0712_ | _0960_;
	assign _0714_ = _0713_ | _0707_;
	assign _0715_ = _0701_ & ~_0714_;
	assign \mchip.stophold0.buttoncount.D [24] = _0715_ ^ \mchip.stophold0.buttoncount.Q [24];
	assign _1323_[1] = \mchip.clock_count [0] ^ \mchip.clock_count [1];
	assign _0716_ = \mchip.clock_count [0] & \mchip.clock_count [1];
	assign _1323_[2] = _0716_ ^ \mchip.clock_count [2];
	assign _0717_ = _0716_ & \mchip.clock_count [2];
	assign _1323_[3] = _0717_ ^ \mchip.clock_count [3];
	assign _0718_ = ~(\mchip.clock_count [2] & \mchip.clock_count [3]);
	assign _0719_ = _0716_ & ~_0718_;
	assign _1323_[4] = _0719_ ^ \mchip.clock_count [4];
	assign _0720_ = _0719_ & \mchip.clock_count [4];
	assign _1323_[5] = _0720_ ^ \mchip.clock_count [5];
	assign _0721_ = ~(\mchip.clock_count [4] & \mchip.clock_count [5]);
	assign _0722_ = _0719_ & ~_0721_;
	assign _1323_[6] = _0722_ ^ \mchip.clock_count [6];
	assign _0723_ = _0722_ & \mchip.clock_count [6];
	assign _1323_[7] = _0723_ ^ \mchip.clock_count [7];
	assign _0724_ = ~(\mchip.clock_count [6] & \mchip.clock_count [7]);
	assign _0725_ = _0724_ | _0721_;
	assign _0726_ = _0719_ & ~_0725_;
	assign _1323_[8] = _0726_ ^ \mchip.clock_count [8];
	assign _0727_ = _0726_ & \mchip.clock_count [8];
	assign _1323_[9] = _0727_ ^ \mchip.clock_count [9];
	assign _0728_ = ~(\mchip.clock_count [9] & \mchip.clock_count [8]);
	assign _0729_ = _0726_ & ~_0728_;
	assign _1323_[10] = _0729_ ^ \mchip.clock_count [10];
	assign _0730_ = _0729_ & \mchip.clock_count [10];
	assign _1323_[11] = _0730_ ^ \mchip.clock_count [11];
	assign _0731_ = ~(\mchip.clock_count [10] & \mchip.clock_count [11]);
	assign _0732_ = _0731_ | _0728_;
	assign _0733_ = _0726_ & ~_0732_;
	assign _1323_[12] = _0733_ ^ \mchip.clock_count [12];
	assign _0734_ = _0733_ & \mchip.clock_count [12];
	assign _1323_[13] = _0734_ ^ \mchip.clock_count [13];
	assign _0735_ = ~(\mchip.clock_count [12] & \mchip.clock_count [13]);
	assign _0736_ = _0733_ & ~_0735_;
	assign _1323_[14] = _0736_ ^ \mchip.clock_count [14];
	assign _0737_ = _0736_ & \mchip.clock_count [14];
	assign _1323_[15] = _0737_ ^ \mchip.clock_count [15];
	assign _0738_ = ~(\mchip.clock_count [14] & \mchip.clock_count [15]);
	assign _0739_ = _0738_ | _0735_;
	assign _0740_ = ~(_0739_ | _0732_);
	assign _0741_ = ~(_0740_ & _0726_);
	assign _1323_[16] = ~(_0741_ ^ \mchip.clock_count [16]);
	assign _0742_ = \mchip.clock_count [16] & ~_0741_;
	assign _1323_[17] = _0742_ ^ \mchip.clock_count [17];
	assign _0743_ = ~(_0741_ | _0862_);
	assign _1323_[18] = _0743_ ^ \mchip.clock_count [18];
	assign _0744_ = _0743_ & \mchip.clock_count [18];
	assign _1323_[19] = _0744_ ^ \mchip.clock_count [19];
	assign _0745_ = ~(\mchip.clock_count [18] & \mchip.clock_count [19]);
	assign _0746_ = _0745_ | _0862_;
	assign _0747_ = ~(_0746_ | _0741_);
	assign _1323_[20] = _0747_ ^ \mchip.clock_count [20];
	assign _0748_ = _0747_ & \mchip.clock_count [20];
	assign _1323_[21] = _0748_ ^ \mchip.clock_count [21];
	assign _0749_ = ~(\mchip.clock_count [20] & \mchip.clock_count [21]);
	assign _0750_ = _0747_ & ~_0749_;
	assign _1323_[22] = _0750_ ^ \mchip.clock_count [22];
	assign _0751_ = _0750_ & \mchip.clock_count [22];
	assign _1323_[23] = _0751_ ^ \mchip.clock_count [23];
	assign _0752_ = _0749_ | _0858_;
	assign _0753_ = _0752_ | _0746_;
	assign _0754_ = _0753_ | _0741_;
	assign _1323_[24] = ~(_0754_ ^ \mchip.clock_count [24]);
	assign _0755_ = \mchip.clock_count [24] & ~_0754_;
	assign _1323_[25] = _0755_ ^ \mchip.clock_count [25];
	assign _0756_ = ~(_0754_ | _0855_);
	assign _1323_[26] = _0756_ ^ \mchip.clock_count [26];
	assign _0757_ = _0756_ & \mchip.clock_count [26];
	assign _1323_[27] = _0757_ ^ \mchip.clock_count [27];
	assign _0758_ = ~(\mchip.clock_count [26] & \mchip.clock_count [27]);
	assign _0759_ = _0758_ | _0855_;
	assign _0760_ = ~(_0759_ | _0754_);
	assign _1323_[28] = _0760_ ^ \mchip.clock_count [28];
	assign _0761_ = _0760_ & \mchip.clock_count [28];
	assign _1323_[29] = _0761_ ^ \mchip.clock_count [29];
	assign _1322_[1] = \mchip.button_count [0] ^ \mchip.button_count [1];
	assign _0762_ = \mchip.button_count [0] & \mchip.button_count [1];
	assign _1322_[2] = _0762_ ^ \mchip.button_count [2];
	assign _0763_ = _0762_ & \mchip.button_count [2];
	assign _1322_[3] = _0763_ ^ \mchip.button_count [3];
	assign _0764_ = ~(\mchip.button_count [2] & \mchip.button_count [3]);
	assign _0765_ = _0762_ & ~_0764_;
	assign _1322_[4] = _0765_ ^ \mchip.button_count [4];
	assign _0766_ = _0765_ & \mchip.button_count [4];
	assign _1322_[5] = _0766_ ^ \mchip.button_count [5];
	assign _0767_ = ~(\mchip.button_count [5] & \mchip.button_count [4]);
	assign _0768_ = _0765_ & ~_0767_;
	assign _1322_[6] = _0768_ ^ \mchip.button_count [6];
	assign _0769_ = _0768_ & \mchip.button_count [6];
	assign _1322_[7] = _0769_ ^ \mchip.button_count [7];
	assign _0770_ = ~(\mchip.button_count [6] & \mchip.button_count [7]);
	assign _0771_ = _0770_ | _0767_;
	assign _0772_ = _0765_ & ~_0771_;
	assign _1322_[8] = _0772_ ^ \mchip.button_count [8];
	assign _0773_ = _0772_ & \mchip.button_count [8];
	assign _1322_[9] = _0773_ ^ \mchip.button_count [9];
	assign _0774_ = ~(\mchip.button_count [8] & \mchip.button_count [9]);
	assign _0775_ = _0772_ & ~_0774_;
	assign _1322_[10] = _0775_ ^ \mchip.button_count [10];
	assign _0776_ = _0775_ & \mchip.button_count [10];
	assign _1322_[11] = _0776_ ^ \mchip.button_count [11];
	assign _0777_ = ~(\mchip.button_count [10] & \mchip.button_count [11]);
	assign _0778_ = _0777_ | _0774_;
	assign _0779_ = _0772_ & ~_0778_;
	assign _1322_[12] = _0779_ ^ \mchip.button_count [12];
	assign _0780_ = _0779_ & \mchip.button_count [12];
	assign _1322_[13] = _0780_ ^ \mchip.button_count [13];
	assign _0781_ = ~(\mchip.button_count [13] & \mchip.button_count [12]);
	assign _0782_ = _0779_ & ~_0781_;
	assign _1322_[14] = _0782_ ^ \mchip.button_count [14];
	assign _0783_ = _0782_ & \mchip.button_count [14];
	assign _1322_[15] = _0783_ ^ \mchip.button_count [15];
	assign _0784_ = ~(\mchip.button_count [15] & \mchip.button_count [14]);
	assign _0785_ = _0784_ | _0781_;
	assign _0786_ = ~(_0785_ | _0778_);
	assign _0787_ = ~(_0786_ & _0772_);
	assign _1322_[16] = ~(_0787_ ^ \mchip.button_count [16]);
	assign _0788_ = \mchip.button_count [16] & ~_0787_;
	assign _1322_[17] = _0788_ ^ \mchip.button_count [17];
	assign _0789_ = _1063_ & ~_0787_;
	assign _1322_[18] = _0789_ ^ \mchip.button_count [18];
	assign _1325_[1] = \mchip.leddrive0.out_clockcount [0] ^ \mchip.leddrive0.out_clockcount [1];
	assign _1325_[2] = _1184_ ^ \mchip.leddrive0.out_clockcount [2];
	assign _0790_ = _1184_ & \mchip.leddrive0.out_clockcount [2];
	assign _1325_[3] = _0790_ ^ \mchip.leddrive0.out_clockcount [3];
	assign _1325_[4] = _1186_ ^ \mchip.leddrive0.out_clockcount [4];
	assign _0791_ = _1186_ & \mchip.leddrive0.out_clockcount [4];
	assign _1325_[5] = _0791_ ^ \mchip.leddrive0.out_clockcount [5];
	assign _0792_ = _1186_ & ~_1232_;
	assign _1325_[6] = _0792_ ^ \mchip.leddrive0.out_clockcount [6];
	assign _0793_ = _0792_ & \mchip.leddrive0.out_clockcount [6];
	assign _1325_[7] = _0793_ ^ \mchip.leddrive0.out_clockcount [7];
	assign _0794_ = _1232_ | _1187_;
	assign _0795_ = _0794_ | ~_1186_;
	assign _1325_[8] = ~(_0795_ ^ \mchip.leddrive0.out_clockcount [8]);
	assign _0796_ = \mchip.leddrive0.out_clockcount [8] & ~_0795_;
	assign _1325_[9] = _0796_ ^ \mchip.leddrive0.out_clockcount [9];
	assign _0797_ = ~(_0795_ | _1222_);
	assign _1325_[10] = _0797_ ^ \mchip.leddrive0.out_clockcount [10];
	assign _0798_ = _0797_ & \mchip.leddrive0.out_clockcount [10];
	assign _1325_[11] = _0798_ ^ \mchip.leddrive0.out_clockcount [11];
	assign _0799_ = ~(\mchip.leddrive0.out_clockcount [10] & \mchip.leddrive0.out_clockcount [11]);
	assign _0800_ = _0799_ | _1222_;
	assign _0801_ = _0800_ | _0795_;
	assign _1325_[12] = ~(_0801_ ^ \mchip.leddrive0.out_clockcount [12]);
	assign _0802_ = \mchip.leddrive0.out_clockcount [12] & ~_0801_;
	assign _1325_[13] = _0802_ ^ \mchip.leddrive0.out_clockcount [13];
	assign _0803_ = ~(_0801_ | _1192_);
	assign _1325_[14] = _0803_ ^ \mchip.leddrive0.out_clockcount [14];
	assign _0804_ = _0803_ & \mchip.leddrive0.out_clockcount [14];
	assign _1325_[15] = _0804_ ^ \mchip.leddrive0.out_clockcount [15];
	assign _0805_ = ~(\mchip.leddrive0.out_clockcount [15] & \mchip.leddrive0.out_clockcount [14]);
	assign _0806_ = _0805_ | _1192_;
	assign _0807_ = _0806_ | _0800_;
	assign _0808_ = ~(_0807_ | _0795_);
	assign _1325_[16] = _0808_ ^ \mchip.leddrive0.out_clockcount [16];
	assign _0809_ = _0808_ & \mchip.leddrive0.out_clockcount [16];
	assign _1325_[17] = _0809_ ^ \mchip.leddrive0.out_clockcount [17];
	assign _0810_ = ~(\mchip.leddrive0.out_clockcount [16] & \mchip.leddrive0.out_clockcount [17]);
	assign _0811_ = _0808_ & ~_0810_;
	assign _1325_[18] = _0811_ ^ \mchip.leddrive0.out_clockcount [18];
	assign _0812_ = _0811_ & \mchip.leddrive0.out_clockcount [18];
	assign _1325_[19] = _0812_ ^ \mchip.leddrive0.out_clockcount [19];
	assign _0813_ = _1208_ & ~_0810_;
	assign _0814_ = ~(_0813_ & _0808_);
	assign _1325_[20] = _0814_ ^ _1156_;
	assign _0815_ = \mchip.leddrive0.out_clockcount [20] & ~_0814_;
	assign _1325_[21] = _0815_ ^ \mchip.leddrive0.out_clockcount [21];
	assign _0816_ = ~(_0814_ | _1199_);
	assign _1325_[22] = _0816_ ^ \mchip.leddrive0.out_clockcount [22];
	assign _0817_ = _0816_ & \mchip.leddrive0.out_clockcount [22];
	assign _1325_[23] = _0817_ ^ \mchip.leddrive0.out_clockcount [23];
	assign \mchip.leddrive0.colcount0.D [1] = \mchip.leddrive0.colcount0.Q [0] ^ \mchip.leddrive0.colcount0.Q [1];
	assign _0818_ = \mchip.leddrive0.colcount0.Q [0] & \mchip.leddrive0.colcount0.Q [1];
	assign \mchip.leddrive0.colcount0.D [2] = _0818_ ^ \mchip.leddrive0.colcount0.Q [2];
	assign _0819_ = _0818_ & \mchip.leddrive0.colcount0.Q [2];
	assign \mchip.leddrive0.colcount0.D [3] = _0819_ ^ \mchip.leddrive0.colcount0.Q [3];
	assign _0820_ = _0818_ & _1066_;
	assign \mchip.leddrive0.colcount0.D [4] = _0820_ ^ \mchip.leddrive0.colcount0.Q [4];
	assign _0821_ = _0820_ & \mchip.leddrive0.colcount0.Q [4];
	assign \mchip.leddrive0.colcount0.D [5] = _0821_ ^ \mchip.leddrive0.colcount0.Q [5];
	assign _0822_ = _0820_ & ~_1069_;
	assign \mchip.leddrive0.colcount0.D [6] = _0822_ ^ \mchip.leddrive0.colcount0.Q [6];
	assign _0823_ = _0822_ & \mchip.leddrive0.colcount0.Q [6];
	assign \mchip.leddrive0.colcount0.D [7] = _0823_ ^ \mchip.leddrive0.colcount0.Q [7];
	assign _0824_ = _0820_ & ~_1070_;
	assign \mchip.leddrive0.colcount0.D [8] = _0824_ ^ \mchip.leddrive0.colcount0.Q [8];
	assign _0825_ = _0824_ & \mchip.leddrive0.colcount0.Q [8];
	assign \mchip.leddrive0.colcount0.D [9] = _0825_ ^ \mchip.leddrive0.colcount0.Q [9];
	assign _0826_ = _0824_ & _1072_;
	assign \mchip.leddrive0.colcount0.D [10] = _0826_ ^ \mchip.leddrive0.colcount0.Q [10];
	assign _0827_ = \mchip.mode_buf  | \mchip.modehold0.button_latched ;
	assign _0828_ = \mchip.modehold0.button_state [2] & ~_0827_;
	assign _0829_ = \mchip.modehold0.button_latched  & \mchip.modehold0.button_state [2];
	assign _0830_ = _0829_ | io_in[13];
	assign _0831_ = _0830_ | _0828_;
	assign _0832_ = \mchip.cur_state [1] & ~_0831_;
	assign _0833_ = io_in[13] | ~_0829_;
	assign _0834_ = \mchip.cur_state [1] & ~_0833_;
	assign _0835_ = _0828_ & ~_0830_;
	assign _0836_ = _0835_ & \mchip.cur_state [0];
	assign _0837_ = _0836_ | _0834_;
	assign _0001_ = _0837_ | _0832_;
	assign _0838_ = ~(\mchip.clock_count [0] | \mchip.clock_count [1]);
	assign _0839_ = \mchip.clock_count [2] | \mchip.clock_count [3];
	assign _0840_ = _0838_ & ~_0839_;
	assign _0841_ = \mchip.clock_count [6] | \mchip.clock_count [7];
	assign _0842_ = \mchip.clock_count [4] | \mchip.clock_count [5];
	assign _0843_ = _0842_ | _0841_;
	assign _0844_ = _0840_ & ~_0843_;
	assign _0845_ = \mchip.clock_count [15] | ~\mchip.clock_count [14];
	assign _0846_ = \mchip.clock_count [12] | \mchip.clock_count [13];
	assign _0847_ = _0846_ | _0845_;
	assign _0848_ = \mchip.clock_count [11] | ~\mchip.clock_count [10];
	assign _0849_ = \mchip.clock_count [8] | ~\mchip.clock_count [9];
	assign _0850_ = _0849_ | _0848_;
	assign _0851_ = _0850_ | _0847_;
	assign _0852_ = _0844_ & ~_0851_;
	assign _0853_ = \mchip.clock_count [28] | ~\mchip.clock_count [29];
	assign _0854_ = \mchip.clock_count [26] | \mchip.clock_count [27];
	assign _0855_ = ~(\mchip.clock_count [24] & \mchip.clock_count [25]);
	assign _0856_ = _0855_ | _0854_;
	assign _0857_ = _0856_ | _0853_;
	assign _0858_ = ~(\mchip.clock_count [22] & \mchip.clock_count [23]);
	assign _0859_ = \mchip.clock_count [20] | \mchip.clock_count [21];
	assign _0860_ = _0859_ | _0858_;
	assign _0861_ = \mchip.clock_count [18] | \mchip.clock_count [19];
	assign _0862_ = ~(\mchip.clock_count [16] & \mchip.clock_count [17]);
	assign _0863_ = _0862_ | _0861_;
	assign _0864_ = _0863_ | _0860_;
	assign _0865_ = _0864_ | _0857_;
	assign _0866_ = _0852_ & ~_0865_;
	assign _0867_ = _0866_ | io_in[13];
	assign _0026_ = _0867_ | \mchip.cur_state [2];
	assign _0868_ = \mchip.start_buf  | ~\mchip.start_state ;
	assign _0018_ = \mchip.cur_state [2] & ~_0868_;
	assign _0869_ = ~(\mchip.modehold0.buttoncount.Q [22] | \mchip.modehold0.buttoncount.Q [23]);
	assign _0870_ = ~(\mchip.modehold0.buttoncount.Q [20] & \mchip.modehold0.buttoncount.Q [21]);
	assign _0871_ = _0869_ & ~_0870_;
	assign _0872_ = \mchip.modehold0.buttoncount.Q [18] | \mchip.modehold0.buttoncount.Q [19];
	assign _0873_ = ~(_0872_ | \mchip.modehold0.buttoncount.Q [17]);
	assign _0874_ = _0871_ & ~_0873_;
	assign _0875_ = _0869_ & ~_0874_;
	assign _0876_ = \mchip.modehold0.buttoncount.Q [17] | ~\mchip.modehold0.buttoncount.Q [16];
	assign _0877_ = _0876_ | _0872_;
	assign _0878_ = _0871_ & ~_0877_;
	assign _0879_ = ~(\mchip.modehold0.buttoncount.Q [14] | \mchip.modehold0.buttoncount.Q [15]);
	assign _0880_ = \mchip.modehold0.buttoncount.Q [13] & \mchip.modehold0.buttoncount.Q [12];
	assign _0881_ = _0879_ & ~_0880_;
	assign _0882_ = \mchip.modehold0.buttoncount.Q [12] | ~\mchip.modehold0.buttoncount.Q [13];
	assign _0883_ = _0879_ & ~_0882_;
	assign _0884_ = ~(\mchip.modehold0.buttoncount.Q [8] | \mchip.modehold0.buttoncount.Q [9]);
	assign _0885_ = ~(\mchip.modehold0.buttoncount.Q [10] & \mchip.modehold0.buttoncount.Q [11]);
	assign _0886_ = _0885_ | _0884_;
	assign _0887_ = _0883_ & ~_0886_;
	assign _0888_ = _0881_ & ~_0887_;
	assign _0889_ = _0878_ & ~_0888_;
	assign _0890_ = _0875_ & ~_0889_;
	assign _0891_ = \mchip.modehold0.buttoncount.Q [24] & ~_0890_;
	assign _0892_ = ~(\mchip.modehold0.buttoncount.Q [0] | \mchip.modehold0.buttoncount.Q [1]);
	assign _0893_ = \mchip.modehold0.buttoncount.Q [2] | \mchip.modehold0.buttoncount.Q [3];
	assign _0894_ = _0892_ & ~_0893_;
	assign _0895_ = \mchip.modehold0.buttoncount.Q [6] | \mchip.modehold0.buttoncount.Q [7];
	assign _0896_ = \mchip.modehold0.buttoncount.Q [4] | \mchip.modehold0.buttoncount.Q [5];
	assign _0897_ = _0896_ | _0895_;
	assign _0898_ = _0894_ & ~_0897_;
	assign _0899_ = \mchip.modehold0.buttoncount.Q [9] | ~\mchip.modehold0.buttoncount.Q [8];
	assign _0900_ = ~(_0899_ | _0885_);
	assign _0901_ = ~(_0900_ & _0883_);
	assign _0902_ = _0898_ & ~_0901_;
	assign _0903_ = ~(_0878_ & \mchip.modehold0.buttoncount.Q [24]);
	assign _0904_ = _0902_ & ~_0903_;
	assign \mchip.modehold0.en_buttonlatch  = _0904_ | _0891_;
	assign \mchip.stophold0.buttoncount.D [0] = ~\mchip.stophold0.buttoncount.Q [0];
	assign _0905_ = ~\mchip.cur_state [2];
	assign _0906_ = ~(\mchip.clock_digit_sel [0] | \mchip.clock_digit_sel [1]);
	assign _0907_ = _0906_ | _0905_;
	assign _0908_ = ~(\mchip.stop_buf  | \mchip.stophold0.button_latched );
	assign _0909_ = ~(_0908_ & \mchip.stophold0.button_state [2]);
	assign _0910_ = _0868_ & ~_0909_;
	assign _0911_ = _0907_ | ~_0910_;
	assign _0912_ = _0905_ & ~_0866_;
	assign _0913_ = _0911_ & ~_0912_;
	assign _0914_ = _0909_ & ~_0905_;
	assign _0915_ = (_0868_ ? _0914_ : \mchip.cur_state [2]);
	assign _0017_ = _0913_ & ~_0915_;
	assign _0025_ = \mchip.cur_state [2] | io_in[13];
	assign _0032_ = ~\mchip.run_chrono ;
	assign _0916_ = (\mchip.run_chrono  ? _0909_ : _0868_);
	assign _0031_ = \mchip.cur_state [1] & ~_0916_;
	assign _0917_ = \mchip.chrono_count [22] | ~\mchip.chrono_count [23];
	assign _0918_ = \mchip.chrono_count [21] | ~\mchip.chrono_count [20];
	assign _0919_ = _0918_ | _0917_;
	assign _0920_ = \mchip.chrono_count [18] | ~\mchip.chrono_count [19];
	assign _0921_ = \mchip.chrono_count [16] | \mchip.chrono_count [17];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [1] <= 1'h0;
		else
			\mchip.clock_count [1] <= _1323_[1];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [2] <= 1'h0;
		else
			\mchip.clock_count [2] <= _1323_[2];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [3] <= 1'h0;
		else
			\mchip.clock_count [3] <= _1323_[3];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [4] <= 1'h0;
		else
			\mchip.clock_count [4] <= _1323_[4];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [5] <= 1'h0;
		else
			\mchip.clock_count [5] <= _1323_[5];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [6] <= 1'h0;
		else
			\mchip.clock_count [6] <= _1323_[6];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [7] <= 1'h0;
		else
			\mchip.clock_count [7] <= _1323_[7];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [8] <= 1'h0;
		else
			\mchip.clock_count [8] <= _1323_[8];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [9] <= 1'h0;
		else
			\mchip.clock_count [9] <= _1323_[9];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [10] <= 1'h0;
		else
			\mchip.clock_count [10] <= _1323_[10];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [11] <= 1'h0;
		else
			\mchip.clock_count [11] <= _1323_[11];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [12] <= 1'h0;
		else
			\mchip.clock_count [12] <= _1323_[12];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [13] <= 1'h0;
		else
			\mchip.clock_count [13] <= _1323_[13];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [14] <= 1'h0;
		else
			\mchip.clock_count [14] <= _1323_[14];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [15] <= 1'h0;
		else
			\mchip.clock_count [15] <= _1323_[15];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [16] <= 1'h0;
		else
			\mchip.clock_count [16] <= _1323_[16];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [17] <= 1'h0;
		else
			\mchip.clock_count [17] <= _1323_[17];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [18] <= 1'h0;
		else
			\mchip.clock_count [18] <= _1323_[18];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [19] <= 1'h0;
		else
			\mchip.clock_count [19] <= _1323_[19];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [20] <= 1'h0;
		else
			\mchip.clock_count [20] <= _1323_[20];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [21] <= 1'h0;
		else
			\mchip.clock_count [21] <= _1323_[21];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [22] <= 1'h0;
		else
			\mchip.clock_count [22] <= _1323_[22];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [23] <= 1'h0;
		else
			\mchip.clock_count [23] <= _1323_[23];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [24] <= 1'h0;
		else
			\mchip.clock_count [24] <= _1323_[24];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [25] <= 1'h0;
		else
			\mchip.clock_count [25] <= _1323_[25];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [26] <= 1'h0;
		else
			\mchip.clock_count [26] <= _1323_[26];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [27] <= 1'h0;
		else
			\mchip.clock_count [27] <= _1323_[27];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [28] <= 1'h0;
		else
			\mchip.clock_count [28] <= _1323_[28];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.clock_count [29] <= 1'h0;
		else
			\mchip.clock_count [29] <= _1323_[29];
	always @(posedge io_in[12]) \mchip.modehold0.button_state [0] <= _0009_;
	always @(posedge io_in[12]) \mchip.modehold0.button_state [1] <= _0010_;
	always @(posedge io_in[12]) \mchip.modehold0.button_state [2] <= _0011_;
	always @(posedge io_in[12]) \mchip.stophold0.button_state [0] <= _0012_;
	always @(posedge io_in[12]) \mchip.stophold0.button_state [1] <= _0013_;
	always @(posedge io_in[12]) \mchip.stophold0.button_state [2] <= _0014_;
	always @(posedge io_in[12]) \mchip.cur_state [0] <= _0000_;
	always @(posedge io_in[12]) \mchip.cur_state [1] <= _0001_;
	always @(posedge io_in[12]) \mchip.cur_state [2] <= _0002_;
	always @(posedge io_in[12])
		if (_0091_)
			\mchip.leddrive0.col_sel [0] <= 1'h0;
		else if (_0095_)
			\mchip.leddrive0.col_sel [0] <= _1326_[0];
	always @(posedge io_in[12])
		if (_0091_)
			\mchip.leddrive0.col_sel [1] <= 1'h0;
		else if (_0095_)
			\mchip.leddrive0.col_sel [1] <= _1327_[1];
	always @(posedge io_in[12])
		if (_0091_)
			\mchip.leddrive0.col_sel [2] <= 1'h0;
		else if (_0095_)
			\mchip.leddrive0.col_sel [2] <= _1327_[2];
	always @(posedge io_in[12])
		if (_0091_)
			\mchip.leddrive0.col_sel [3] <= 1'h0;
		else if (_0095_)
			\mchip.leddrive0.col_sel [3] <= _1327_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.power_bounce  <= 1'h0;
		else
			\mchip.power_bounce  <= \mchip.power_tmp1 ;
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [0] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [0] <= _1324_[0];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [1] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [1] <= _1325_[1];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [2] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [2] <= _1325_[2];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [3] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [3] <= _1325_[3];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [4] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [4] <= _1325_[4];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [5] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [5] <= _1325_[5];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [6] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [6] <= _1325_[6];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [7] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [7] <= _1325_[7];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [8] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [8] <= _1325_[8];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [9] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [9] <= _1325_[9];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [10] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [10] <= _1325_[10];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [11] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [11] <= _1325_[11];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [12] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [12] <= _1325_[12];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [13] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [13] <= _1325_[13];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [14] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [14] <= _1325_[14];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [15] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [15] <= _1325_[15];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [16] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [16] <= _1325_[16];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [17] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [17] <= _1325_[17];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [18] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [18] <= _1325_[18];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [19] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [19] <= _1325_[19];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [20] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [20] <= _1325_[20];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [21] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [21] <= _1325_[21];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [22] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [22] <= _1325_[22];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.leddrive0.out_clockcount [23] <= 1'h0;
		else
			\mchip.leddrive0.out_clockcount [23] <= _1325_[23];
	always @(posedge io_in[12])
		if (_0092_)
			\mchip.modehold0.button_latched  <= 1'h0;
		else if (\mchip.modehold0.en_buttonlatch )
			\mchip.modehold0.button_latched  <= 1'h1;
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [0] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [0] <= \mchip.modehold0.buttoncount.D [0];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [1] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [1] <= \mchip.modehold0.buttoncount.D [1];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [2] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [2] <= \mchip.modehold0.buttoncount.D [2];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [3] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [3] <= \mchip.modehold0.buttoncount.D [3];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [4] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [4] <= \mchip.modehold0.buttoncount.D [4];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [5] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [5] <= \mchip.modehold0.buttoncount.D [5];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [6] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [6] <= \mchip.modehold0.buttoncount.D [6];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [7] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [7] <= \mchip.modehold0.buttoncount.D [7];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [8] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [8] <= \mchip.modehold0.buttoncount.D [8];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [9] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [9] <= \mchip.modehold0.buttoncount.D [9];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [10] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [10] <= \mchip.modehold0.buttoncount.D [10];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [11] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [11] <= \mchip.modehold0.buttoncount.D [11];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [12] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [12] <= \mchip.modehold0.buttoncount.D [12];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [13] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [13] <= \mchip.modehold0.buttoncount.D [13];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [14] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [14] <= \mchip.modehold0.buttoncount.D [14];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [15] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [15] <= \mchip.modehold0.buttoncount.D [15];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [16] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [16] <= \mchip.modehold0.buttoncount.D [16];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [17] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [17] <= \mchip.modehold0.buttoncount.D [17];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [18] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [18] <= \mchip.modehold0.buttoncount.D [18];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [19] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [19] <= \mchip.modehold0.buttoncount.D [19];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [20] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [20] <= \mchip.modehold0.buttoncount.D [20];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [21] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [21] <= \mchip.modehold0.buttoncount.D [21];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [22] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [22] <= \mchip.modehold0.buttoncount.D [22];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [23] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [23] <= \mchip.modehold0.buttoncount.D [23];
	always @(posedge io_in[12])
		if (\mchip.modehold0.buttoncount.reset )
			\mchip.modehold0.buttoncount.Q [24] <= 1'h0;
		else if (\mchip.modehold0.button_state [2])
			\mchip.modehold0.buttoncount.Q [24] <= \mchip.modehold0.buttoncount.D [24];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [0] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [0] <= \mchip.leddrive0.colcount0.D [0];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [1] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [1] <= \mchip.leddrive0.colcount0.D [1];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [2] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [2] <= \mchip.leddrive0.colcount0.D [2];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [3] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [3] <= \mchip.leddrive0.colcount0.D [3];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [4] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [4] <= \mchip.leddrive0.colcount0.D [4];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [5] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [5] <= \mchip.leddrive0.colcount0.D [5];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [6] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [6] <= \mchip.leddrive0.colcount0.D [6];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [7] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [7] <= \mchip.leddrive0.colcount0.D [7];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [8] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [8] <= \mchip.leddrive0.colcount0.D [8];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [9] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [9] <= \mchip.leddrive0.colcount0.D [9];
	always @(posedge io_in[12])
		if (\mchip.leddrive0.colcount0.reset )
			\mchip.leddrive0.colcount0.Q [10] <= 1'h0;
		else
			\mchip.leddrive0.colcount0.Q [10] <= \mchip.leddrive0.colcount0.D [10];
	always @(posedge io_in[12])
		if (_0093_)
			\mchip.stophold0.button_latched  <= 1'h0;
		else if (\mchip.stophold0.en_buttonlatch )
			\mchip.stophold0.button_latched  <= 1'h1;
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [0] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [0] <= \mchip.stophold0.buttoncount.D [0];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [1] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [1] <= \mchip.stophold0.buttoncount.D [1];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [2] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [2] <= \mchip.stophold0.buttoncount.D [2];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [3] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [3] <= \mchip.stophold0.buttoncount.D [3];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [4] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [4] <= \mchip.stophold0.buttoncount.D [4];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [5] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [5] <= \mchip.stophold0.buttoncount.D [5];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [6] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [6] <= \mchip.stophold0.buttoncount.D [6];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [7] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [7] <= \mchip.stophold0.buttoncount.D [7];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [8] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [8] <= \mchip.stophold0.buttoncount.D [8];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [9] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [9] <= \mchip.stophold0.buttoncount.D [9];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [10] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [10] <= \mchip.stophold0.buttoncount.D [10];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [11] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [11] <= \mchip.stophold0.buttoncount.D [11];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [12] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [12] <= \mchip.stophold0.buttoncount.D [12];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [13] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [13] <= \mchip.stophold0.buttoncount.D [13];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [14] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [14] <= \mchip.stophold0.buttoncount.D [14];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [15] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [15] <= \mchip.stophold0.buttoncount.D [15];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [16] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [16] <= \mchip.stophold0.buttoncount.D [16];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [17] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [17] <= \mchip.stophold0.buttoncount.D [17];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [18] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [18] <= \mchip.stophold0.buttoncount.D [18];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [19] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [19] <= \mchip.stophold0.buttoncount.D [19];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [20] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [20] <= \mchip.stophold0.buttoncount.D [20];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [21] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [21] <= \mchip.stophold0.buttoncount.D [21];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [22] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [22] <= \mchip.stophold0.buttoncount.D [22];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [23] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [23] <= \mchip.stophold0.buttoncount.D [23];
	always @(posedge io_in[12])
		if (\mchip.stophold0.buttoncount.reset )
			\mchip.stophold0.buttoncount.Q [24] <= 1'h0;
		else if (\mchip.stophold0.button_state [2])
			\mchip.stophold0.buttoncount.Q [24] <= \mchip.stophold0.buttoncount.D [24];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.power_tmp0  <= 1'h0;
		else
			\mchip.power_tmp0  <= io_in[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.stop_tmp0  <= 1'h0;
		else
			\mchip.stop_tmp0  <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.start_tmp0  <= 1'h0;
		else
			\mchip.start_tmp0  <= io_in[3];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [0] <= 1'h0;
		else
			\mchip.button_count [0] <= _1321_[0];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [1] <= 1'h0;
		else
			\mchip.button_count [1] <= _1322_[1];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [2] <= 1'h0;
		else
			\mchip.button_count [2] <= _1322_[2];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [3] <= 1'h0;
		else
			\mchip.button_count [3] <= _1322_[3];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [4] <= 1'h0;
		else
			\mchip.button_count [4] <= _1322_[4];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [5] <= 1'h0;
		else
			\mchip.button_count [5] <= _1322_[5];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [6] <= 1'h0;
		else
			\mchip.button_count [6] <= _1322_[6];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [7] <= 1'h0;
		else
			\mchip.button_count [7] <= _1322_[7];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [8] <= 1'h0;
		else
			\mchip.button_count [8] <= _1322_[8];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [9] <= 1'h0;
		else
			\mchip.button_count [9] <= _1322_[9];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [10] <= 1'h0;
		else
			\mchip.button_count [10] <= _1322_[10];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [11] <= 1'h0;
		else
			\mchip.button_count [11] <= _1322_[11];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [12] <= 1'h0;
		else
			\mchip.button_count [12] <= _1322_[12];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [13] <= 1'h0;
		else
			\mchip.button_count [13] <= _1322_[13];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [14] <= 1'h0;
		else
			\mchip.button_count [14] <= _1322_[14];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [15] <= 1'h0;
		else
			\mchip.button_count [15] <= _1322_[15];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [16] <= 1'h0;
		else
			\mchip.button_count [16] <= _1322_[16];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [17] <= 1'h0;
		else
			\mchip.button_count [17] <= _1322_[17];
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.button_count [18] <= 1'h0;
		else
			\mchip.button_count [18] <= _1322_[18];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.power_buf  <= 1'h0;
		else if (_0094_)
			\mchip.power_buf  <= \mchip.power_bounce ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.mode_buf  <= 1'h0;
		else if (_0094_)
			\mchip.mode_buf  <= \mchip.mode_bounce ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.stop_buf  <= 1'h0;
		else if (_0094_)
			\mchip.stop_buf  <= \mchip.stop_bounce ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.start_buf  <= 1'h0;
		else if (_0094_)
			\mchip.start_buf  <= \mchip.start_bounce ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.power_state  <= 1'h0;
		else
			\mchip.power_state  <= \mchip.power_buf ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.start_state  <= 1'h0;
		else
			\mchip.start_state  <= \mchip.start_buf ;
	always @(posedge io_in[12])
		if (_0025_)
			\mchip.clock_count [0] <= 1'h0;
		else
			\mchip.clock_count [0] <= _0071_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time3 [0] <= 1'h1;
		else if (_0015_)
			\mchip.clock_time3 [0] <= _0072_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time3 [1] <= 1'h0;
		else if (_0015_)
			\mchip.clock_time3 [1] <= _0073_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time3 [2] <= 1'h0;
		else if (_0015_)
			\mchip.clock_time3 [2] <= _0074_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time3 [3] <= 1'h0;
		else if (_0015_)
			\mchip.clock_time3 [3] <= _0075_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time2 [0] <= 1'h0;
		else if (_0015_)
			\mchip.clock_time2 [0] <= _0076_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time2 [1] <= 1'h0;
		else if (_0015_)
			\mchip.clock_time2 [1] <= _0077_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time2 [2] <= 1'h0;
		else if (_0015_)
			\mchip.clock_time2 [2] <= _0078_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time2 [3] <= 1'h0;
		else if (_0015_)
			\mchip.clock_time2 [3] <= _0079_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time1 [0] <= 1'h1;
		else if (_0016_)
			\mchip.clock_time1 [0] <= _0080_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time1 [1] <= 1'h1;
		else if (_0016_)
			\mchip.clock_time1 [1] <= _0081_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time1 [2] <= 1'h0;
		else if (_0016_)
			\mchip.clock_time1 [2] <= _0082_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time1 [3] <= 1'h0;
		else if (_0016_)
			\mchip.clock_time1 [3] <= _0083_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time0 [0] <= 1'h0;
		else if (_0017_)
			\mchip.clock_time0 [0] <= _0084_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time0 [1] <= 1'h0;
		else if (_0017_)
			\mchip.clock_time0 [1] <= _0085_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time0 [2] <= 1'h1;
		else if (_0017_)
			\mchip.clock_time0 [2] <= _0086_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_time0 [3] <= 1'h0;
		else if (_0017_)
			\mchip.clock_time0 [3] <= _0087_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_digit_sel [0] <= 1'h0;
		else if (_0018_)
			\mchip.clock_digit_sel [0] <= _0088_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.clock_digit_sel [1] <= 1'h1;
		else if (_0018_)
			\mchip.clock_digit_sel [1] <= _0089_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.pm  <= 1'h0;
		else if (_0015_)
			\mchip.pm  <= _0034_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time3 [0] <= 1'h0;
		else if (_0019_)
			\mchip.chrono_time3 [0] <= _0035_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time3 [1] <= 1'h0;
		else if (_0019_)
			\mchip.chrono_time3 [1] <= _0036_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time3 [2] <= 1'h0;
		else if (_0019_)
			\mchip.chrono_time3 [2] <= _0037_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time3 [3] <= 1'h0;
		else if (_0019_)
			\mchip.chrono_time3 [3] <= _0038_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time2 [0] <= 1'h0;
		else if (_0020_)
			\mchip.chrono_time2 [0] <= _0027_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time2 [1] <= 1'h0;
		else if (_0020_)
			\mchip.chrono_time2 [1] <= _0028_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time2 [2] <= 1'h0;
		else if (_0020_)
			\mchip.chrono_time2 [2] <= _0029_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time2 [3] <= 1'h0;
		else if (_0020_)
			\mchip.chrono_time2 [3] <= _0030_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time1 [0] <= 1'h0;
		else if (_0021_)
			\mchip.chrono_time1 [0] <= _0039_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time1 [1] <= 1'h0;
		else if (_0021_)
			\mchip.chrono_time1 [1] <= _0040_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time1 [2] <= 1'h0;
		else if (_0021_)
			\mchip.chrono_time1 [2] <= _0041_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time1 [3] <= 1'h0;
		else if (_0021_)
			\mchip.chrono_time1 [3] <= _0042_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time0 [0] <= 1'h0;
		else if (_0022_)
			\mchip.chrono_time0 [0] <= _0043_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time0 [1] <= 1'h0;
		else if (_0022_)
			\mchip.chrono_time0 [1] <= _0044_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time0 [2] <= 1'h0;
		else if (_0022_)
			\mchip.chrono_time0 [2] <= _0045_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_time0 [3] <= 1'h0;
		else if (_0022_)
			\mchip.chrono_time0 [3] <= _0046_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [0] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [0] <= _0047_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [1] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [1] <= _0058_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [2] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [2] <= _0063_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [3] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [3] <= _0064_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [4] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [4] <= _0065_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [5] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [5] <= _0066_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [6] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [6] <= _0067_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [7] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [7] <= _0068_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [8] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [8] <= _0069_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [9] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [9] <= _0070_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [10] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [10] <= _0048_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [11] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [11] <= _0049_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [12] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [12] <= _0050_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [13] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [13] <= _0051_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [14] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [14] <= _0052_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [15] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [15] <= _0053_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [16] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [16] <= _0054_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [17] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [17] <= _0055_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [18] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [18] <= _0056_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [19] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [19] <= _0057_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [20] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [20] <= _0059_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [21] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [21] <= _0060_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [22] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [22] <= _0061_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.chrono_count [23] <= 1'h0;
		else if (_0023_)
			\mchip.chrono_count [23] <= _0062_;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.run_chrono  <= 1'h0;
		else if (_0031_)
			\mchip.run_chrono  <= _0032_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.stop_bounce  <= 1'h0;
		else
			\mchip.stop_bounce  <= \mchip.stop_tmp1 ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.mode_tmp0  <= 1'h0;
		else
			\mchip.mode_tmp0  <= io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.start_tmp1  <= 1'h0;
		else
			\mchip.start_tmp1  <= \mchip.start_tmp0 ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.mode_bounce  <= 1'h0;
		else
			\mchip.mode_bounce  <= \mchip.mode_tmp1 ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.stop_tmp1  <= 1'h0;
		else
			\mchip.stop_tmp1  <= \mchip.stop_tmp0 ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.power_tmp1  <= 1'h0;
		else
			\mchip.power_tmp1  <= \mchip.power_tmp0 ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.mode_tmp1  <= 1'h0;
		else
			\mchip.mode_tmp1  <= \mchip.mode_tmp0 ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.start_bounce  <= 1'h0;
		else
			\mchip.start_bounce  <= \mchip.start_tmp1 ;
	always @(posedge io_in[12]) \mchip.leddrive0.power_mode [0] <= _0003_;
	always @(posedge io_in[12]) \mchip.leddrive0.power_mode [1] <= _0004_;
	always @(posedge io_in[12]) \mchip.leddrive0.power_mode [2] <= _0005_;
	always @(posedge io_in[12]) \mchip.leddrive0.power_mode [3] <= _0006_;
	always @(posedge io_in[12]) \mchip.leddrive0.power_mode [4] <= _0007_;
	always @(posedge io_in[12]) \mchip.leddrive0.power_mode [5] <= _0008_;
	assign _1321_[18:1] = \mchip.button_count [18:1];
	assign _1322_[0] = _1321_[0];
	assign _1323_[0] = 1'h0;
	assign _1324_[23:1] = \mchip.leddrive0.out_clockcount [23:1];
	assign _1325_[0] = _1324_[0];
	assign _1326_[3:1] = \mchip.leddrive0.col_sel [3:1];
	assign _1327_[0] = _1326_[0];
	assign {io_out[13:9], io_out[3:0]} = {5'h00, \mchip.leddrive0.col_sel };
	assign \mchip.blink_drive  = \mchip.cur_state [2];
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {3'h0, io_out[8:4], \mchip.leddrive0.col_sel };
	assign \mchip.leddrive0.blink  = \mchip.cur_state [2];
	assign \mchip.leddrive0.blink_sel  = \mchip.clock_digit_sel ;
	assign \mchip.leddrive0.cd0.col0  = 5'h10;
	assign \mchip.leddrive0.cd0.col1  = 5'h00;
	assign \mchip.leddrive0.cd0.col2  = 5'h01;
	assign \mchip.leddrive0.cd1.col0  = 5'h10;
	assign \mchip.leddrive0.cd1.col1  = 5'h00;
	assign \mchip.leddrive0.cd1.col2  = 5'h01;
	assign \mchip.leddrive0.cd2.col0  = 5'h10;
	assign \mchip.leddrive0.cd2.col1  = 5'h00;
	assign \mchip.leddrive0.cd2.col2  = 5'h01;
	assign \mchip.leddrive0.cd3.col0  = 5'h10;
	assign \mchip.leddrive0.cd3.col1  = 5'h00;
	assign \mchip.leddrive0.cd3.col2  = 5'h01;
	assign \mchip.leddrive0.clock  = io_in[12];
	assign \mchip.leddrive0.colcount0.clock  = io_in[12];
	assign \mchip.leddrive0.colcount0.en  = 1'h1;
	assign \mchip.leddrive0.dig0col0  = 5'h10;
	assign \mchip.leddrive0.dig0col1  = 5'h00;
	assign \mchip.leddrive0.dig0col2  = 5'h01;
	assign \mchip.leddrive0.dig1col0  = 5'h10;
	assign \mchip.leddrive0.dig1col1  = 5'h00;
	assign \mchip.leddrive0.dig1col2  = 5'h01;
	assign \mchip.leddrive0.dig2col0  = 5'h10;
	assign \mchip.leddrive0.dig2col1  = 5'h00;
	assign \mchip.leddrive0.dig2col2  = 5'h01;
	assign \mchip.leddrive0.dig3col0  = 5'h10;
	assign \mchip.leddrive0.dig3col1  = 5'h00;
	assign \mchip.leddrive0.dig3col2  = 5'h01;
	assign \mchip.leddrive0.in_colcount  = \mchip.leddrive0.colcount0.D ;
	assign \mchip.leddrive0.out_colcount  = \mchip.leddrive0.colcount0.Q ;
	assign \mchip.leddrive0.reset  = io_in[13];
	assign \mchip.leddrive0.reset_colcount  = \mchip.leddrive0.colcount0.reset ;
	assign \mchip.leddrive0.row_L  = io_out[8:4];
	assign \mchip.modehold0.button  = \mchip.mode_buf ;
	assign \mchip.modehold0.buttoncount.clock  = io_in[12];
	assign \mchip.modehold0.buttoncount.en  = \mchip.modehold0.button_state [2];
	assign \mchip.modehold0.clear_buttoncount  = \mchip.modehold0.button_state [0];
	assign \mchip.modehold0.clock  = io_in[12];
	assign \mchip.modehold0.en_buttoncount  = \mchip.modehold0.button_state [2];
	assign \mchip.modehold0.in_buttoncount  = \mchip.modehold0.buttoncount.D ;
	assign \mchip.modehold0.out_buttoncount  = \mchip.modehold0.buttoncount.Q ;
	assign \mchip.modehold0.reset  = io_in[13];
	assign \mchip.modehold0.reset_buttoncount  = \mchip.modehold0.buttoncount.reset ;
	assign \mchip.power_state_next  = \mchip.power_buf ;
	assign \mchip.reset  = io_in[13];
	assign \mchip.start_state_next  = \mchip.start_buf ;
	assign \mchip.stophold0.button  = \mchip.stop_buf ;
	assign \mchip.stophold0.buttoncount.clock  = io_in[12];
	assign \mchip.stophold0.buttoncount.en  = \mchip.stophold0.button_state [2];
	assign \mchip.stophold0.clear_buttoncount  = \mchip.stophold0.button_state [0];
	assign \mchip.stophold0.clock  = io_in[12];
	assign \mchip.stophold0.en_buttoncount  = \mchip.stophold0.button_state [2];
	assign \mchip.stophold0.in_buttoncount  = \mchip.stophold0.buttoncount.D ;
	assign \mchip.stophold0.out_buttoncount  = \mchip.stophold0.buttoncount.Q ;
	assign \mchip.stophold0.reset  = io_in[13];
	assign \mchip.stophold0.reset_buttoncount  = \mchip.stophold0.buttoncount.reset ;
endmodule
module d18_vrajesh_motorcontroller (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	reg _0060_;
	reg _0061_;
	reg _0062_;
	reg _0063_;
	reg _0064_;
	reg _0065_;
	reg _0066_;
	reg _0067_;
	reg _0068_;
	reg _0069_;
	reg _0070_;
	reg _0071_;
	reg _0072_;
	reg _0073_;
	reg _0074_;
	reg _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire [7:0] _1004_;
	wire [7:0] _1005_;
	wire [9:0] _1006_;
	wire [9:0] _1007_;
	wire [9:0] _1008_;
	wire [9:0] _1009_;
	wire [4:0] _1010_;
	wire [4:0] _1011_;
	wire [4:0] _1012_;
	wire [4:0] _1013_;
	wire [8:0] _1014_;
	wire [8:0] _1015_;
	wire [8:0] _1016_;
	wire [17:0] _1017_;
	wire [31:0] _1018_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire \mchip.dut.adc_spi_clk ;
	wire \mchip.dut.adc_spi_cs_n ;
	wire \mchip.dut.adc_spi_miso ;
	wire \mchip.dut.adc_spi_mosi ;
	wire \mchip.dut.clk ;
	wire \mchip.dut.driver.a.clk ;
	reg [9:0] \mchip.dut.driver.a.counter ;
	wire [7:0] \mchip.dut.driver.a.duty_cycle ;
	reg \mchip.dut.driver.a.pwm_out ;
	wire [9:0] \mchip.dut.driver.a.switch_threshold ;
	wire \mchip.dut.driver.b.clk ;
	reg [9:0] \mchip.dut.driver.b.counter ;
	wire [7:0] \mchip.dut.driver.b.duty_cycle ;
	reg \mchip.dut.driver.b.pwm_out ;
	wire [9:0] \mchip.dut.driver.b.switch_threshold ;
	wire \mchip.dut.driver.clk ;
	reg [7:0] \mchip.dut.driver.motor_a_duty_cycle ;
	wire [7:0] \mchip.dut.driver.motor_b_duty_cycle ;
	wire \mchip.dut.driver.pwm_a ;
	wire \mchip.dut.driver.pwm_b ;
	wire [7:0] \mchip.dut.driver.setpoint ;
	wire [15:0] \mchip.dut.input_mosi_buffer ;
	wire \mchip.dut.input_spi_clk ;
	wire \mchip.dut.input_spi_cs_n ;
	wire \mchip.dut.input_spi_interface.clk.clk ;
	reg [2:0] \mchip.dut.input_spi_interface.clk.data_buffer ;
	wire \mchip.dut.input_spi_interface.clk.data_in ;
	reg \mchip.dut.input_spi_interface.clk.data_out ;
	wire \mchip.dut.input_spi_interface.cs_n.clk ;
	reg [2:0] \mchip.dut.input_spi_interface.cs_n.data_buffer ;
	wire \mchip.dut.input_spi_interface.cs_n.data_in ;
	reg \mchip.dut.input_spi_interface.cs_n.data_out ;
	wire \mchip.dut.input_spi_interface.internal_reset_n ;
	wire \mchip.dut.input_spi_interface.mosi.clk ;
	reg [2:0] \mchip.dut.input_spi_interface.mosi.data_buffer ;
	wire \mchip.dut.input_spi_interface.mosi.data_in ;
	reg \mchip.dut.input_spi_interface.mosi.data_out ;
	wire [15:0] \mchip.dut.input_spi_interface.mosi_buffer ;
	wire [4:0] \mchip.dut.input_spi_interface.mosi_buffer_counter ;
	wire \mchip.dut.input_spi_interface.spi_clk ;
	wire \mchip.dut.input_spi_interface.spi_cs_n ;
	wire \mchip.dut.input_spi_interface.spi_mosi ;
	wire \mchip.dut.input_spi_interface.sync_spi_clk ;
	wire \mchip.dut.input_spi_interface.sync_spi_cs_n ;
	wire \mchip.dut.input_spi_interface.sync_spi_mosi ;
	wire \mchip.dut.input_spi_interface.sys_clk ;
	wire \mchip.dut.input_spi_mosi ;
	reg [4:0] \mchip.dut.mcp3202.counter ;
	reg [8:0] \mchip.dut.mcp3202.done_counter ;
	wire [31:0] \mchip.dut.mcp3202.next_state ;
	reg \mchip.dut.mcp3202.reading_valid ;
	wire [11:0] \mchip.dut.mcp3202.sensor_reading ;
	reg \mchip.dut.mcp3202.spi_clk ;
	reg \mchip.dut.mcp3202.spi_cs_n ;
	wire \mchip.dut.mcp3202.spi_miso ;
	reg \mchip.dut.mcp3202.spi_mosi ;
	reg [20:0] \mchip.dut.mcp3202.state ;
	wire \mchip.dut.mcp3202.sys_clk ;
	wire [7:0] \mchip.dut.motor_setpoint ;
	wire [7:0] \mchip.dut.p ;
	wire \mchip.dut.p_cont.clk ;
	reg [8:0] \mchip.dut.p_cont.error ;
	wire [17:0] \mchip.dut.p_cont.internal_output_setpoint ;
	reg [7:0] \mchip.dut.p_cont.output_setpoint ;
	wire [7:0] \mchip.dut.p_cont.p ;
	reg [7:0] \mchip.dut.p_cont.round_reading ;
	wire [11:0] \mchip.dut.p_cont.sensor_reading ;
	wire [7:0] \mchip.dut.p_cont.setpoint ;
	wire \mchip.dut.p_setpoint_storage.address ;
	wire \mchip.dut.p_setpoint_storage.clk ;
	reg [7:0] \mchip.dut.p_setpoint_storage.p ;
	wire [7:0] \mchip.dut.p_setpoint_storage.param ;
	reg [7:0] \mchip.dut.p_setpoint_storage.setpoint ;
	wire \mchip.dut.param_address ;
	wire [7:0] \mchip.dut.param_value ;
	wire \mchip.dut.pwm_a ;
	wire \mchip.dut.pwm_b ;
	wire [11:0] \mchip.dut.sensor_reading ;
	wire [11:0] \mchip.dut.sensor_reading_captured ;
	wire \mchip.dut.sensor_reading_valid ;
	wire [7:0] \mchip.dut.setpoint ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _1004_[0] = ~\mchip.dut.p_cont.output_setpoint [0];
	assign _1016_[0] = \mchip.dut.p_cont.round_reading [0] ^ \mchip.dut.p_setpoint_storage.setpoint [0];
	assign _1004_[1] = ~\mchip.dut.p_cont.output_setpoint [1];
	assign _1004_[2] = ~\mchip.dut.p_cont.output_setpoint [2];
	assign _1004_[3] = ~\mchip.dut.p_cont.output_setpoint [3];
	assign _1004_[4] = ~\mchip.dut.p_cont.output_setpoint [4];
	assign _1004_[5] = ~\mchip.dut.p_cont.output_setpoint [5];
	assign _1004_[6] = ~\mchip.dut.p_cont.output_setpoint [6];
	assign _0419_ = \mchip.dut.mcp3202.counter [2] | \mchip.dut.mcp3202.counter [3];
	assign _0420_ = \mchip.dut.mcp3202.counter [0] | \mchip.dut.mcp3202.counter [1];
	assign _0421_ = _0420_ | _0419_;
	assign _0422_ = _0421_ | \mchip.dut.mcp3202.counter [4];
	assign _0423_ = _0422_ & ~io_in[13];
	assign _0424_ = ~\mchip.dut.mcp3202.state [20];
	assign _0425_ = \mchip.dut.mcp3202.state [19] | \mchip.dut.mcp3202.state [15];
	assign _0426_ = \mchip.dut.mcp3202.state [14] | \mchip.dut.mcp3202.state [10];
	assign _0427_ = _0426_ | _0425_;
	assign _0428_ = \mchip.dut.mcp3202.state [9] | \mchip.dut.mcp3202.state [5];
	assign _0429_ = \mchip.dut.mcp3202.state [4] | \mchip.dut.mcp3202.state [3];
	assign _0430_ = _0429_ | _0428_;
	assign _0431_ = _0430_ | _0427_;
	assign _0432_ = _0424_ & ~_0431_;
	assign _0433_ = _0423_ & ~_0432_;
	assign _0434_ = \mchip.dut.mcp3202.done_counter [0] & \mchip.dut.mcp3202.done_counter [1];
	assign _0435_ = ~(\mchip.dut.mcp3202.done_counter [2] & \mchip.dut.mcp3202.done_counter [3]);
	assign _0436_ = _0434_ & ~_0435_;
	assign _0437_ = ~(\mchip.dut.mcp3202.done_counter [6] & \mchip.dut.mcp3202.done_counter [7]);
	assign _0438_ = ~(\mchip.dut.mcp3202.done_counter [4] & \mchip.dut.mcp3202.done_counter [5]);
	assign _0439_ = ~(_0438_ | _0437_);
	assign _0440_ = ~(_0439_ & _0436_);
	assign _0441_ = \mchip.dut.mcp3202.done_counter [8] & ~_0440_;
	assign _0442_ = _0441_ | io_in[13];
	assign _0443_ = _0442_ | _0422_;
	assign _0444_ = \mchip.dut.mcp3202.state [4] & ~_0443_;
	assign _0445_ = ~(_0422_ | io_in[13]);
	assign _0446_ = ~(\mchip.dut.mcp3202.state [17] | \mchip.dut.mcp3202.state [16]);
	assign _0447_ = ~(\mchip.dut.mcp3202.state [15] | \mchip.dut.mcp3202.state [14]);
	assign _0448_ = ~(_0447_ & _0446_);
	assign _0449_ = ~(\mchip.dut.mcp3202.state [10] | \mchip.dut.mcp3202.state [9]);
	assign _0450_ = ~(\mchip.dut.mcp3202.state [5] | \mchip.dut.mcp3202.state [3]);
	assign _0451_ = ~(_0450_ & _0449_);
	assign _0452_ = ~(_0451_ | _0448_);
	assign _0453_ = _0452_ & ~\mchip.dut.mcp3202.state [18];
	assign _0454_ = _0445_ & ~_0453_;
	assign _0455_ = _0454_ | _0444_;
	assign _0046_ = _0455_ | _0433_;
	assign _0456_ = ~(\mchip.dut.mcp3202.state [2] | \mchip.dut.mcp3202.state [5]);
	assign _0457_ = \mchip.dut.mcp3202.state [8] | \mchip.dut.mcp3202.state [10];
	assign _0458_ = _0456_ & ~_0457_;
	assign _0459_ = \mchip.dut.mcp3202.state [19] | \mchip.dut.mcp3202.state [18];
	assign _0460_ = \mchip.dut.mcp3202.state [13] | \mchip.dut.mcp3202.state [15];
	assign _0461_ = _0460_ | _0459_;
	assign _0462_ = _0458_ & ~_0461_;
	assign _0463_ = _0445_ & ~_0462_;
	assign _0464_ = \mchip.dut.mcp3202.state [20] | \mchip.dut.mcp3202.state [18];
	assign _0465_ = _0464_ | _0460_;
	assign _0466_ = _0458_ & ~_0465_;
	assign _0467_ = _0423_ & ~_0466_;
	assign _0047_ = _0467_ | _0463_;
	assign _0468_ = \mchip.dut.mcp3202.state [12] | \mchip.dut.mcp3202.state [17];
	assign _0469_ = \mchip.dut.mcp3202.state [7] | \mchip.dut.mcp3202.state [1];
	assign _0470_ = _0469_ | _0468_;
	assign _0471_ = _0424_ & ~_0470_;
	assign _0472_ = _0445_ & ~_0471_;
	assign _0473_ = ~(\mchip.dut.mcp3202.state [7] | \mchip.dut.mcp3202.state [12]);
	assign _0474_ = ~(\mchip.dut.mcp3202.state [1] | \mchip.dut.mcp3202.state [4]);
	assign _0475_ = _0474_ & _0473_;
	assign _0476_ = _0475_ & ~\mchip.dut.mcp3202.state [17];
	assign _0477_ = _0423_ & ~_0476_;
	assign _0478_ = _0477_ | _0472_;
	assign _0048_ = _0478_ | _0444_;
	assign _1006_[0] = ~\mchip.dut.driver.a.counter [0];
	assign _0043_ = _0421_ | ~\mchip.dut.mcp3202.counter [4];
	assign _0479_ = ~_1018_[4];
	assign _0480_ = \mchip.dut.mcp3202.state [4] & ~_0441_;
	assign _0481_ = _0480_ | \mchip.dut.mcp3202.state [17];
	assign _0482_ = _0473_ & ~_0481_;
	assign _0483_ = \mchip.dut.mcp3202.state [1] | \mchip.dut.mcp3202.state [20];
	assign _0484_ = _0482_ & ~_0483_;
	assign _0485_ = \mchip.dut.mcp3202.state [4] | \mchip.dut.mcp3202.state [17];
	assign _0486_ = _0473_ & ~_0485_;
	assign _0487_ = \mchip.dut.mcp3202.state [15] | \mchip.dut.mcp3202.state [10];
	assign _0488_ = _0487_ | _0483_;
	assign _0489_ = _0486_ & ~_0488_;
	assign _0490_ = \mchip.dut.mcp3202.state [14] | \mchip.dut.mcp3202.state [9];
	assign _0491_ = \mchip.dut.mcp3202.state [2] | \mchip.dut.mcp3202.state [19];
	assign _0492_ = _0491_ | _0490_;
	assign _0493_ = \mchip.dut.mcp3202.state [13] | \mchip.dut.mcp3202.state [8];
	assign _0494_ = \mchip.dut.mcp3202.state [18] | \mchip.dut.mcp3202.state [5];
	assign _0495_ = _0494_ | _0493_;
	assign _0496_ = _0495_ | _0492_;
	assign _0497_ = _0489_ & ~_0496_;
	assign _0498_ = \mchip.dut.mcp3202.state [11] | \mchip.dut.mcp3202.state [6];
	assign _0499_ = \mchip.dut.mcp3202.state [16] | \mchip.dut.mcp3202.state [3];
	assign _0500_ = _0499_ | _0498_;
	assign _0501_ = _0500_ | \mchip.dut.mcp3202.state [0];
	assign _0502_ = _0497_ & ~_0501_;
	assign _0503_ = (_0502_ ? _0479_ : _0484_);
	assign _0504_ = (_0422_ ? _0479_ : _0503_);
	assign _0505_ = ~_1018_[1];
	assign _0506_ = _0493_ | _0490_;
	assign _0507_ = _0487_ | ~_0473_;
	assign _0508_ = _0507_ | _0506_;
	assign _0509_ = ~(_0508_ | _0498_);
	assign _0510_ = (_0502_ ? _0505_ : _0509_);
	assign _0511_ = (_0422_ ? _0505_ : _0510_);
	assign _0512_ = \mchip.dut.mcp3202.state [1] | \mchip.dut.mcp3202.state [10];
	assign _0513_ = _0512_ | \mchip.dut.mcp3202.state [7];
	assign _0514_ = \mchip.dut.mcp3202.state [2] | \mchip.dut.mcp3202.state [9];
	assign _0515_ = \mchip.dut.mcp3202.state [8] | \mchip.dut.mcp3202.state [5];
	assign _0516_ = _0515_ | _0514_;
	assign _0517_ = _0516_ | _0513_;
	assign _0518_ = \mchip.dut.mcp3202.state [6] | \mchip.dut.mcp3202.state [3];
	assign _0519_ = _0518_ | \mchip.dut.mcp3202.state [0];
	assign _0520_ = _0519_ | _0517_;
	assign _0521_ = (_0502_ ? _1018_[0] : _0520_);
	assign _0522_ = (_0422_ ? _1018_[0] : _0521_);
	assign _0523_ = ~(_0522_ & _0511_);
	assign _0524_ = ~_1018_[3];
	assign _0525_ = _0495_ | _0491_;
	assign _0526_ = ~(_0525_ | _0487_);
	assign _0527_ = (_0502_ ? _0524_ : _0526_);
	assign _0528_ = (_0422_ ? _0524_ : _0527_);
	assign _0529_ = ~_1018_[2];
	assign _0530_ = _0494_ | _0490_;
	assign _0531_ = _0487_ | _0481_;
	assign _0532_ = _0531_ | _0530_;
	assign _0533_ = ~(_0532_ | _0499_);
	assign _0534_ = (_0502_ ? _0529_ : _0533_);
	assign _0535_ = (_0422_ ? _0529_ : _0534_);
	assign _0536_ = _0528_ | ~_0535_;
	assign _0537_ = _0536_ | _0523_;
	assign _0538_ = _0537_ | ~_0504_;
	assign _0539_ = _0522_ | _0511_;
	assign _0540_ = _0535_ | ~_0528_;
	assign _0541_ = _0540_ | _0539_;
	assign _0542_ = _0504_ & ~_0541_;
	assign _0543_ = _0538_ & ~_0542_;
	assign _0544_ = _0511_ | ~_0522_;
	assign _0545_ = _0544_ | _0540_;
	assign _0546_ = _0504_ & ~_0545_;
	assign _0547_ = _0522_ | ~_0511_;
	assign _0548_ = _0547_ | _0536_;
	assign _0549_ = _0504_ & ~_0548_;
	assign _0550_ = _0549_ | _0546_;
	assign _0551_ = _0543_ & ~_0550_;
	assign _0552_ = _0535_ | _0528_;
	assign _0553_ = _0552_ | _0523_;
	assign _0554_ = _0504_ & ~_0553_;
	assign _0555_ = _0552_ | _0547_;
	assign _0556_ = _0504_ & ~_0555_;
	assign _0557_ = _0556_ | _0554_;
	assign _0558_ = _0544_ | _0536_;
	assign _0559_ = _0504_ & ~_0558_;
	assign _0560_ = _0539_ | _0536_;
	assign _0561_ = _0504_ & ~_0560_;
	assign _0562_ = _0561_ | _0559_;
	assign _0563_ = _0562_ | _0557_;
	assign _0564_ = _0551_ & ~_0563_;
	assign _0565_ = _0552_ | _0539_;
	assign _0566_ = _0504_ & ~_0565_;
	assign _0567_ = _0043_ | ~_0566_;
	assign _0028_ = _0564_ & ~_0567_;
	assign _0568_ = _0556_ | ~_0554_;
	assign _0569_ = _0568_ | _0562_;
	assign _0570_ = _0569_ | ~_0551_;
	assign _0029_ = ~(_0570_ | _0043_);
	assign _0571_ = _0043_ | ~_0556_;
	assign _0572_ = _0571_ | _0562_;
	assign _0030_ = _0551_ & ~_0572_;
	assign _0573_ = _0561_ | ~_0559_;
	assign _0574_ = _0573_ | _0043_;
	assign _0031_ = _0551_ & ~_0574_;
	assign _0575_ = _0043_ | ~_0561_;
	assign _0032_ = _0551_ & ~_0575_;
	assign _0576_ = _0542_ | _0538_;
	assign _0577_ = _0576_ | _0550_;
	assign _0021_ = ~(_0577_ | _0043_);
	assign _0578_ = ~(_0546_ | _0542_);
	assign _0579_ = _0043_ | ~_0549_;
	assign _0022_ = _0578_ & ~_0579_;
	assign _0580_ = _0542_ | ~_0546_;
	assign _0023_ = ~(_0580_ | _0043_);
	assign _0024_ = _0542_ & ~_0043_;
	assign _0581_ = ~(\mchip.dut.mcp3202.state [19] | \mchip.dut.mcp3202.state [20]);
	assign _0582_ = \mchip.dut.mcp3202.state [18] | \mchip.dut.mcp3202.state [17];
	assign _0583_ = \mchip.dut.mcp3202.state [16] | \mchip.dut.mcp3202.state [10];
	assign _0584_ = _0583_ | _0582_;
	assign _0585_ = \mchip.dut.mcp3202.state [6] | \mchip.dut.mcp3202.state [7];
	assign _0586_ = \mchip.dut.mcp3202.state [8] | \mchip.dut.mcp3202.state [9];
	assign _0587_ = _0586_ | _0585_;
	assign _0588_ = _0587_ | _0584_;
	assign _0589_ = _0581_ & ~_0588_;
	assign _0590_ = _0423_ & ~_0589_;
	assign _0591_ = \mchip.dut.mcp3202.state [12] | \mchip.dut.mcp3202.state [13];
	assign _0592_ = \mchip.dut.mcp3202.state [11] | \mchip.dut.mcp3202.state [10];
	assign _0593_ = _0592_ | _0591_;
	assign _0594_ = _0593_ | _0587_;
	assign _0595_ = _0447_ & ~_0594_;
	assign _0596_ = _0445_ & ~_0595_;
	assign _0045_ = _0596_ | _0590_;
	assign _0597_ = \mchip.dut.mcp3202.state [16] | \mchip.dut.mcp3202.state [15];
	assign _0598_ = _0597_ | _0582_;
	assign _0599_ = \mchip.dut.mcp3202.state [13] | \mchip.dut.mcp3202.state [14];
	assign _0600_ = \mchip.dut.mcp3202.state [11] | \mchip.dut.mcp3202.state [12];
	assign _0601_ = _0600_ | _0599_;
	assign _0602_ = _0601_ | _0598_;
	assign _0603_ = _0581_ & ~_0602_;
	assign _0604_ = _0423_ & ~_0603_;
	assign _0605_ = \mchip.dut.mcp3202.state [7] | \mchip.dut.mcp3202.state [8];
	assign _0606_ = \mchip.dut.mcp3202.state [6] | \mchip.dut.mcp3202.state [5];
	assign _0607_ = _0606_ | _0605_;
	assign _0608_ = \mchip.dut.mcp3202.state [2] | \mchip.dut.mcp3202.state [3];
	assign _0609_ = \mchip.dut.mcp3202.state [0] | \mchip.dut.mcp3202.state [1];
	assign _0610_ = _0609_ | _0608_;
	assign _0611_ = _0610_ | _0607_;
	assign _0612_ = _0449_ & ~_0611_;
	assign _0613_ = _0445_ & ~_0612_;
	assign _0044_ = _0613_ | _0604_;
	assign _0614_ = _0423_ & ~_0424_;
	assign _0615_ = _0445_ & \mchip.dut.mcp3202.state [10];
	assign _0012_ = _0615_ | _0614_;
	assign _0616_ = _0423_ & \mchip.dut.mcp3202.state [19];
	assign _0617_ = _0445_ & \mchip.dut.mcp3202.state [9];
	assign _0010_ = _0617_ | _0616_;
	assign _1008_[0] = ~\mchip.dut.driver.b.counter [0];
	assign _0618_ = _0423_ & \mchip.dut.mcp3202.state [18];
	assign _0619_ = _0445_ & \mchip.dut.mcp3202.state [8];
	assign _0009_ = _0619_ | _0618_;
	assign _0620_ = _0423_ & \mchip.dut.mcp3202.state [17];
	assign _0621_ = _0445_ & \mchip.dut.mcp3202.state [7];
	assign _0008_ = _0621_ | _0620_;
	assign _0622_ = ~(_0535_ & _0528_);
	assign _0623_ = _0622_ | _0523_;
	assign _0624_ = ~(_0623_ | _0504_);
	assign _0625_ = _0622_ | _0539_;
	assign _0626_ = _0625_ | _0504_;
	assign _0627_ = ~(_0622_ | _0547_);
	assign _0628_ = _0627_ & ~_0504_;
	assign _0629_ = _0628_ | _0626_;
	assign _0630_ = _0552_ | _0544_;
	assign _0631_ = _0504_ & ~_0630_;
	assign _0632_ = _0631_ | _0566_;
	assign _0633_ = _0632_ | _0629_;
	assign _0634_ = _0633_ | _0624_;
	assign _0027_ = _0564_ & ~_0634_;
	assign _0635_ = _0423_ & \mchip.dut.mcp3202.state [16];
	assign _0636_ = _0445_ & \mchip.dut.mcp3202.state [6];
	assign _0007_ = _0636_ | _0635_;
	assign _0637_ = _0423_ & \mchip.dut.mcp3202.state [15];
	assign _0638_ = _0445_ & \mchip.dut.mcp3202.state [5];
	assign _0006_ = _0638_ | _0637_;
	assign _0639_ = _0423_ & \mchip.dut.mcp3202.state [14];
	assign _0640_ = _0445_ & \mchip.dut.mcp3202.state [3];
	assign _0005_ = _0640_ | _0639_;
	assign _0641_ = _0423_ & \mchip.dut.mcp3202.state [13];
	assign _0642_ = _0445_ & \mchip.dut.mcp3202.state [2];
	assign _0004_ = _0642_ | _0641_;
	assign _0643_ = _0423_ & \mchip.dut.mcp3202.state [12];
	assign _0644_ = _0445_ & \mchip.dut.mcp3202.state [1];
	assign _0003_ = _0644_ | _0643_;
	assign _0645_ = _0423_ & \mchip.dut.mcp3202.state [11];
	assign _0646_ = _0445_ & \mchip.dut.mcp3202.state [0];
	assign _0002_ = _0646_ | _0645_;
	assign _0647_ = _0423_ & \mchip.dut.mcp3202.state [10];
	assign _0648_ = _0445_ & \mchip.dut.mcp3202.state [15];
	assign _0001_ = _0648_ | _0647_;
	assign _0649_ = _0423_ & \mchip.dut.mcp3202.state [9];
	assign _0650_ = _0445_ & \mchip.dut.mcp3202.state [14];
	assign _0020_ = _0650_ | _0649_;
	assign _0651_ = _0423_ & \mchip.dut.mcp3202.state [8];
	assign _0652_ = _0445_ & \mchip.dut.mcp3202.state [13];
	assign _0019_ = _0652_ | _0651_;
	assign _0653_ = _0423_ & \mchip.dut.mcp3202.state [7];
	assign _0654_ = _0445_ & \mchip.dut.mcp3202.state [12];
	assign _0018_ = _0654_ | _0653_;
	assign _0655_ = _0423_ & \mchip.dut.mcp3202.state [6];
	assign _0656_ = _0445_ & \mchip.dut.mcp3202.state [11];
	assign _0017_ = _0656_ | _0655_;
	assign _0657_ = _0423_ & \mchip.dut.mcp3202.state [5];
	assign _0658_ = _0445_ & \mchip.dut.mcp3202.state [18];
	assign _0016_ = _0658_ | _0657_;
	assign _0659_ = io_in[13] | ~_0441_;
	assign _0660_ = _0659_ | _0422_;
	assign _0661_ = \mchip.dut.mcp3202.state [4] & ~_0660_;
	assign _0662_ = _0423_ & \mchip.dut.mcp3202.state [0];
	assign _0663_ = _0662_ | io_in[13];
	assign _0000_ = _0663_ | _0661_;
	assign \mchip.dut.input_spi_interface.internal_reset_n  = _0075_ & ~io_in[13];
	assign _0664_ = \mchip.dut.input_spi_interface.internal_reset_n  & _0064_;
	assign _0665_ = \mchip.dut.input_spi_interface.internal_reset_n  & _0063_;
	assign _0666_ = ~(_0665_ | _0664_);
	assign _0667_ = \mchip.dut.input_spi_interface.internal_reset_n  & _0062_;
	assign _0668_ = \mchip.dut.input_spi_interface.internal_reset_n  & _0061_;
	assign _0669_ = _0668_ | _0667_;
	assign _0670_ = _0669_ | ~_0666_;
	assign _0671_ = \mchip.dut.input_spi_interface.internal_reset_n  & _0065_;
	assign _0672_ = _0671_ & ~_0670_;
	assign _0673_ = \mchip.dut.input_spi_interface.internal_reset_n  & _0074_;
	assign _0025_ = _0672_ & ~_0673_;
	assign _0674_ = _0423_ & \mchip.dut.mcp3202.state [4];
	assign _0675_ = _0445_ & \mchip.dut.mcp3202.state [17];
	assign _0676_ = _0675_ | _0674_;
	assign _0015_ = _0676_ | _0444_;
	assign _0677_ = _0504_ & ~_0623_;
	assign _0678_ = _0504_ & ~_0625_;
	assign _0034_ = _0678_ | _0677_;
	assign _0679_ = \mchip.dut.input_spi_interface.cs_n.data_buffer [0] & \mchip.dut.input_spi_interface.cs_n.data_buffer [1];
	assign _0040_ = ~(_0679_ & \mchip.dut.input_spi_interface.cs_n.data_buffer [2]);
	assign _0680_ = \mchip.dut.input_spi_interface.mosi.data_buffer [0] & \mchip.dut.input_spi_interface.mosi.data_buffer [1];
	assign _0041_ = ~(_0680_ & \mchip.dut.input_spi_interface.mosi.data_buffer [2]);
	assign _0681_ = \mchip.dut.input_spi_interface.clk.data_buffer [0] & \mchip.dut.input_spi_interface.clk.data_buffer [1];
	assign _0042_ = ~(_0681_ & \mchip.dut.input_spi_interface.clk.data_buffer [2]);
	assign _0682_ = _0423_ & \mchip.dut.mcp3202.state [3];
	assign _0683_ = _0445_ & \mchip.dut.mcp3202.state [16];
	assign _0014_ = _0683_ | _0682_;
	assign _0033_ = \mchip.dut.mcp3202.state [17] | io_in[13];
	assign _0684_ = _0423_ & \mchip.dut.mcp3202.state [2];
	assign _0685_ = _0445_ & \mchip.dut.mcp3202.state [19];
	assign _0013_ = _0685_ | _0684_;
	assign _0026_ = _0673_ & _0672_;
	assign _0686_ = _0445_ & ~_0424_;
	assign _0687_ = _0423_ & \mchip.dut.mcp3202.state [1];
	assign _0011_ = _0687_ | _0686_;
	assign _0688_ = \mchip.dut.input_spi_interface.cs_n.data_buffer [0] | \mchip.dut.input_spi_interface.cs_n.data_buffer [1];
	assign _0037_ = _0688_ | \mchip.dut.input_spi_interface.cs_n.data_buffer [2];
	assign _0689_ = \mchip.dut.input_spi_interface.mosi.data_buffer [0] | \mchip.dut.input_spi_interface.mosi.data_buffer [1];
	assign _0038_ = _0689_ | \mchip.dut.input_spi_interface.mosi.data_buffer [2];
	assign _0690_ = \mchip.dut.input_spi_interface.clk.data_buffer [0] | \mchip.dut.input_spi_interface.clk.data_buffer [1];
	assign _0039_ = _0690_ | \mchip.dut.input_spi_interface.clk.data_buffer [2];
	assign _0691_ = ~(_0547_ | _0540_);
	assign _0050_ = (_0504_ ? _0627_ : _0691_);
	assign _0692_ = _0691_ & _0504_;
	assign _0693_ = _0622_ | _0544_;
	assign _0694_ = _0504_ & ~_0693_;
	assign _0051_ = _0692_ & ~_0694_;
	assign _0695_ = \mchip.dut.sensor_reading_captured [11] & \mchip.dut.sensor_reading_captured [10];
	assign _0696_ = ~(\mchip.dut.sensor_reading_captured [8] & \mchip.dut.sensor_reading_captured [9]);
	assign _0697_ = _0695_ & ~_0696_;
	assign _0698_ = \mchip.dut.sensor_reading_captured [4] & \mchip.dut.sensor_reading_captured [5];
	assign _0699_ = \mchip.dut.sensor_reading_captured [6] & \mchip.dut.sensor_reading_captured [7];
	assign _0700_ = ~(_0699_ & _0698_);
	assign _0701_ = _0700_ | ~_0697_;
	assign _0702_ = ~(_0701_ & \mchip.dut.sensor_reading_captured [3]);
	assign _0052_ = ~(_0702_ ^ \mchip.dut.sensor_reading_captured [4]);
	assign _0703_ = \mchip.dut.sensor_reading_captured [4] ^ \mchip.dut.sensor_reading_captured [5];
	assign _0053_ = (_0702_ ? \mchip.dut.sensor_reading_captured [5] : _0703_);
	assign _0704_ = _0698_ ^ \mchip.dut.sensor_reading_captured [6];
	assign _0054_ = (_0702_ ? \mchip.dut.sensor_reading_captured [6] : _0704_);
	assign _0705_ = _0698_ & \mchip.dut.sensor_reading_captured [6];
	assign _0706_ = _0705_ ^ \mchip.dut.sensor_reading_captured [7];
	assign _0055_ = (_0702_ ? \mchip.dut.sensor_reading_captured [7] : _0706_);
	assign _0707_ = ~(_0700_ ^ \mchip.dut.sensor_reading_captured [8]);
	assign _0056_ = (_0702_ ? \mchip.dut.sensor_reading_captured [8] : _0707_);
	assign _0708_ = \mchip.dut.sensor_reading_captured [8] & ~_0700_;
	assign _0709_ = _0708_ ^ \mchip.dut.sensor_reading_captured [9];
	assign _0057_ = (_0702_ ? \mchip.dut.sensor_reading_captured [9] : _0709_);
	assign _0710_ = ~(_0700_ | _0696_);
	assign _0711_ = _0710_ ^ \mchip.dut.sensor_reading_captured [10];
	assign _0058_ = (_0702_ ? \mchip.dut.sensor_reading_captured [10] : _0711_);
	assign _0712_ = _0710_ & \mchip.dut.sensor_reading_captured [10];
	assign _0713_ = _0712_ ^ \mchip.dut.sensor_reading_captured [11];
	assign _0059_ = (_0702_ ? \mchip.dut.sensor_reading_captured [11] : _0713_);
	assign _0714_ = ~(_0060_ | io_in[13]);
	assign _0049_ = _0714_ | \mchip.dut.input_spi_interface.cs_n.data_out ;
	assign _1014_[0] = ~\mchip.dut.mcp3202.done_counter [0];
	assign _1010_[0] = ~_0668_;
	assign _1012_[0] = ~\mchip.dut.mcp3202.counter [0];
	assign _0715_ = ~(\mchip.dut.driver.a.counter [9] ^ \mchip.dut.driver.motor_a_duty_cycle [7]);
	assign _0716_ = \mchip.dut.driver.a.counter [8] ^ \mchip.dut.driver.motor_a_duty_cycle [6];
	assign _0717_ = _0715_ & ~_0716_;
	assign _0718_ = \mchip.dut.driver.motor_a_duty_cycle [4] ^ \mchip.dut.driver.a.counter [6];
	assign _0719_ = \mchip.dut.driver.a.counter [7] ^ \mchip.dut.driver.motor_a_duty_cycle [5];
	assign _0720_ = _0719_ | _0718_;
	assign _0721_ = ~(\mchip.dut.driver.a.counter [5] ^ \mchip.dut.driver.motor_a_duty_cycle [3]);
	assign _0722_ = \mchip.dut.driver.a.counter [4] ^ \mchip.dut.driver.motor_a_duty_cycle [2];
	assign _0723_ = _0721_ & ~_0722_;
	assign _0724_ = _0720_ | ~_0723_;
	assign _0725_ = \mchip.dut.driver.motor_a_duty_cycle [0] ^ \mchip.dut.driver.a.counter [2];
	assign _0726_ = \mchip.dut.driver.a.counter [3] ^ \mchip.dut.driver.motor_a_duty_cycle [1];
	assign _0727_ = _0726_ | _0725_;
	assign _0728_ = \mchip.dut.driver.a.counter [1] | \mchip.dut.driver.a.counter [0];
	assign _0729_ = _0728_ | _0727_;
	assign _0730_ = _0729_ | _0724_;
	assign _0731_ = _0717_ & ~_0730_;
	assign _0732_ = \mchip.dut.driver.motor_a_duty_cycle [7] | ~\mchip.dut.driver.a.counter [9];
	assign _0733_ = \mchip.dut.driver.motor_a_duty_cycle [6] | ~\mchip.dut.driver.a.counter [8];
	assign _0734_ = _0715_ & ~_0733_;
	assign _0735_ = _0732_ & ~_0734_;
	assign _0736_ = \mchip.dut.driver.motor_a_duty_cycle [5] | ~\mchip.dut.driver.a.counter [7];
	assign _0737_ = \mchip.dut.driver.a.counter [6] & ~\mchip.dut.driver.motor_a_duty_cycle [4];
	assign _0738_ = _0737_ & ~_0719_;
	assign _0739_ = _0736_ & ~_0738_;
	assign _0740_ = _0717_ & ~_0739_;
	assign _0741_ = _0735_ & ~_0740_;
	assign _0742_ = _0717_ & ~_0720_;
	assign _0743_ = \mchip.dut.driver.motor_a_duty_cycle [3] | ~\mchip.dut.driver.a.counter [5];
	assign _0744_ = \mchip.dut.driver.motor_a_duty_cycle [2] | ~\mchip.dut.driver.a.counter [4];
	assign _0745_ = _0721_ & ~_0744_;
	assign _0746_ = _0743_ & ~_0745_;
	assign _0747_ = \mchip.dut.driver.motor_a_duty_cycle [1] | ~\mchip.dut.driver.a.counter [3];
	assign _0748_ = \mchip.dut.driver.a.counter [2] | ~\mchip.dut.driver.motor_a_duty_cycle [0];
	assign _0749_ = _0748_ & ~_0726_;
	assign _0750_ = _0747_ & ~_0749_;
	assign _0751_ = _0723_ & ~_0750_;
	assign _0752_ = _0746_ & ~_0751_;
	assign _0753_ = _0742_ & ~_0752_;
	assign _0754_ = _0741_ & ~_0753_;
	assign _0036_ = _0754_ | _0731_;
	assign _0755_ = ~(\mchip.dut.driver.b.counter [9] ^ \mchip.dut.driver.motor_b_duty_cycle [7]);
	assign _0756_ = \mchip.dut.driver.b.counter [8] ^ \mchip.dut.driver.motor_b_duty_cycle [6];
	assign _0757_ = _0755_ & ~_0756_;
	assign _0758_ = \mchip.dut.driver.motor_b_duty_cycle [4] ^ \mchip.dut.driver.b.counter [6];
	assign _0759_ = \mchip.dut.driver.b.counter [7] ^ \mchip.dut.driver.motor_b_duty_cycle [5];
	assign _0760_ = _0759_ | _0758_;
	assign _0761_ = ~(\mchip.dut.driver.b.counter [5] ^ \mchip.dut.driver.motor_b_duty_cycle [3]);
	assign _0762_ = \mchip.dut.driver.b.counter [4] ^ \mchip.dut.driver.motor_b_duty_cycle [2];
	assign _0763_ = _0761_ & ~_0762_;
	assign _0764_ = _0760_ | ~_0763_;
	assign _0765_ = \mchip.dut.driver.b.counter [2] ^ \mchip.dut.driver.motor_a_duty_cycle [0];
	assign _0766_ = \mchip.dut.driver.b.counter [3] ^ \mchip.dut.driver.motor_b_duty_cycle [1];
	assign _0767_ = _0766_ | _0765_;
	assign _0768_ = \mchip.dut.driver.b.counter [1] | \mchip.dut.driver.b.counter [0];
	assign _0769_ = _0768_ | _0767_;
	assign _0770_ = _0769_ | _0764_;
	assign _0771_ = _0757_ & ~_0770_;
	assign _0772_ = \mchip.dut.driver.motor_b_duty_cycle [7] | ~\mchip.dut.driver.b.counter [9];
	assign _0773_ = \mchip.dut.driver.motor_b_duty_cycle [6] | ~\mchip.dut.driver.b.counter [8];
	assign _0774_ = _0755_ & ~_0773_;
	assign _0775_ = _0772_ & ~_0774_;
	assign _0776_ = \mchip.dut.driver.motor_b_duty_cycle [5] | ~\mchip.dut.driver.b.counter [7];
	assign _0777_ = \mchip.dut.driver.b.counter [6] & ~\mchip.dut.driver.motor_b_duty_cycle [4];
	assign _0778_ = _0777_ & ~_0759_;
	assign _0779_ = _0776_ & ~_0778_;
	assign _0780_ = _0757_ & ~_0779_;
	assign _0781_ = _0775_ & ~_0780_;
	assign _0782_ = _0757_ & ~_0760_;
	assign _0783_ = \mchip.dut.driver.motor_b_duty_cycle [3] | ~\mchip.dut.driver.b.counter [5];
	assign _0784_ = \mchip.dut.driver.motor_b_duty_cycle [2] | ~\mchip.dut.driver.b.counter [4];
	assign _0785_ = _0761_ & ~_0784_;
	assign _0786_ = _0783_ & ~_0785_;
	assign _0787_ = \mchip.dut.driver.motor_b_duty_cycle [1] | ~\mchip.dut.driver.b.counter [3];
	assign _0788_ = \mchip.dut.driver.b.counter [2] | ~\mchip.dut.driver.motor_a_duty_cycle [0];
	assign _0789_ = _0788_ & ~_0766_;
	assign _0790_ = _0787_ & ~_0789_;
	assign _0791_ = _0763_ & ~_0790_;
	assign _0792_ = _0786_ & ~_0791_;
	assign _0793_ = _0782_ & ~_0792_;
	assign _0794_ = _0781_ & ~_0793_;
	assign _0035_ = _0794_ | _0771_;
	assign _1009_[1] = \mchip.dut.driver.b.counter [1] ^ \mchip.dut.driver.b.counter [0];
	assign _0795_ = \mchip.dut.driver.b.counter [1] & \mchip.dut.driver.b.counter [0];
	assign _1009_[2] = _0795_ ^ \mchip.dut.driver.b.counter [2];
	assign _0796_ = _0795_ & \mchip.dut.driver.b.counter [2];
	assign _1009_[3] = _0796_ ^ \mchip.dut.driver.b.counter [3];
	assign _0797_ = ~(\mchip.dut.driver.b.counter [2] & \mchip.dut.driver.b.counter [3]);
	assign _0798_ = _0795_ & ~_0797_;
	assign _1009_[4] = _0798_ ^ \mchip.dut.driver.b.counter [4];
	assign _0799_ = _0798_ & \mchip.dut.driver.b.counter [4];
	assign _1009_[5] = _0799_ ^ \mchip.dut.driver.b.counter [5];
	assign _0800_ = ~(\mchip.dut.driver.b.counter [4] & \mchip.dut.driver.b.counter [5]);
	assign _0801_ = _0798_ & ~_0800_;
	assign _1009_[6] = _0801_ ^ \mchip.dut.driver.b.counter [6];
	assign _0802_ = _0801_ & \mchip.dut.driver.b.counter [6];
	assign _1009_[7] = _0802_ ^ \mchip.dut.driver.b.counter [7];
	assign _0803_ = ~(\mchip.dut.driver.b.counter [6] & \mchip.dut.driver.b.counter [7]);
	assign _0804_ = _0803_ | _0800_;
	assign _0805_ = _0798_ & ~_0804_;
	assign _1009_[8] = _0805_ ^ \mchip.dut.driver.b.counter [8];
	assign _0806_ = _0805_ & \mchip.dut.driver.b.counter [8];
	assign _1009_[9] = _0806_ ^ \mchip.dut.driver.b.counter [9];
	assign _1005_[1] = ~(\mchip.dut.p_cont.output_setpoint [1] ^ \mchip.dut.p_cont.output_setpoint [0]);
	assign _0807_ = ~(\mchip.dut.p_cont.output_setpoint [1] | \mchip.dut.p_cont.output_setpoint [0]);
	assign _1005_[2] = _0807_ ^ \mchip.dut.p_cont.output_setpoint [2];
	assign _0808_ = _0807_ & ~\mchip.dut.p_cont.output_setpoint [2];
	assign _1005_[3] = _0808_ ^ \mchip.dut.p_cont.output_setpoint [3];
	assign _0809_ = \mchip.dut.p_cont.output_setpoint [3] | \mchip.dut.p_cont.output_setpoint [2];
	assign _0810_ = _0807_ & ~_0809_;
	assign _1005_[4] = _0810_ ^ \mchip.dut.p_cont.output_setpoint [4];
	assign _0811_ = _0810_ & ~\mchip.dut.p_cont.output_setpoint [4];
	assign _1005_[5] = _0811_ ^ \mchip.dut.p_cont.output_setpoint [5];
	assign _0812_ = \mchip.dut.p_cont.output_setpoint [5] | \mchip.dut.p_cont.output_setpoint [4];
	assign _0813_ = _0810_ & ~_0812_;
	assign _1005_[6] = _0813_ ^ \mchip.dut.p_cont.output_setpoint [6];
	assign _0814_ = ~(_0813_ & _1004_[6]);
	assign _1005_[7] = _0814_ ^ \mchip.dut.p_cont.output_setpoint [7];
	assign _1015_[1] = \mchip.dut.mcp3202.done_counter [0] ^ \mchip.dut.mcp3202.done_counter [1];
	assign _1015_[2] = _0434_ ^ \mchip.dut.mcp3202.done_counter [2];
	assign _0815_ = _0434_ & \mchip.dut.mcp3202.done_counter [2];
	assign _1015_[3] = _0815_ ^ \mchip.dut.mcp3202.done_counter [3];
	assign _1015_[4] = _0436_ ^ \mchip.dut.mcp3202.done_counter [4];
	assign _0816_ = _0436_ & \mchip.dut.mcp3202.done_counter [4];
	assign _1015_[5] = _0816_ ^ \mchip.dut.mcp3202.done_counter [5];
	assign _0817_ = _0436_ & ~_0438_;
	assign _1015_[6] = _0817_ ^ \mchip.dut.mcp3202.done_counter [6];
	assign _0818_ = _0817_ & \mchip.dut.mcp3202.done_counter [6];
	assign _1015_[7] = _0818_ ^ \mchip.dut.mcp3202.done_counter [7];
	assign _1015_[8] = ~(_0440_ ^ \mchip.dut.mcp3202.done_counter [8]);
	assign _1007_[1] = \mchip.dut.driver.a.counter [1] ^ \mchip.dut.driver.a.counter [0];
	assign _0819_ = \mchip.dut.driver.a.counter [1] & \mchip.dut.driver.a.counter [0];
	assign _1007_[2] = _0819_ ^ \mchip.dut.driver.a.counter [2];
	assign _0820_ = _0819_ & \mchip.dut.driver.a.counter [2];
	assign _1007_[3] = _0820_ ^ \mchip.dut.driver.a.counter [3];
	assign _0821_ = ~(\mchip.dut.driver.a.counter [2] & \mchip.dut.driver.a.counter [3]);
	assign _0822_ = _0819_ & ~_0821_;
	assign _1007_[4] = _0822_ ^ \mchip.dut.driver.a.counter [4];
	assign _0823_ = _0822_ & \mchip.dut.driver.a.counter [4];
	assign _1007_[5] = _0823_ ^ \mchip.dut.driver.a.counter [5];
	assign _0824_ = ~(\mchip.dut.driver.a.counter [4] & \mchip.dut.driver.a.counter [5]);
	assign _0825_ = _0822_ & ~_0824_;
	assign _1007_[6] = _0825_ ^ \mchip.dut.driver.a.counter [6];
	assign _0826_ = _0825_ & \mchip.dut.driver.a.counter [6];
	assign _1007_[7] = _0826_ ^ \mchip.dut.driver.a.counter [7];
	assign _0827_ = ~(\mchip.dut.driver.a.counter [6] & \mchip.dut.driver.a.counter [7]);
	assign _0828_ = _0827_ | _0824_;
	assign _0829_ = _0822_ & ~_0828_;
	assign _1007_[8] = _0829_ ^ \mchip.dut.driver.a.counter [8];
	assign _0830_ = _0829_ & \mchip.dut.driver.a.counter [8];
	assign _1007_[9] = _0830_ ^ \mchip.dut.driver.a.counter [9];
	assign _0831_ = \mchip.dut.p_setpoint_storage.setpoint [0] | ~\mchip.dut.p_cont.round_reading [0];
	assign _0832_ = ~(\mchip.dut.p_cont.round_reading [1] ^ \mchip.dut.p_setpoint_storage.setpoint [1]);
	assign _1016_[1] = _0832_ ^ _0831_;
	assign _0833_ = \mchip.dut.p_setpoint_storage.setpoint [1] & ~\mchip.dut.p_cont.round_reading [1];
	assign _0834_ = _0832_ & _0831_;
	assign _0835_ = _0834_ | _0833_;
	assign _0836_ = ~(\mchip.dut.p_cont.round_reading [2] ^ \mchip.dut.p_setpoint_storage.setpoint [2]);
	assign _1016_[2] = _0836_ ^ _0835_;
	assign _0837_ = \mchip.dut.p_setpoint_storage.setpoint [2] & ~\mchip.dut.p_cont.round_reading [2];
	assign _0838_ = _0836_ & _0835_;
	assign _0839_ = _0838_ | _0837_;
	assign _0840_ = ~(\mchip.dut.p_cont.round_reading [3] ^ \mchip.dut.p_setpoint_storage.setpoint [3]);
	assign _1016_[3] = _0840_ ^ _0839_;
	assign _0841_ = \mchip.dut.p_setpoint_storage.setpoint [3] & ~\mchip.dut.p_cont.round_reading [3];
	assign _0842_ = _0840_ & _0837_;
	assign _0843_ = _0842_ | _0841_;
	assign _0844_ = ~(_0840_ & _0836_);
	assign _0845_ = _0835_ & ~_0844_;
	assign _0846_ = _0845_ | _0843_;
	assign _0847_ = ~(\mchip.dut.p_cont.round_reading [4] ^ \mchip.dut.p_setpoint_storage.setpoint [4]);
	assign _1016_[4] = _0847_ ^ _0846_;
	assign _0848_ = \mchip.dut.p_setpoint_storage.setpoint [4] & ~\mchip.dut.p_cont.round_reading [4];
	assign _0849_ = _0847_ & _0846_;
	assign _0850_ = _0849_ | _0848_;
	assign _0851_ = ~(\mchip.dut.p_cont.round_reading [5] ^ \mchip.dut.p_setpoint_storage.setpoint [5]);
	assign _1016_[5] = _0851_ ^ _0850_;
	assign _0852_ = \mchip.dut.p_setpoint_storage.setpoint [5] & ~\mchip.dut.p_cont.round_reading [5];
	assign _0853_ = _0851_ & _0848_;
	assign _0854_ = _0853_ | _0852_;
	assign _0855_ = ~(_0851_ & _0847_);
	assign _0856_ = _0846_ & ~_0855_;
	assign _0857_ = _0856_ | _0854_;
	assign _0858_ = ~(\mchip.dut.p_cont.round_reading [6] ^ \mchip.dut.p_setpoint_storage.setpoint [6]);
	assign _1016_[6] = _0858_ ^ _0857_;
	assign _0859_ = \mchip.dut.p_setpoint_storage.setpoint [6] & ~\mchip.dut.p_cont.round_reading [6];
	assign _0860_ = _0858_ & _0857_;
	assign _0861_ = _0860_ | _0859_;
	assign _0862_ = ~(\mchip.dut.p_cont.round_reading [7] ^ \mchip.dut.p_setpoint_storage.setpoint [7]);
	assign _1016_[7] = _0862_ ^ _0861_;
	assign _0863_ = \mchip.dut.p_cont.round_reading [7] | ~\mchip.dut.p_setpoint_storage.setpoint [7];
	assign _0864_ = _0862_ & _0859_;
	assign _0865_ = _0863_ & ~_0864_;
	assign _0866_ = ~(_0862_ & _0858_);
	assign _0867_ = _0854_ & ~_0866_;
	assign _0868_ = _0865_ & ~_0867_;
	assign _0869_ = _0866_ | _0855_;
	assign _0870_ = _0846_ & ~_0869_;
	assign _0871_ = _0870_ | ~_0868_;
	assign _1016_[8] = _0871_ ^ _0862_;
	assign _1011_[1] = _0668_ ^ _0667_;
	assign _0872_ = _0668_ & _0667_;
	assign _1011_[2] = _0872_ ^ _0665_;
	assign _0873_ = _0872_ & _0665_;
	assign _1011_[3] = _0873_ ^ _0664_;
	assign _0874_ = ~(_0665_ & _0664_);
	assign _0875_ = _0872_ & ~_0874_;
	assign _1011_[4] = _0875_ ^ _0671_;
	assign _1013_[1] = \mchip.dut.mcp3202.counter [0] ^ \mchip.dut.mcp3202.counter [1];
	assign _0876_ = \mchip.dut.mcp3202.counter [0] & \mchip.dut.mcp3202.counter [1];
	assign _1013_[2] = _0876_ ^ \mchip.dut.mcp3202.counter [2];
	assign _0877_ = _0876_ & \mchip.dut.mcp3202.counter [2];
	assign _1013_[3] = _0877_ ^ \mchip.dut.mcp3202.counter [3];
	assign _0878_ = ~(\mchip.dut.mcp3202.counter [2] & \mchip.dut.mcp3202.counter [3]);
	assign _0879_ = _0876_ & ~_0878_;
	assign _1013_[4] = _0879_ ^ \mchip.dut.mcp3202.counter [4];
	assign _0880_ = \mchip.dut.p_cont.error [4] & \mchip.dut.p_setpoint_storage.p [0];
	assign _0881_ = \mchip.dut.p_cont.error [3] & \mchip.dut.p_setpoint_storage.p [1];
	assign _0882_ = ~(_0881_ & _0880_);
	assign _0883_ = ~(\mchip.dut.p_cont.error [2] & \mchip.dut.p_setpoint_storage.p [2]);
	assign _0884_ = _0881_ ^ _0880_;
	assign _0885_ = _0884_ & ~_0883_;
	assign _0886_ = _0882_ & ~_0885_;
	assign _0887_ = \mchip.dut.p_cont.error [4] & \mchip.dut.p_setpoint_storage.p [1];
	assign _0888_ = \mchip.dut.p_cont.error [5] & \mchip.dut.p_setpoint_storage.p [0];
	assign _0889_ = _0888_ ^ _0887_;
	assign _0890_ = ~(\mchip.dut.p_cont.error [3] & \mchip.dut.p_setpoint_storage.p [2]);
	assign _0891_ = _0890_ ^ _0889_;
	assign _0892_ = _0891_ | _0886_;
	assign _0893_ = ~(\mchip.dut.p_cont.error [0] & \mchip.dut.p_setpoint_storage.p [5]);
	assign _0894_ = \mchip.dut.p_cont.error [1] & \mchip.dut.p_setpoint_storage.p [4];
	assign _0895_ = ~(\mchip.dut.p_cont.error [2] & \mchip.dut.p_setpoint_storage.p [3]);
	assign _0896_ = _0895_ ^ _0894_;
	assign _0897_ = _0896_ ^ _0893_;
	assign _0898_ = ~_0897_;
	assign _0899_ = _0891_ ^ _0886_;
	assign _0900_ = _0899_ & ~_0898_;
	assign _0901_ = _0892_ & ~_0900_;
	assign _0902_ = ~(_0888_ & _0887_);
	assign _0903_ = _0889_ & ~_0890_;
	assign _0904_ = _0902_ & ~_0903_;
	assign _0905_ = \mchip.dut.p_cont.error [5] & \mchip.dut.p_setpoint_storage.p [1];
	assign _0906_ = \mchip.dut.p_cont.error [6] & \mchip.dut.p_setpoint_storage.p [0];
	assign _0907_ = _0906_ ^ _0905_;
	assign _0908_ = ~(\mchip.dut.p_cont.error [4] & \mchip.dut.p_setpoint_storage.p [2]);
	assign _0909_ = _0908_ ^ _0907_;
	assign _0910_ = _0909_ ^ _0904_;
	assign _0911_ = \mchip.dut.p_cont.error [1] & \mchip.dut.p_setpoint_storage.p [5];
	assign _0912_ = ~(\mchip.dut.p_cont.error [2] & \mchip.dut.p_setpoint_storage.p [4]);
	assign _0913_ = ~(\mchip.dut.p_cont.error [3] & \mchip.dut.p_setpoint_storage.p [3]);
	assign _0914_ = ~(_0913_ ^ _0912_);
	assign _0915_ = _0914_ ^ _0911_;
	assign _0916_ = _0915_ ^ _0910_;
	assign _0917_ = _0916_ | _0901_;
	assign _0918_ = \mchip.dut.p_cont.error [0] & \mchip.dut.p_setpoint_storage.p [6];
	assign _0919_ = ~_0918_;
	assign _0920_ = _0896_ | _0893_;
	assign _0921_ = _0894_ & ~_0895_;
	assign _0922_ = _0920_ & ~_0921_;
	assign _0923_ = _0922_ ^ _0919_;
	assign _0924_ = _0916_ ^ _0901_;
	assign _0925_ = _0924_ & _0923_;
	assign _0926_ = _0925_ | ~_0917_;
	assign _0927_ = _0909_ | _0904_;
	assign _0928_ = _0910_ & ~_0915_;
	assign _0929_ = _0927_ & ~_0928_;
	assign _0930_ = ~(_0906_ & _0905_);
	assign _0931_ = _0907_ & ~_0908_;
	assign _0932_ = _0930_ & ~_0931_;
	assign _0933_ = \mchip.dut.p_cont.error [6] & \mchip.dut.p_setpoint_storage.p [1];
	assign _0934_ = \mchip.dut.p_cont.error [7] & \mchip.dut.p_setpoint_storage.p [0];
	assign _0935_ = _0934_ ^ _0933_;
	assign _0936_ = ~(\mchip.dut.p_cont.error [5] & \mchip.dut.p_setpoint_storage.p [2]);
	assign _0937_ = _0936_ ^ _0935_;
	assign _0938_ = _0937_ ^ _0932_;
	assign _0939_ = ~(\mchip.dut.p_cont.error [2] & \mchip.dut.p_setpoint_storage.p [5]);
	assign _0940_ = \mchip.dut.p_cont.error [3] & \mchip.dut.p_setpoint_storage.p [4];
	assign _0941_ = ~(\mchip.dut.p_cont.error [4] & \mchip.dut.p_setpoint_storage.p [3]);
	assign _0942_ = _0941_ ^ _0940_;
	assign _0943_ = ~(_0942_ ^ _0939_);
	assign _0944_ = _0943_ ^ _0938_;
	assign _0945_ = _0944_ ^ _0929_;
	assign _0946_ = \mchip.dut.p_cont.error [0] & \mchip.dut.p_setpoint_storage.p [7];
	assign _0947_ = \mchip.dut.p_cont.error [1] & \mchip.dut.p_setpoint_storage.p [6];
	assign _0948_ = _0947_ ^ _0946_;
	assign _0949_ = _0913_ | _0912_;
	assign _0950_ = _0911_ & ~_0914_;
	assign _0951_ = _0949_ & ~_0950_;
	assign _0952_ = _0951_ ^ _0948_;
	assign _0953_ = _0952_ ^ _0945_;
	assign _0954_ = _0926_ & ~_0953_;
	assign _0955_ = _0918_ & ~_0922_;
	assign _0956_ = ~_0955_;
	assign _0957_ = ~(_0953_ ^ _0926_);
	assign _0958_ = _0957_ & ~_0956_;
	assign _0959_ = _0958_ | _0954_;
	assign _0960_ = _0944_ | _0929_;
	assign _0961_ = _0945_ & ~_0952_;
	assign _0962_ = _0960_ & ~_0961_;
	assign _0963_ = _0937_ | _0932_;
	assign _0964_ = _0938_ & ~_0943_;
	assign _0965_ = _0963_ & ~_0964_;
	assign _0966_ = ~(_0934_ & _0933_);
	assign _0967_ = _0935_ & ~_0936_;
	assign _0968_ = _0966_ & ~_0967_;
	assign _0969_ = ~(\mchip.dut.p_cont.error [7] & \mchip.dut.p_setpoint_storage.p [1]);
	assign _0970_ = ~(\mchip.dut.p_cont.error [8] & \mchip.dut.p_setpoint_storage.p [0]);
	assign _0971_ = _0970_ ^ _0969_;
	assign _0972_ = ~(\mchip.dut.p_cont.error [6] & \mchip.dut.p_setpoint_storage.p [2]);
	assign _0973_ = _0972_ ^ _0971_;
	assign _0974_ = _0973_ ^ _0968_;
	assign _0975_ = \mchip.dut.p_cont.error [3] & \mchip.dut.p_setpoint_storage.p [5];
	assign _0976_ = ~(\mchip.dut.p_cont.error [4] & \mchip.dut.p_setpoint_storage.p [4]);
	assign _0977_ = ~(\mchip.dut.p_cont.error [5] & \mchip.dut.p_setpoint_storage.p [3]);
	assign _0978_ = ~(_0977_ ^ _0976_);
	assign _0979_ = _0978_ ^ _0975_;
	assign _0980_ = _0979_ ^ _0974_;
	assign _0981_ = _0980_ ^ _0965_;
	assign _0982_ = _0947_ & _0946_;
	assign _0983_ = \mchip.dut.p_cont.error [1] & \mchip.dut.p_setpoint_storage.p [7];
	assign _0984_ = \mchip.dut.p_cont.error [2] & \mchip.dut.p_setpoint_storage.p [6];
	assign _0985_ = _0984_ ^ _0983_;
	assign _0986_ = _0942_ | _0939_;
	assign _0987_ = _0940_ & ~_0941_;
	assign _0988_ = _0986_ & ~_0987_;
	assign _0989_ = _0988_ ^ _0985_;
	assign _0990_ = _0989_ ^ _0982_;
	assign _0991_ = _0990_ ^ _0981_;
	assign _0992_ = _0991_ ^ _0962_;
	assign _0993_ = _0948_ & ~_0951_;
	assign _0994_ = ~_0993_;
	assign _0995_ = _0994_ ^ _0992_;
	assign _0996_ = _0995_ ^ _0959_;
	assign _0997_ = _0991_ | _0962_;
	assign _0998_ = _0992_ & ~_0994_;
	assign _0999_ = _0998_ | ~_0997_;
	assign _1000_ = _0980_ | _0965_;
	assign _1001_ = _0981_ & ~_0990_;
	assign _1002_ = _1000_ & ~_1001_;
	assign _1003_ = _0973_ | _0968_;
	assign _0076_ = _0974_ & ~_0979_;
	assign _0077_ = _1003_ & ~_0076_;
	assign _0078_ = _0970_ | _0969_;
	assign _0079_ = _0971_ & ~_0972_;
	assign _0080_ = _0078_ & ~_0079_;
	assign _0081_ = \mchip.dut.p_cont.error [7] & \mchip.dut.p_setpoint_storage.p [2];
	assign _0082_ = \mchip.dut.p_setpoint_storage.p [1] & \mchip.dut.p_cont.error [8];
	assign _0083_ = _0082_ ^ _0970_;
	assign _0084_ = _0083_ ^ _0081_;
	assign _0085_ = _0084_ ^ _0080_;
	assign _0086_ = \mchip.dut.p_cont.error [4] & \mchip.dut.p_setpoint_storage.p [5];
	assign _0087_ = ~(\mchip.dut.p_cont.error [5] & \mchip.dut.p_setpoint_storage.p [4]);
	assign _0088_ = ~(\mchip.dut.p_cont.error [6] & \mchip.dut.p_setpoint_storage.p [3]);
	assign _0089_ = ~(_0088_ ^ _0087_);
	assign _0090_ = _0089_ ^ _0086_;
	assign _0091_ = _0090_ ^ _0085_;
	assign _0092_ = _0091_ ^ _0077_;
	assign _0093_ = _0984_ & _0983_;
	assign _0094_ = \mchip.dut.p_cont.error [2] & \mchip.dut.p_setpoint_storage.p [7];
	assign _0095_ = \mchip.dut.p_cont.error [3] & \mchip.dut.p_setpoint_storage.p [6];
	assign _0096_ = _0095_ ^ _0094_;
	assign _0097_ = _0977_ | _0976_;
	assign _0098_ = _0975_ & ~_0978_;
	assign _0099_ = _0097_ & ~_0098_;
	assign _0100_ = _0099_ ^ _0096_;
	assign _0101_ = _0100_ ^ _0093_;
	assign _0102_ = _0101_ ^ _0092_;
	assign _0103_ = _0102_ ^ _1002_;
	assign _0104_ = _0989_ | ~_0982_;
	assign _0105_ = _0985_ & ~_0988_;
	assign _0106_ = _0104_ & ~_0105_;
	assign _0107_ = _0106_ ^ _0103_;
	assign _0108_ = _0107_ ^ _0999_;
	assign _0109_ = _0108_ | _0996_;
	assign _0110_ = _0924_ ^ _0923_;
	assign _0111_ = ~(\mchip.dut.p_cont.error [3] & \mchip.dut.p_setpoint_storage.p [0]);
	assign _0112_ = \mchip.dut.p_cont.error [2] & \mchip.dut.p_setpoint_storage.p [1];
	assign _0113_ = _0111_ | ~_0112_;
	assign _0114_ = \mchip.dut.p_cont.error [1] & \mchip.dut.p_setpoint_storage.p [2];
	assign _0115_ = _0112_ ^ _0111_;
	assign _0116_ = _0114_ & ~_0115_;
	assign _0117_ = _0113_ & ~_0116_;
	assign _0118_ = _0884_ ^ _0883_;
	assign _0119_ = _0118_ | _0117_;
	assign _0120_ = \mchip.dut.p_cont.error [0] & \mchip.dut.p_setpoint_storage.p [4];
	assign _0121_ = \mchip.dut.p_cont.error [1] & \mchip.dut.p_setpoint_storage.p [3];
	assign _0122_ = _0121_ ^ _0120_;
	assign _0123_ = _0118_ ^ _0117_;
	assign _0124_ = _0123_ & _0122_;
	assign _0125_ = _0119_ & ~_0124_;
	assign _0126_ = _0899_ ^ _0898_;
	assign _0127_ = _0126_ | _0125_;
	assign _0128_ = _0121_ & _0120_;
	assign _0129_ = _0126_ ^ _0125_;
	assign _0130_ = _0129_ & _0128_;
	assign _0131_ = _0127_ & ~_0130_;
	assign _0132_ = _0110_ & ~_0131_;
	assign _0133_ = _0957_ ^ _0956_;
	assign _0134_ = ~(_0133_ ^ _0132_);
	assign _0135_ = ~(\mchip.dut.p_cont.error [2] & \mchip.dut.p_setpoint_storage.p [0]);
	assign _0136_ = \mchip.dut.p_cont.error [1] & \mchip.dut.p_setpoint_storage.p [1];
	assign _0137_ = _0136_ & ~_0135_;
	assign _0138_ = \mchip.dut.p_cont.error [0] & \mchip.dut.p_setpoint_storage.p [2];
	assign _0139_ = _0136_ ^ _0135_;
	assign _0140_ = _0138_ & ~_0139_;
	assign _0141_ = ~(_0140_ | _0137_);
	assign _0142_ = ~(_0115_ ^ _0114_);
	assign _0143_ = _0141_ | ~_0142_;
	assign _0144_ = \mchip.dut.p_cont.error [0] & \mchip.dut.p_setpoint_storage.p [3];
	assign _0145_ = _0142_ ^ _0141_;
	assign _0146_ = _0144_ & ~_0145_;
	assign _0147_ = _0143_ & ~_0146_;
	assign _0148_ = _0123_ ^ _0122_;
	assign _0149_ = _0147_ | ~_0148_;
	assign _0150_ = _0129_ ^ _0128_;
	assign _0151_ = _0149_ | ~_0150_;
	assign _0152_ = ~(_0131_ ^ _0110_);
	assign _0153_ = _0152_ ^ _0151_;
	assign _0154_ = _0134_ & ~_0153_;
	assign _0155_ = ~(\mchip.dut.p_cont.error [0] & \mchip.dut.p_setpoint_storage.p [1]);
	assign _0156_ = ~(\mchip.dut.p_cont.error [1] & \mchip.dut.p_setpoint_storage.p [0]);
	assign _0157_ = _0156_ | _0155_;
	assign _0158_ = _0139_ ^ _0138_;
	assign _0159_ = _0158_ | _0157_;
	assign _0160_ = _0145_ ^ _0144_;
	assign _0161_ = _0160_ | _0159_;
	assign _0162_ = _0148_ ^ _0147_;
	assign _0163_ = _0162_ | _0161_;
	assign _0164_ = _0150_ ^ _0149_;
	assign _0165_ = _0164_ | _0163_;
	assign _0166_ = _0154_ & ~_0165_;
	assign _0167_ = _0151_ | ~_0152_;
	assign _0168_ = _0134_ & ~_0167_;
	assign _0169_ = _0132_ & ~_0133_;
	assign _0170_ = _0169_ | _0168_;
	assign _0171_ = _0170_ | _0166_;
	assign _0172_ = _0171_ & ~_0109_;
	assign _0173_ = _0959_ & ~_0995_;
	assign _0174_ = _0173_ & ~_0108_;
	assign _0175_ = _0999_ & ~_0107_;
	assign _0176_ = _0175_ | _0174_;
	assign _0177_ = _0176_ | _0172_;
	assign _0178_ = ~(_0102_ | _1002_);
	assign _0179_ = _0103_ & ~_0106_;
	assign _0180_ = _0179_ | _0178_;
	assign _0181_ = _0096_ & ~_0099_;
	assign _0182_ = _0093_ & ~_0100_;
	assign _0183_ = ~(_0182_ | _0181_);
	assign _0184_ = _0091_ | _0077_;
	assign _0185_ = _0092_ & ~_0101_;
	assign _0186_ = _0185_ | ~_0184_;
	assign _0187_ = _0095_ & _0094_;
	assign _0188_ = \mchip.dut.p_cont.error [3] & \mchip.dut.p_setpoint_storage.p [7];
	assign _0189_ = \mchip.dut.p_setpoint_storage.p [6] & \mchip.dut.p_cont.error [4];
	assign _0190_ = _0189_ ^ _0188_;
	assign _0191_ = _0088_ | _0087_;
	assign _0192_ = _0086_ & ~_0089_;
	assign _0193_ = _0191_ & ~_0192_;
	assign _0194_ = ~(_0193_ ^ _0190_);
	assign _0195_ = ~(_0194_ ^ _0187_);
	assign _0196_ = _0084_ | _0080_;
	assign _0197_ = _0085_ & ~_0090_;
	assign _0198_ = _0197_ | ~_0196_;
	assign _0199_ = ~(\mchip.dut.p_cont.error [5] & \mchip.dut.p_setpoint_storage.p [5]);
	assign _0200_ = \mchip.dut.p_cont.error [6] & \mchip.dut.p_setpoint_storage.p [4];
	assign _0201_ = ~(\mchip.dut.p_setpoint_storage.p [3] & \mchip.dut.p_cont.error [7]);
	assign _0202_ = _0201_ ^ _0200_;
	assign _0203_ = _0202_ ^ _0199_;
	assign _0204_ = _0970_ | ~_0082_;
	assign _0205_ = _0081_ & ~_0083_;
	assign _0206_ = _0205_ | ~_0204_;
	assign _0207_ = \mchip.dut.p_setpoint_storage.p [2] & \mchip.dut.p_cont.error [8];
	assign _0208_ = ~(_0207_ ^ _0083_);
	assign _0209_ = ~_0208_;
	assign _0210_ = _0209_ ^ _0206_;
	assign _0211_ = _0210_ ^ _0203_;
	assign _0212_ = _0211_ ^ _0198_;
	assign _0213_ = ~(_0212_ ^ _0195_);
	assign _0214_ = _0213_ ^ _0186_;
	assign _0215_ = _0214_ ^ _0183_;
	assign _0216_ = ~(_0215_ ^ _0180_);
	assign _1017_[10] = ~(_0216_ ^ _0177_);
	assign _0217_ = _0215_ & _0180_;
	assign _0218_ = _0177_ & ~_0216_;
	assign _0219_ = ~(_0218_ | _0217_);
	assign _0220_ = ~(_0214_ | _0183_);
	assign _0221_ = _0186_ & ~_0213_;
	assign _0222_ = _0221_ | _0220_;
	assign _0223_ = _0190_ & ~_0193_;
	assign _0224_ = _0194_ & _0187_;
	assign _0225_ = _0224_ | _0223_;
	assign _0226_ = _0212_ | _0195_;
	assign _0227_ = _0198_ & ~_0211_;
	assign _0228_ = _0226_ & ~_0227_;
	assign _0229_ = _0189_ & _0188_;
	assign _0230_ = \mchip.dut.p_setpoint_storage.p [7] & \mchip.dut.p_cont.error [4];
	assign _0231_ = \mchip.dut.p_setpoint_storage.p [6] & \mchip.dut.p_cont.error [5];
	assign _0232_ = _0231_ ^ _0230_;
	assign _0233_ = _0202_ | _0199_;
	assign _0234_ = _0200_ & ~_0201_;
	assign _0235_ = _0233_ & ~_0234_;
	assign _0236_ = ~(_0235_ ^ _0232_);
	assign _0237_ = _0236_ ^ _0229_;
	assign _0238_ = _0210_ | ~_0203_;
	assign _0239_ = _0206_ & ~_0209_;
	assign _0240_ = _0239_ | ~_0238_;
	assign _0241_ = ~(\mchip.dut.p_setpoint_storage.p [5] & \mchip.dut.p_cont.error [6]);
	assign _0242_ = ~(\mchip.dut.p_setpoint_storage.p [4] & \mchip.dut.p_cont.error [7]);
	assign _0243_ = \mchip.dut.p_setpoint_storage.p [3] & \mchip.dut.p_cont.error [8];
	assign _0244_ = _0243_ ^ _0242_;
	assign _0245_ = ~(_0244_ ^ _0241_);
	assign _0246_ = _0207_ & ~_0083_;
	assign _0247_ = _0204_ & ~_0246_;
	assign _0248_ = _0247_ ^ _0208_;
	assign _0249_ = ~(_0248_ ^ _0245_);
	assign _0250_ = _0249_ ^ _0240_;
	assign _0251_ = _0250_ ^ _0237_;
	assign _0252_ = ~(_0251_ ^ _0228_);
	assign _0253_ = _0252_ ^ _0225_;
	assign _0254_ = _0253_ ^ _0222_;
	assign _1017_[11] = _0254_ ^ _0219_;
	assign _0255_ = _0254_ | _0216_;
	assign _0256_ = _0255_ | _0109_;
	assign _0257_ = _0171_ & ~_0256_;
	assign _0258_ = _0176_ & ~_0255_;
	assign _0259_ = _0222_ & ~_0253_;
	assign _0260_ = _0217_ & ~_0254_;
	assign _0261_ = _0260_ | _0259_;
	assign _0262_ = _0261_ | _0258_;
	assign _0263_ = _0262_ | _0257_;
	assign _0264_ = ~(_0251_ | _0228_);
	assign _0265_ = _0225_ & ~_0252_;
	assign _0266_ = _0265_ | _0264_;
	assign _0267_ = _0232_ & ~_0235_;
	assign _0268_ = _0236_ & _0229_;
	assign _0269_ = ~(_0268_ | _0267_);
	assign _0270_ = _0250_ | ~_0237_;
	assign _0271_ = _0240_ & ~_0249_;
	assign _0272_ = _0271_ | ~_0270_;
	assign _0273_ = _0231_ & _0230_;
	assign _0274_ = \mchip.dut.p_setpoint_storage.p [7] & \mchip.dut.p_cont.error [5];
	assign _0275_ = \mchip.dut.p_setpoint_storage.p [6] & \mchip.dut.p_cont.error [6];
	assign _0276_ = _0275_ ^ _0274_;
	assign _0277_ = _0244_ | _0241_;
	assign _0278_ = _0243_ & ~_0242_;
	assign _0279_ = _0277_ & ~_0278_;
	assign _0280_ = ~(_0279_ ^ _0276_);
	assign _0281_ = ~(_0280_ ^ _0273_);
	assign _0282_ = _0248_ | _0245_;
	assign _0283_ = _0208_ & ~_0247_;
	assign _0284_ = ~_0283_;
	assign _0285_ = ~(_0284_ & _0282_);
	assign _0286_ = \mchip.dut.p_setpoint_storage.p [5] & \mchip.dut.p_cont.error [7];
	assign _0287_ = \mchip.dut.p_setpoint_storage.p [4] & \mchip.dut.p_cont.error [8];
	assign _0288_ = _0287_ ^ _0243_;
	assign _0289_ = _0288_ ^ _0286_;
	assign _0290_ = _0289_ ^ _0248_;
	assign _0291_ = _0290_ ^ _0285_;
	assign _0292_ = ~(_0291_ ^ _0281_);
	assign _0293_ = _0292_ ^ _0272_;
	assign _0294_ = _0293_ ^ _0269_;
	assign _0295_ = ~(_0294_ ^ _0266_);
	assign _1017_[12] = ~(_0295_ ^ _0263_);
	assign _0296_ = _0294_ & _0266_;
	assign _0297_ = _0263_ & ~_0295_;
	assign _0298_ = ~(_0297_ | _0296_);
	assign _0299_ = ~(_0293_ | _0269_);
	assign _0300_ = _0272_ & ~_0292_;
	assign _0301_ = _0300_ | _0299_;
	assign _0302_ = _0276_ & ~_0279_;
	assign _0303_ = _0280_ & _0273_;
	assign _0304_ = _0303_ | _0302_;
	assign _0305_ = _0291_ | _0281_;
	assign _0306_ = _0285_ & ~_0290_;
	assign _0307_ = _0306_ | ~_0305_;
	assign _0308_ = _0275_ & _0274_;
	assign _0309_ = \mchip.dut.p_setpoint_storage.p [7] & \mchip.dut.p_cont.error [6];
	assign _0310_ = \mchip.dut.p_setpoint_storage.p [6] & \mchip.dut.p_cont.error [7];
	assign _0311_ = _0310_ ^ _0309_;
	assign _0312_ = ~(_0287_ & _0243_);
	assign _0313_ = _0288_ & _0286_;
	assign _0314_ = _0312_ & ~_0313_;
	assign _0315_ = ~(_0314_ ^ _0311_);
	assign _0316_ = ~(_0315_ ^ _0308_);
	assign _0317_ = _0289_ & ~_0248_;
	assign _0318_ = _0317_ | _0283_;
	assign _0319_ = \mchip.dut.p_setpoint_storage.p [5] & \mchip.dut.p_cont.error [8];
	assign _0320_ = _0319_ ^ _0288_;
	assign _0321_ = ~(_0320_ ^ _0248_);
	assign _0322_ = ~_0321_;
	assign _0323_ = _0322_ ^ _0318_;
	assign _0324_ = ~(_0323_ ^ _0316_);
	assign _0325_ = _0324_ ^ _0307_;
	assign _0326_ = _0325_ ^ _0304_;
	assign _0327_ = _0326_ ^ _0301_;
	assign _1017_[13] = _0327_ ^ _0298_;
	assign _0328_ = _0327_ | _0295_;
	assign _0329_ = _0263_ & ~_0328_;
	assign _0330_ = _0301_ & ~_0326_;
	assign _0331_ = _0296_ & ~_0327_;
	assign _0332_ = _0331_ | _0330_;
	assign _0333_ = _0332_ | _0329_;
	assign _0334_ = _0307_ & ~_0324_;
	assign _0335_ = _0304_ & ~_0325_;
	assign _0336_ = _0335_ | _0334_;
	assign _0337_ = _0311_ & ~_0314_;
	assign _0338_ = _0315_ & _0308_;
	assign _0339_ = ~(_0338_ | _0337_);
	assign _0340_ = _0323_ | _0316_;
	assign _0341_ = _0318_ & ~_0322_;
	assign _0342_ = _0341_ | ~_0340_;
	assign _0343_ = _0310_ & _0309_;
	assign _0344_ = \mchip.dut.p_setpoint_storage.p [7] & \mchip.dut.p_cont.error [7];
	assign _0345_ = \mchip.dut.p_setpoint_storage.p [6] & \mchip.dut.p_cont.error [8];
	assign _0346_ = _0345_ ^ _0344_;
	assign _0347_ = _0319_ & _0288_;
	assign _0348_ = _0312_ & ~_0347_;
	assign _0349_ = ~(_0348_ ^ _0346_);
	assign _0350_ = _0349_ ^ _0343_;
	assign _0351_ = _0320_ & ~_0248_;
	assign _0352_ = _0284_ & ~_0351_;
	assign _0353_ = _0352_ ^ _0321_;
	assign _0354_ = _0353_ ^ _0350_;
	assign _0355_ = _0354_ ^ _0342_;
	assign _0356_ = _0355_ ^ _0339_;
	assign _0357_ = ~(_0356_ ^ _0336_);
	assign _1017_[14] = ~(_0357_ ^ _0333_);
	assign _0358_ = _0356_ & _0336_;
	assign _0359_ = _0333_ & ~_0357_;
	assign _0360_ = ~(_0359_ | _0358_);
	assign _0361_ = ~(_0355_ | _0339_);
	assign _0362_ = _0342_ & ~_0354_;
	assign _0363_ = _0362_ | _0361_;
	assign _0364_ = _0346_ & ~_0348_;
	assign _0365_ = _0349_ & _0343_;
	assign _0366_ = ~(_0365_ | _0364_);
	assign _0367_ = _0353_ | ~_0350_;
	assign _0368_ = _0321_ & ~_0352_;
	assign _0369_ = _0367_ & ~_0368_;
	assign _0370_ = _0345_ & _0344_;
	assign _0371_ = \mchip.dut.p_setpoint_storage.p [7] & \mchip.dut.p_cont.error [8];
	assign _0372_ = _0371_ ^ _0345_;
	assign _0373_ = ~(_0372_ ^ _0348_);
	assign _0374_ = _0373_ ^ _0370_;
	assign _0375_ = ~(_0374_ ^ _0353_);
	assign _0376_ = _0375_ ^ _0369_;
	assign _0377_ = _0376_ ^ _0366_;
	assign _0378_ = ~(_0377_ ^ _0363_);
	assign _1017_[15] = _0378_ ^ _0360_;
	assign _0379_ = _0377_ & _0363_;
	assign _0380_ = _0358_ & ~_0378_;
	assign _0381_ = _0380_ | _0379_;
	assign _0382_ = _0378_ | _0357_;
	assign _0383_ = _0332_ & ~_0382_;
	assign _0384_ = _0383_ | _0381_;
	assign _0385_ = _0382_ | _0328_;
	assign _0386_ = _0262_ & ~_0385_;
	assign _0387_ = _0386_ | _0384_;
	assign _0388_ = _0385_ | _0256_;
	assign _0389_ = _0171_ & ~_0388_;
	assign _0390_ = _0389_ | _0387_;
	assign _0391_ = ~(_0376_ | _0366_);
	assign _0392_ = _0375_ & ~_0369_;
	assign _0393_ = _0392_ | _0391_;
	assign _0394_ = _0372_ & ~_0348_;
	assign _0395_ = _0373_ & _0370_;
	assign _0396_ = _0395_ | _0394_;
	assign _0397_ = _0374_ & ~_0353_;
	assign _0398_ = ~(_0397_ | _0368_);
	assign _0399_ = _0371_ & _0345_;
	assign _0400_ = _0373_ ^ _0399_;
	assign _0401_ = ~(_0400_ ^ _0353_);
	assign _0402_ = ~_0401_;
	assign _0403_ = _0402_ ^ _0398_;
	assign _0404_ = _0403_ ^ _0396_;
	assign _0405_ = _0404_ ^ _0393_;
	assign _1017_[16] = _0405_ ^ _0390_;
	assign _0406_ = _0404_ & _0393_;
	assign _0407_ = _0405_ & _0390_;
	assign _0408_ = _0407_ | _0406_;
	assign _0409_ = _0402_ | _0398_;
	assign _0410_ = _0403_ & _0396_;
	assign _0411_ = _0409_ & ~_0410_;
	assign _0412_ = ~(_0373_ & _0399_);
	assign _0413_ = _0412_ & ~_0394_;
	assign _0414_ = _0353_ | ~_0400_;
	assign _0415_ = _0414_ & ~_0368_;
	assign _0416_ = _0415_ ^ _0402_;
	assign _0417_ = _0416_ ^ _0413_;
	assign _0418_ = _0417_ ^ _0411_;
	assign _1017_[17] = _0418_ ^ _0408_;
	assign \mchip.dut.input_spi_interface.mosi_buffer [0] = \mchip.dut.input_spi_interface.internal_reset_n  & _0066_;
	assign \mchip.dut.input_spi_interface.mosi_buffer [1] = \mchip.dut.input_spi_interface.internal_reset_n  & _0067_;
	assign \mchip.dut.input_spi_interface.mosi_buffer [2] = \mchip.dut.input_spi_interface.internal_reset_n  & _0068_;
	assign \mchip.dut.input_spi_interface.mosi_buffer [3] = \mchip.dut.input_spi_interface.internal_reset_n  & _0069_;
	assign \mchip.dut.input_spi_interface.mosi_buffer [4] = \mchip.dut.input_spi_interface.internal_reset_n  & _0070_;
	assign \mchip.dut.input_spi_interface.mosi_buffer [5] = \mchip.dut.input_spi_interface.internal_reset_n  & _0071_;
	assign \mchip.dut.input_spi_interface.mosi_buffer [6] = \mchip.dut.input_spi_interface.internal_reset_n  & _0072_;
	assign \mchip.dut.input_spi_interface.mosi_buffer [7] = \mchip.dut.input_spi_interface.internal_reset_n  & _0073_;
	reg \mchip.dut.mcp3202.sensor_reading_reg[3] ;
	always @(posedge io_in[12])
		if (_0028_)
			\mchip.dut.mcp3202.sensor_reading_reg[3]  <= io_in[8];
	assign \mchip.dut.mcp3202.sensor_reading [3] = \mchip.dut.mcp3202.sensor_reading_reg[3] ;
	reg \mchip.dut.mcp3202.sensor_reading_reg[4] ;
	always @(posedge io_in[12])
		if (_0029_)
			\mchip.dut.mcp3202.sensor_reading_reg[4]  <= io_in[8];
	assign \mchip.dut.mcp3202.sensor_reading [4] = \mchip.dut.mcp3202.sensor_reading_reg[4] ;
	reg \mchip.dut.mcp3202.sensor_reading_reg[5] ;
	always @(posedge io_in[12])
		if (_0030_)
			\mchip.dut.mcp3202.sensor_reading_reg[5]  <= io_in[8];
	assign \mchip.dut.mcp3202.sensor_reading [5] = \mchip.dut.mcp3202.sensor_reading_reg[5] ;
	reg \mchip.dut.mcp3202.sensor_reading_reg[6] ;
	always @(posedge io_in[12])
		if (_0031_)
			\mchip.dut.mcp3202.sensor_reading_reg[6]  <= io_in[8];
	assign \mchip.dut.mcp3202.sensor_reading [6] = \mchip.dut.mcp3202.sensor_reading_reg[6] ;
	reg \mchip.dut.mcp3202.sensor_reading_reg[7] ;
	always @(posedge io_in[12])
		if (_0032_)
			\mchip.dut.mcp3202.sensor_reading_reg[7]  <= io_in[8];
	assign \mchip.dut.mcp3202.sensor_reading [7] = \mchip.dut.mcp3202.sensor_reading_reg[7] ;
	reg \mchip.dut.mcp3202.sensor_reading_reg[8] ;
	always @(posedge io_in[12])
		if (_0021_)
			\mchip.dut.mcp3202.sensor_reading_reg[8]  <= io_in[8];
	assign \mchip.dut.mcp3202.sensor_reading [8] = \mchip.dut.mcp3202.sensor_reading_reg[8] ;
	reg _2092_;
	always @(posedge io_in[12]) _2092_ <= _0044_;
	assign _1018_[0] = _2092_;
	reg _2093_;
	always @(posedge io_in[12]) _2093_ <= _0045_;
	assign _1018_[1] = _2093_;
	reg _2094_;
	always @(posedge io_in[12]) _2094_ <= _0046_;
	assign _1018_[2] = _2094_;
	reg _2095_;
	always @(posedge io_in[12]) _2095_ <= _0047_;
	assign _1018_[3] = _2095_;
	reg _2096_;
	always @(posedge io_in[12]) _2096_ <= _0048_;
	assign _1018_[4] = _2096_;
	reg \mchip.dut.mcp3202.sensor_reading_reg[9] ;
	always @(posedge io_in[12])
		if (_0022_)
			\mchip.dut.mcp3202.sensor_reading_reg[9]  <= io_in[8];
	assign \mchip.dut.mcp3202.sensor_reading [9] = \mchip.dut.mcp3202.sensor_reading_reg[9] ;
	reg \mchip.dut.mcp3202.sensor_reading_reg[10] ;
	always @(posedge io_in[12])
		if (_0023_)
			\mchip.dut.mcp3202.sensor_reading_reg[10]  <= io_in[8];
	assign \mchip.dut.mcp3202.sensor_reading [10] = \mchip.dut.mcp3202.sensor_reading_reg[10] ;
	reg \mchip.dut.mcp3202.sensor_reading_reg[11] ;
	always @(posedge io_in[12])
		if (_0024_)
			\mchip.dut.mcp3202.sensor_reading_reg[11]  <= io_in[8];
	assign \mchip.dut.mcp3202.sensor_reading [11] = \mchip.dut.mcp3202.sensor_reading_reg[11] ;
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.dut.mcp3202.done_counter [0] <= 1'h0;
		else
			\mchip.dut.mcp3202.done_counter [0] <= _1014_[0];
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.dut.mcp3202.done_counter [1] <= 1'h0;
		else
			\mchip.dut.mcp3202.done_counter [1] <= _1015_[1];
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.dut.mcp3202.done_counter [2] <= 1'h0;
		else
			\mchip.dut.mcp3202.done_counter [2] <= _1015_[2];
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.dut.mcp3202.done_counter [3] <= 1'h0;
		else
			\mchip.dut.mcp3202.done_counter [3] <= _1015_[3];
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.dut.mcp3202.done_counter [4] <= 1'h0;
		else
			\mchip.dut.mcp3202.done_counter [4] <= _1015_[4];
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.dut.mcp3202.done_counter [5] <= 1'h0;
		else
			\mchip.dut.mcp3202.done_counter [5] <= _1015_[5];
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.dut.mcp3202.done_counter [6] <= 1'h0;
		else
			\mchip.dut.mcp3202.done_counter [6] <= _1015_[6];
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.dut.mcp3202.done_counter [7] <= 1'h0;
		else
			\mchip.dut.mcp3202.done_counter [7] <= _1015_[7];
	always @(posedge io_in[12])
		if (_0033_)
			\mchip.dut.mcp3202.done_counter [8] <= 1'h0;
		else
			\mchip.dut.mcp3202.done_counter [8] <= _1015_[8];
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [0] <= _0000_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [1] <= _0011_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [2] <= _0013_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [3] <= _0014_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [4] <= _0015_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [5] <= _0016_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [6] <= _0017_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [7] <= _0018_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [8] <= _0019_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [9] <= _0020_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [10] <= _0001_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [11] <= _0002_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [12] <= _0003_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [13] <= _0004_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [14] <= _0005_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [15] <= _0006_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [16] <= _0007_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [17] <= _0008_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [18] <= _0009_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [19] <= _0010_;
	always @(posedge io_in[12]) \mchip.dut.mcp3202.state [20] <= _0012_;
	always @(posedge io_in[12]) \mchip.dut.p_cont.round_reading [0] <= _0052_;
	always @(posedge io_in[12]) \mchip.dut.p_cont.round_reading [1] <= _0053_;
	always @(posedge io_in[12]) \mchip.dut.p_cont.round_reading [2] <= _0054_;
	always @(posedge io_in[12]) \mchip.dut.p_cont.round_reading [3] <= _0055_;
	always @(posedge io_in[12]) \mchip.dut.p_cont.round_reading [4] <= _0056_;
	always @(posedge io_in[12]) \mchip.dut.p_cont.round_reading [5] <= _0057_;
	always @(posedge io_in[12]) \mchip.dut.p_cont.round_reading [6] <= _0058_;
	always @(posedge io_in[12]) \mchip.dut.p_cont.round_reading [7] <= _0059_;
	always @(posedge io_in[12])
		if (!_0040_)
			\mchip.dut.input_spi_interface.cs_n.data_out  <= 1'h1;
		else if (!_0037_)
			\mchip.dut.input_spi_interface.cs_n.data_out  <= 1'h0;
	always @(posedge io_in[12]) \mchip.dut.input_spi_interface.cs_n.data_buffer [0] <= io_in[9];
	always @(posedge io_in[12]) \mchip.dut.input_spi_interface.cs_n.data_buffer [1] <= \mchip.dut.input_spi_interface.cs_n.data_buffer [0];
	always @(posedge io_in[12]) \mchip.dut.input_spi_interface.cs_n.data_buffer [2] <= \mchip.dut.input_spi_interface.cs_n.data_buffer [1];
	always @(posedge io_in[12])
		if (!_0041_)
			\mchip.dut.input_spi_interface.mosi.data_out  <= 1'h1;
		else if (!_0038_)
			\mchip.dut.input_spi_interface.mosi.data_out  <= 1'h0;
	always @(posedge io_in[12]) \mchip.dut.input_spi_interface.mosi.data_buffer [0] <= io_in[10];
	always @(posedge io_in[12]) \mchip.dut.input_spi_interface.mosi.data_buffer [1] <= \mchip.dut.input_spi_interface.mosi.data_buffer [0];
	always @(posedge io_in[12]) \mchip.dut.input_spi_interface.mosi.data_buffer [2] <= \mchip.dut.input_spi_interface.mosi.data_buffer [1];
	always @(posedge io_in[12])
		if (!_0042_)
			\mchip.dut.input_spi_interface.clk.data_out  <= 1'h1;
		else if (!_0039_)
			\mchip.dut.input_spi_interface.clk.data_out  <= 1'h0;
	always @(posedge io_in[12]) \mchip.dut.input_spi_interface.clk.data_buffer [0] <= io_in[11];
	always @(posedge io_in[12]) \mchip.dut.input_spi_interface.clk.data_buffer [1] <= \mchip.dut.input_spi_interface.clk.data_buffer [0];
	always @(posedge io_in[12]) \mchip.dut.input_spi_interface.clk.data_buffer [2] <= \mchip.dut.input_spi_interface.clk.data_buffer [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0060_ <= 1'h1;
		else
			_0060_ <= \mchip.dut.input_spi_interface.cs_n.data_out ;
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0061_ <= 1'h0;
		else
			_0061_ <= _1010_[0];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0062_ <= 1'h0;
		else
			_0062_ <= _1011_[1];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0063_ <= 1'h0;
		else
			_0063_ <= _1011_[2];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0064_ <= 1'h0;
		else
			_0064_ <= _1011_[3];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0065_ <= 1'h0;
		else
			_0065_ <= _1011_[4];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0066_ <= 1'h0;
		else
			_0066_ <= \mchip.dut.input_spi_interface.mosi.data_out ;
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0067_ <= 1'h0;
		else
			_0067_ <= \mchip.dut.input_spi_interface.mosi_buffer [0];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0068_ <= 1'h0;
		else
			_0068_ <= \mchip.dut.input_spi_interface.mosi_buffer [1];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0069_ <= 1'h0;
		else
			_0069_ <= \mchip.dut.input_spi_interface.mosi_buffer [2];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0070_ <= 1'h0;
		else
			_0070_ <= \mchip.dut.input_spi_interface.mosi_buffer [3];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0071_ <= 1'h0;
		else
			_0071_ <= \mchip.dut.input_spi_interface.mosi_buffer [4];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0072_ <= 1'h0;
		else
			_0072_ <= \mchip.dut.input_spi_interface.mosi_buffer [5];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0073_ <= 1'h0;
		else
			_0073_ <= \mchip.dut.input_spi_interface.mosi_buffer [6];
	always @(posedge \mchip.dut.input_spi_interface.clk.data_out )
		if (!\mchip.dut.input_spi_interface.internal_reset_n )
			_0074_ <= 1'h0;
		else
			_0074_ <= \mchip.dut.input_spi_interface.mosi_buffer [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0075_ <= 1'h0;
		else
			_0075_ <= _0049_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.setpoint [0] <= 1'h1;
		else if (_0026_)
			\mchip.dut.p_setpoint_storage.setpoint [0] <= \mchip.dut.input_spi_interface.mosi_buffer [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.setpoint [1] <= 1'h1;
		else if (_0026_)
			\mchip.dut.p_setpoint_storage.setpoint [1] <= \mchip.dut.input_spi_interface.mosi_buffer [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.setpoint [2] <= 1'h1;
		else if (_0026_)
			\mchip.dut.p_setpoint_storage.setpoint [2] <= \mchip.dut.input_spi_interface.mosi_buffer [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.setpoint [3] <= 1'h1;
		else if (_0026_)
			\mchip.dut.p_setpoint_storage.setpoint [3] <= \mchip.dut.input_spi_interface.mosi_buffer [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.setpoint [4] <= 1'h1;
		else if (_0026_)
			\mchip.dut.p_setpoint_storage.setpoint [4] <= \mchip.dut.input_spi_interface.mosi_buffer [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.setpoint [5] <= 1'h1;
		else if (_0026_)
			\mchip.dut.p_setpoint_storage.setpoint [5] <= \mchip.dut.input_spi_interface.mosi_buffer [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.setpoint [6] <= 1'h1;
		else if (_0026_)
			\mchip.dut.p_setpoint_storage.setpoint [6] <= \mchip.dut.input_spi_interface.mosi_buffer [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.setpoint [7] <= 1'h0;
		else if (_0026_)
			\mchip.dut.p_setpoint_storage.setpoint [7] <= \mchip.dut.input_spi_interface.mosi_buffer [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.p [0] <= 1'h0;
		else if (_0025_)
			\mchip.dut.p_setpoint_storage.p [0] <= \mchip.dut.input_spi_interface.mosi_buffer [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.p [1] <= 1'h0;
		else if (_0025_)
			\mchip.dut.p_setpoint_storage.p [1] <= \mchip.dut.input_spi_interface.mosi_buffer [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.p [2] <= 1'h0;
		else if (_0025_)
			\mchip.dut.p_setpoint_storage.p [2] <= \mchip.dut.input_spi_interface.mosi_buffer [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.p [3] <= 1'h0;
		else if (_0025_)
			\mchip.dut.p_setpoint_storage.p [3] <= \mchip.dut.input_spi_interface.mosi_buffer [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.p [4] <= 1'h1;
		else if (_0025_)
			\mchip.dut.p_setpoint_storage.p [4] <= \mchip.dut.input_spi_interface.mosi_buffer [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.p [5] <= 1'h0;
		else if (_0025_)
			\mchip.dut.p_setpoint_storage.p [5] <= \mchip.dut.input_spi_interface.mosi_buffer [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.p [6] <= 1'h0;
		else if (_0025_)
			\mchip.dut.p_setpoint_storage.p [6] <= \mchip.dut.input_spi_interface.mosi_buffer [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.p_setpoint_storage.p [7] <= 1'h0;
		else if (_0025_)
			\mchip.dut.p_setpoint_storage.p [7] <= \mchip.dut.input_spi_interface.mosi_buffer [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.mcp3202.counter [0] <= 1'h0;
		else
			\mchip.dut.mcp3202.counter [0] <= _1012_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.mcp3202.counter [1] <= 1'h0;
		else
			\mchip.dut.mcp3202.counter [1] <= _1013_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.mcp3202.counter [2] <= 1'h0;
		else
			\mchip.dut.mcp3202.counter [2] <= _1013_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.mcp3202.counter [3] <= 1'h0;
		else
			\mchip.dut.mcp3202.counter [3] <= _1013_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.mcp3202.counter [4] <= 1'h0;
		else
			\mchip.dut.mcp3202.counter [4] <= _1013_[4];
	always @(posedge io_in[12])
		if (_0050_)
			\mchip.dut.mcp3202.spi_clk  <= 1'h0;
		else
			\mchip.dut.mcp3202.spi_clk  <= \mchip.dut.mcp3202.counter [4];
	always @(posedge io_in[12]) \mchip.dut.mcp3202.spi_cs_n  <= _0050_;
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.dut.mcp3202.spi_mosi  <= 1'h1;
		else
			\mchip.dut.mcp3202.spi_mosi  <= _0051_;
	always @(posedge io_in[12])
		if (_0043_)
			\mchip.dut.mcp3202.reading_valid  <= 1'h0;
		else if (_0027_)
			\mchip.dut.mcp3202.reading_valid  <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [0] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [0] <= _1008_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [1] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [1] <= _1009_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [2] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [2] <= _1009_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [3] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [3] <= _1009_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [4] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [4] <= _1009_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [5] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [5] <= _1009_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [6] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [6] <= _1009_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [7] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [7] <= _1009_[7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [8] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [8] <= _1009_[8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.b.counter [9] <= 1'h0;
		else
			\mchip.dut.driver.b.counter [9] <= _1009_[9];
	reg \mchip.dut.p_cont.internal_output_setpoint_reg[10] ;
	always @(posedge io_in[12]) \mchip.dut.p_cont.internal_output_setpoint_reg[10]  <= _1017_[10];
	assign \mchip.dut.p_cont.internal_output_setpoint [10] = \mchip.dut.p_cont.internal_output_setpoint_reg[10] ;
	reg \mchip.dut.p_cont.internal_output_setpoint_reg[11] ;
	always @(posedge io_in[12]) \mchip.dut.p_cont.internal_output_setpoint_reg[11]  <= _1017_[11];
	assign \mchip.dut.p_cont.internal_output_setpoint [11] = \mchip.dut.p_cont.internal_output_setpoint_reg[11] ;
	reg \mchip.dut.p_cont.internal_output_setpoint_reg[12] ;
	always @(posedge io_in[12]) \mchip.dut.p_cont.internal_output_setpoint_reg[12]  <= _1017_[12];
	assign \mchip.dut.p_cont.internal_output_setpoint [12] = \mchip.dut.p_cont.internal_output_setpoint_reg[12] ;
	reg \mchip.dut.p_cont.internal_output_setpoint_reg[13] ;
	always @(posedge io_in[12]) \mchip.dut.p_cont.internal_output_setpoint_reg[13]  <= _1017_[13];
	assign \mchip.dut.p_cont.internal_output_setpoint [13] = \mchip.dut.p_cont.internal_output_setpoint_reg[13] ;
	reg \mchip.dut.p_cont.internal_output_setpoint_reg[14] ;
	always @(posedge io_in[12]) \mchip.dut.p_cont.internal_output_setpoint_reg[14]  <= _1017_[14];
	assign \mchip.dut.p_cont.internal_output_setpoint [14] = \mchip.dut.p_cont.internal_output_setpoint_reg[14] ;
	reg \mchip.dut.p_cont.internal_output_setpoint_reg[15] ;
	always @(posedge io_in[12]) \mchip.dut.p_cont.internal_output_setpoint_reg[15]  <= _1017_[15];
	assign \mchip.dut.p_cont.internal_output_setpoint [15] = \mchip.dut.p_cont.internal_output_setpoint_reg[15] ;
	reg \mchip.dut.p_cont.internal_output_setpoint_reg[16] ;
	always @(posedge io_in[12]) \mchip.dut.p_cont.internal_output_setpoint_reg[16]  <= _1017_[16];
	assign \mchip.dut.p_cont.internal_output_setpoint [16] = \mchip.dut.p_cont.internal_output_setpoint_reg[16] ;
	reg \mchip.dut.p_cont.internal_output_setpoint_reg[17] ;
	always @(posedge io_in[12]) \mchip.dut.p_cont.internal_output_setpoint_reg[17]  <= _1017_[17];
	assign \mchip.dut.p_cont.internal_output_setpoint [17] = \mchip.dut.p_cont.internal_output_setpoint_reg[17] ;
	always @(posedge io_in[12]) \mchip.dut.p_cont.output_setpoint [0] <= \mchip.dut.p_cont.internal_output_setpoint [10];
	always @(posedge io_in[12]) \mchip.dut.p_cont.output_setpoint [1] <= \mchip.dut.p_cont.internal_output_setpoint [11];
	always @(posedge io_in[12]) \mchip.dut.p_cont.output_setpoint [2] <= \mchip.dut.p_cont.internal_output_setpoint [12];
	always @(posedge io_in[12]) \mchip.dut.p_cont.output_setpoint [3] <= \mchip.dut.p_cont.internal_output_setpoint [13];
	always @(posedge io_in[12]) \mchip.dut.p_cont.output_setpoint [4] <= \mchip.dut.p_cont.internal_output_setpoint [14];
	always @(posedge io_in[12]) \mchip.dut.p_cont.output_setpoint [5] <= \mchip.dut.p_cont.internal_output_setpoint [15];
	always @(posedge io_in[12]) \mchip.dut.p_cont.output_setpoint [6] <= \mchip.dut.p_cont.internal_output_setpoint [16];
	always @(posedge io_in[12]) \mchip.dut.p_cont.output_setpoint [7] <= \mchip.dut.p_cont.internal_output_setpoint [17];
	always @(posedge io_in[12]) \mchip.dut.p_cont.error [0] <= _1016_[0];
	always @(posedge io_in[12]) \mchip.dut.p_cont.error [1] <= _1016_[1];
	always @(posedge io_in[12]) \mchip.dut.p_cont.error [2] <= _1016_[2];
	always @(posedge io_in[12]) \mchip.dut.p_cont.error [3] <= _1016_[3];
	always @(posedge io_in[12]) \mchip.dut.p_cont.error [4] <= _1016_[4];
	always @(posedge io_in[12]) \mchip.dut.p_cont.error [5] <= _1016_[5];
	always @(posedge io_in[12]) \mchip.dut.p_cont.error [6] <= _1016_[6];
	always @(posedge io_in[12]) \mchip.dut.p_cont.error [7] <= _1016_[7];
	always @(posedge io_in[12]) \mchip.dut.p_cont.error [8] <= _1016_[8];
	always @(posedge io_in[12]) \mchip.dut.driver.b.pwm_out  <= _0035_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [0] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [0] <= _1006_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [1] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [1] <= _1007_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [2] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [2] <= _1007_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [3] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [3] <= _1007_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [4] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [4] <= _1007_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [5] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [5] <= _1007_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [6] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [6] <= _1007_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [7] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [7] <= _1007_[7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [8] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [8] <= _1007_[8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.a.counter [9] <= 1'h0;
		else
			\mchip.dut.driver.a.counter [9] <= _1007_[9];
	always @(posedge io_in[12]) \mchip.dut.driver.a.pwm_out  <= _0036_;
	reg \mchip.dut.driver.motor_b_duty_cycle_reg[1] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_b_duty_cycle_reg[1]  <= 1'h1;
		else
			\mchip.dut.driver.motor_b_duty_cycle_reg[1]  <= _1004_[1];
	assign \mchip.dut.driver.motor_b_duty_cycle [1] = \mchip.dut.driver.motor_b_duty_cycle_reg[1] ;
	reg \mchip.dut.driver.motor_b_duty_cycle_reg[2] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_b_duty_cycle_reg[2]  <= 1'h1;
		else
			\mchip.dut.driver.motor_b_duty_cycle_reg[2]  <= _1004_[2];
	assign \mchip.dut.driver.motor_b_duty_cycle [2] = \mchip.dut.driver.motor_b_duty_cycle_reg[2] ;
	reg \mchip.dut.driver.motor_b_duty_cycle_reg[3] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_b_duty_cycle_reg[3]  <= 1'h1;
		else
			\mchip.dut.driver.motor_b_duty_cycle_reg[3]  <= _1004_[3];
	assign \mchip.dut.driver.motor_b_duty_cycle [3] = \mchip.dut.driver.motor_b_duty_cycle_reg[3] ;
	reg \mchip.dut.driver.motor_b_duty_cycle_reg[4] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_b_duty_cycle_reg[4]  <= 1'h1;
		else
			\mchip.dut.driver.motor_b_duty_cycle_reg[4]  <= _1004_[4];
	assign \mchip.dut.driver.motor_b_duty_cycle [4] = \mchip.dut.driver.motor_b_duty_cycle_reg[4] ;
	reg \mchip.dut.driver.motor_b_duty_cycle_reg[5] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_b_duty_cycle_reg[5]  <= 1'h1;
		else
			\mchip.dut.driver.motor_b_duty_cycle_reg[5]  <= _1004_[5];
	assign \mchip.dut.driver.motor_b_duty_cycle [5] = \mchip.dut.driver.motor_b_duty_cycle_reg[5] ;
	reg \mchip.dut.driver.motor_b_duty_cycle_reg[6] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_b_duty_cycle_reg[6]  <= 1'h1;
		else
			\mchip.dut.driver.motor_b_duty_cycle_reg[6]  <= _1004_[6];
	assign \mchip.dut.driver.motor_b_duty_cycle [6] = \mchip.dut.driver.motor_b_duty_cycle_reg[6] ;
	reg \mchip.dut.driver.motor_b_duty_cycle_reg[7] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_b_duty_cycle_reg[7]  <= 1'h0;
		else
			\mchip.dut.driver.motor_b_duty_cycle_reg[7]  <= \mchip.dut.p_cont.output_setpoint [7];
	assign \mchip.dut.driver.motor_b_duty_cycle [7] = \mchip.dut.driver.motor_b_duty_cycle_reg[7] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_a_duty_cycle [0] <= 1'h1;
		else
			\mchip.dut.driver.motor_a_duty_cycle [0] <= _1004_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_a_duty_cycle [1] <= 1'h1;
		else
			\mchip.dut.driver.motor_a_duty_cycle [1] <= _1005_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_a_duty_cycle [2] <= 1'h1;
		else
			\mchip.dut.driver.motor_a_duty_cycle [2] <= _1005_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_a_duty_cycle [3] <= 1'h1;
		else
			\mchip.dut.driver.motor_a_duty_cycle [3] <= _1005_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_a_duty_cycle [4] <= 1'h1;
		else
			\mchip.dut.driver.motor_a_duty_cycle [4] <= _1005_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_a_duty_cycle [5] <= 1'h1;
		else
			\mchip.dut.driver.motor_a_duty_cycle [5] <= _1005_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_a_duty_cycle [6] <= 1'h1;
		else
			\mchip.dut.driver.motor_a_duty_cycle [6] <= _1005_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.dut.driver.motor_a_duty_cycle [7] <= 1'h0;
		else
			\mchip.dut.driver.motor_a_duty_cycle [7] <= _1005_[7];
	reg \mchip.dut.sensor_reading_captured_reg[3] ;
	always @(posedge io_in[12])
		if (\mchip.dut.mcp3202.reading_valid )
			\mchip.dut.sensor_reading_captured_reg[3]  <= \mchip.dut.mcp3202.sensor_reading [3];
	assign \mchip.dut.sensor_reading_captured [3] = \mchip.dut.sensor_reading_captured_reg[3] ;
	reg \mchip.dut.sensor_reading_captured_reg[4] ;
	always @(posedge io_in[12])
		if (\mchip.dut.mcp3202.reading_valid )
			\mchip.dut.sensor_reading_captured_reg[4]  <= \mchip.dut.mcp3202.sensor_reading [4];
	assign \mchip.dut.sensor_reading_captured [4] = \mchip.dut.sensor_reading_captured_reg[4] ;
	reg \mchip.dut.sensor_reading_captured_reg[5] ;
	always @(posedge io_in[12])
		if (\mchip.dut.mcp3202.reading_valid )
			\mchip.dut.sensor_reading_captured_reg[5]  <= \mchip.dut.mcp3202.sensor_reading [5];
	assign \mchip.dut.sensor_reading_captured [5] = \mchip.dut.sensor_reading_captured_reg[5] ;
	reg \mchip.dut.sensor_reading_captured_reg[6] ;
	always @(posedge io_in[12])
		if (\mchip.dut.mcp3202.reading_valid )
			\mchip.dut.sensor_reading_captured_reg[6]  <= \mchip.dut.mcp3202.sensor_reading [6];
	assign \mchip.dut.sensor_reading_captured [6] = \mchip.dut.sensor_reading_captured_reg[6] ;
	reg \mchip.dut.sensor_reading_captured_reg[7] ;
	always @(posedge io_in[12])
		if (\mchip.dut.mcp3202.reading_valid )
			\mchip.dut.sensor_reading_captured_reg[7]  <= \mchip.dut.mcp3202.sensor_reading [7];
	assign \mchip.dut.sensor_reading_captured [7] = \mchip.dut.sensor_reading_captured_reg[7] ;
	reg \mchip.dut.sensor_reading_captured_reg[8] ;
	always @(posedge io_in[12])
		if (\mchip.dut.mcp3202.reading_valid )
			\mchip.dut.sensor_reading_captured_reg[8]  <= \mchip.dut.mcp3202.sensor_reading [8];
	assign \mchip.dut.sensor_reading_captured [8] = \mchip.dut.sensor_reading_captured_reg[8] ;
	reg \mchip.dut.sensor_reading_captured_reg[9] ;
	always @(posedge io_in[12])
		if (\mchip.dut.mcp3202.reading_valid )
			\mchip.dut.sensor_reading_captured_reg[9]  <= \mchip.dut.mcp3202.sensor_reading [9];
	assign \mchip.dut.sensor_reading_captured [9] = \mchip.dut.sensor_reading_captured_reg[9] ;
	reg \mchip.dut.sensor_reading_captured_reg[10] ;
	always @(posedge io_in[12])
		if (\mchip.dut.mcp3202.reading_valid )
			\mchip.dut.sensor_reading_captured_reg[10]  <= \mchip.dut.mcp3202.sensor_reading [10];
	assign \mchip.dut.sensor_reading_captured [10] = \mchip.dut.sensor_reading_captured_reg[10] ;
	reg \mchip.dut.sensor_reading_captured_reg[11] ;
	always @(posedge io_in[12])
		if (\mchip.dut.mcp3202.reading_valid )
			\mchip.dut.sensor_reading_captured_reg[11]  <= \mchip.dut.mcp3202.sensor_reading [11];
	assign \mchip.dut.sensor_reading_captured [11] = \mchip.dut.sensor_reading_captured_reg[11] ;
	assign _1004_[7] = \mchip.dut.p_cont.output_setpoint [7];
	assign _1005_[0] = _1004_[0];
	assign _1006_[9:1] = \mchip.dut.driver.a.counter [9:1];
	assign _1007_[0] = _1006_[0];
	assign _1008_[9:1] = \mchip.dut.driver.b.counter [9:1];
	assign _1009_[0] = _1008_[0];
	assign _1010_[4:1] = \mchip.dut.input_spi_interface.mosi_buffer_counter [4:1];
	assign _1011_[0] = _1010_[0];
	assign _1012_[4:1] = \mchip.dut.mcp3202.counter [4:1];
	assign _1013_[0] = _1012_[0];
	assign _1014_[8:1] = \mchip.dut.mcp3202.done_counter [8:1];
	assign _1015_[0] = _1014_[0];
	assign _1017_[9:0] = 10'h000;
	assign _1018_[31:5] = 27'h0000000;
	assign io_out = {2'h0, \mchip.dut.mcp3202.spi_clk , \mchip.dut.mcp3202.spi_mosi , \mchip.dut.mcp3202.spi_cs_n , \mchip.dut.driver.a.pwm_out , \mchip.dut.driver.b.pwm_out , 7'h00};
	assign \mchip.clock  = io_in[12];
	assign \mchip.dut.adc_spi_clk  = \mchip.dut.mcp3202.spi_clk ;
	assign \mchip.dut.adc_spi_cs_n  = \mchip.dut.mcp3202.spi_cs_n ;
	assign \mchip.dut.adc_spi_miso  = io_in[8];
	assign \mchip.dut.adc_spi_mosi  = \mchip.dut.mcp3202.spi_mosi ;
	assign \mchip.dut.clk  = io_in[12];
	assign \mchip.dut.driver.a.clk  = io_in[12];
	assign \mchip.dut.driver.a.duty_cycle  = \mchip.dut.driver.motor_a_duty_cycle ;
	assign \mchip.dut.driver.a.switch_threshold  = {\mchip.dut.driver.motor_a_duty_cycle , 2'h0};
	assign \mchip.dut.driver.b.clk  = io_in[12];
	assign \mchip.dut.driver.b.duty_cycle  = {\mchip.dut.driver.motor_b_duty_cycle [7:1], \mchip.dut.driver.motor_a_duty_cycle [0]};
	assign \mchip.dut.driver.b.switch_threshold  = {\mchip.dut.driver.motor_b_duty_cycle [7:1], \mchip.dut.driver.motor_a_duty_cycle [0], 2'h0};
	assign \mchip.dut.driver.clk  = io_in[12];
	assign \mchip.dut.driver.motor_b_duty_cycle [0] = \mchip.dut.driver.motor_a_duty_cycle [0];
	assign \mchip.dut.driver.pwm_a  = \mchip.dut.driver.a.pwm_out ;
	assign \mchip.dut.driver.pwm_b  = \mchip.dut.driver.b.pwm_out ;
	assign \mchip.dut.driver.setpoint  = \mchip.dut.p_cont.output_setpoint ;
	assign {\mchip.dut.input_mosi_buffer [15:9], \mchip.dut.input_mosi_buffer [7:0]} = {7'h00, \mchip.dut.input_spi_interface.mosi_buffer [7:0]};
	assign \mchip.dut.input_spi_clk  = io_in[11];
	assign \mchip.dut.input_spi_cs_n  = io_in[9];
	assign \mchip.dut.input_spi_interface.clk.clk  = io_in[12];
	assign \mchip.dut.input_spi_interface.clk.data_in  = io_in[11];
	assign \mchip.dut.input_spi_interface.cs_n.clk  = io_in[12];
	assign \mchip.dut.input_spi_interface.cs_n.data_in  = io_in[9];
	assign \mchip.dut.input_spi_interface.mosi.clk  = io_in[12];
	assign \mchip.dut.input_spi_interface.mosi.data_in  = io_in[10];
	assign \mchip.dut.input_spi_interface.mosi_buffer [15:8] = {7'h00, \mchip.dut.input_mosi_buffer [8]};
	assign \mchip.dut.input_spi_interface.spi_clk  = io_in[11];
	assign \mchip.dut.input_spi_interface.spi_cs_n  = io_in[9];
	assign \mchip.dut.input_spi_interface.spi_mosi  = io_in[10];
	assign \mchip.dut.input_spi_interface.sync_spi_clk  = \mchip.dut.input_spi_interface.clk.data_out ;
	assign \mchip.dut.input_spi_interface.sync_spi_cs_n  = \mchip.dut.input_spi_interface.cs_n.data_out ;
	assign \mchip.dut.input_spi_interface.sync_spi_mosi  = \mchip.dut.input_spi_interface.mosi.data_out ;
	assign \mchip.dut.input_spi_interface.sys_clk  = io_in[12];
	assign \mchip.dut.input_spi_mosi  = io_in[10];
	assign \mchip.dut.mcp3202.next_state  = 32'd0;
	assign \mchip.dut.mcp3202.sensor_reading [2:0] = 3'h0;
	assign \mchip.dut.mcp3202.spi_miso  = io_in[8];
	assign \mchip.dut.mcp3202.sys_clk  = io_in[12];
	assign \mchip.dut.motor_setpoint  = \mchip.dut.p_cont.output_setpoint ;
	assign \mchip.dut.p  = \mchip.dut.p_setpoint_storage.p ;
	assign \mchip.dut.p_cont.clk  = io_in[12];
	assign \mchip.dut.p_cont.internal_output_setpoint [9:0] = 10'h000;
	assign \mchip.dut.p_cont.p  = \mchip.dut.p_setpoint_storage.p ;
	assign \mchip.dut.p_cont.sensor_reading  = {\mchip.dut.sensor_reading_captured [11:3], 3'h0};
	assign \mchip.dut.p_cont.setpoint  = \mchip.dut.p_setpoint_storage.setpoint ;
	assign \mchip.dut.p_setpoint_storage.address  = \mchip.dut.input_mosi_buffer [8];
	assign \mchip.dut.p_setpoint_storage.clk  = io_in[12];
	assign \mchip.dut.p_setpoint_storage.param  = \mchip.dut.input_spi_interface.mosi_buffer [7:0];
	assign \mchip.dut.param_address  = \mchip.dut.input_mosi_buffer [8];
	assign \mchip.dut.param_value  = \mchip.dut.input_spi_interface.mosi_buffer [7:0];
	assign \mchip.dut.pwm_a  = \mchip.dut.driver.a.pwm_out ;
	assign \mchip.dut.pwm_b  = \mchip.dut.driver.b.pwm_out ;
	assign \mchip.dut.sensor_reading  = {\mchip.dut.mcp3202.sensor_reading [11:3], 3'h0};
	assign \mchip.dut.sensor_reading_captured [2:0] = 3'h0;
	assign \mchip.dut.sensor_reading_valid  = \mchip.dut.mcp3202.reading_valid ;
	assign \mchip.dut.setpoint  = \mchip.dut.p_setpoint_storage.setpoint ;
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.dut.mcp3202.spi_clk , \mchip.dut.mcp3202.spi_mosi , \mchip.dut.mcp3202.spi_cs_n , \mchip.dut.driver.a.pwm_out , \mchip.dut.driver.b.pwm_out , 7'h00};
	assign \mchip.reset  = io_in[13];
endmodule
module d19_gsavant_16bit_serial_cpu (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire _2025_;
	wire _2026_;
	wire _2027_;
	wire [4:0] _2028_;
	wire [4:0] _2029_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [15:0] \mchip.cpu.alu.result ;
	wire [15:0] \mchip.cpu.alu_result ;
	wire \mchip.cpu.ard_clk ;
	wire \mchip.cpu.ard_data_ready ;
	wire \mchip.cpu.ard_receive_ready ;
	wire \mchip.cpu.bus_mar ;
	wire \mchip.cpu.bus_mdr ;
	wire \mchip.cpu.bus_pc ;
	wire \mchip.cpu.clk ;
	wire [9:0] \mchip.cpu.ctrl ;
	wire \mchip.cpu.ctrl_fsm.ard_data_ready ;
	wire \mchip.cpu.ctrl_fsm.ard_receive_ready ;
	wire \mchip.cpu.ctrl_fsm.bus_mar ;
	wire \mchip.cpu.ctrl_fsm.bus_mdr ;
	wire \mchip.cpu.ctrl_fsm.bus_pc ;
	wire \mchip.cpu.ctrl_fsm.clk ;
	wire [14:0] \mchip.cpu.ctrl_fsm.cs ;
	wire [9:0] \mchip.cpu.ctrl_fsm.ctrl ;
	wire \mchip.cpu.ctrl_fsm.halt ;
	wire \mchip.cpu.ctrl_fsm.rst ;
	wire [43:0] \mchip.cpu.ctrl_fsm.signals ;
	wire [43:0] \mchip.cpu.dec ;
	wire [15:0] \mchip.cpu.dec_instr.instruction ;
	wire [43:0] \mchip.cpu.dec_instr.signals ;
	wire \mchip.cpu.error_instr ;
	wire \mchip.cpu.halt ;
	wire [15:0] \mchip.cpu.imm ;
	wire [7:0] \mchip.cpu.in_bus ;
	wire [15:0] \mchip.cpu.instr ;
	wire \mchip.cpu.instr_shift.clk ;
	reg [4:0] \mchip.cpu.instr_shift.count ;
	wire \mchip.cpu.instr_shift.data_ready ;
	wire \mchip.cpu.instr_shift.error ;
	wire \mchip.cpu.instr_shift.halt ;
	reg [15:0] \mchip.cpu.instr_shift.imm ;
	reg [15:0] \mchip.cpu.instr_shift.instruction ;
	wire [2:0] \mchip.cpu.instr_shift.opcode ;
	wire \mchip.cpu.instr_shift.rst ;
	wire [7:0] \mchip.cpu.instr_shift.serial_in ;
	wire [15:0] \mchip.cpu.mar_in ;
	wire [15:0] \mchip.cpu.mar_out ;
	wire \mchip.cpu.mar_shift_reg.clk ;
	wire \mchip.cpu.mar_shift_reg.load ;
	reg \mchip.cpu.mar_shift_reg.low_b ;
	wire [15:0] \mchip.cpu.mar_shift_reg.prll_in ;
	reg [15:0] \mchip.cpu.mar_shift_reg.prll_out ;
	wire \mchip.cpu.mar_shift_reg.rst ;
	wire [7:0] \mchip.cpu.mar_shift_reg.serial_in ;
	wire \mchip.cpu.mar_shift_reg.shift_in ;
	wire \mchip.cpu.mar_shift_reg.shift_out ;
	wire [15:0] \mchip.cpu.mdr_out ;
	wire \mchip.cpu.mdr_shift_reg.clk ;
	wire \mchip.cpu.mdr_shift_reg.load ;
	reg \mchip.cpu.mdr_shift_reg.low_b ;
	reg [15:0] \mchip.cpu.mdr_shift_reg.prll_out ;
	wire \mchip.cpu.mdr_shift_reg.rst ;
	wire [7:0] \mchip.cpu.mdr_shift_reg.serial_in ;
	wire \mchip.cpu.mdr_shift_reg.shift_in ;
	wire \mchip.cpu.mdr_shift_reg.shift_out ;
	wire [7:0] \mchip.cpu.out_bus ;
	wire [15:0] \mchip.cpu.pc ;
	wire [15:0] \mchip.cpu.pc_in ;
	wire \mchip.cpu.pc_reg.clk ;
	wire \mchip.cpu.pc_reg.load ;
	reg \mchip.cpu.pc_reg.low_b ;
	wire [15:0] \mchip.cpu.pc_reg.prll_in ;
	reg [15:0] \mchip.cpu.pc_reg.prll_out ;
	wire \mchip.cpu.pc_reg.rst ;
	wire \mchip.cpu.pc_reg.shift_out ;
	wire [15:0] \mchip.cpu.rd_data ;
	wire \mchip.cpu.rf.clk ;
	wire [2:0] \mchip.cpu.rf.rd ;
	wire [15:0] \mchip.cpu.rf.rd_data ;
	reg [15:0] \mchip.cpu.rf.reg_file[0] ;
	reg [15:0] \mchip.cpu.rf.reg_file[1] ;
	reg [15:0] \mchip.cpu.rf.reg_file[2] ;
	reg [15:0] \mchip.cpu.rf.reg_file[3] ;
	reg [15:0] \mchip.cpu.rf.reg_file[4] ;
	reg [15:0] \mchip.cpu.rf.reg_file[5] ;
	reg [15:0] \mchip.cpu.rf.reg_file[6] ;
	reg [15:0] \mchip.cpu.rf.reg_file[7] ;
	wire [2:0] \mchip.cpu.rf.rs1 ;
	wire [2:0] \mchip.cpu.rf.rs2 ;
	wire \mchip.cpu.rf.rst ;
	wire \mchip.cpu.rst ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _1039_ = (_0842_ ? _1023_ : _1025_);
	assign _1040_ = _0872_ & ~_1039_;
	assign _1041_ = _1040_ | _1038_;
	assign _1042_ = _1036_ & ~_1041_;
	assign _1043_ = (_0881_ ? _1023_ : _1042_);
	assign _1044_ = _0759_ & ~_1043_;
	assign _1045_ = ~(\mchip.cpu.pc_reg.prll_out [4] & \mchip.cpu.pc_reg.prll_out [3]);
	assign _1046_ = _0983_ & ~_1045_;
	assign _1047_ = _1046_ ^ _1739_;
	assign _1048_ = _1462_ & ~_1047_;
	assign _1049_ = _1048_ | _1044_;
	assign \mchip.cpu.pc_reg.prll_in [5] = (_0885_ ? _1022_ : _1049_);
	assign _1050_ = ~(\mchip.cpu.pc_reg.prll_out [5] & \mchip.cpu.pc_reg.prll_out [4]);
	assign _1051_ = _0988_ & ~_1050_;
	assign _1052_ = _1051_ ^ \mchip.cpu.pc_reg.prll_out [6];
	assign _1053_ = ~_1052_;
	assign _1054_ = ~(_1050_ | _0996_);
	assign _1055_ = _1054_ ^ _1789_;
	assign _1056_ = (_0843_ ? _1055_ : _1053_);
	assign _1057_ = _1056_ | _0850_;
	assign _1058_ = (_0837_ ? _1055_ : _1053_);
	assign _1059_ = _0853_ & ~_1058_;
	assign _1060_ = _1057_ & ~_1059_;
	assign _1061_ = (_0859_ ? _1055_ : _1053_);
	assign _1062_ = _0858_ & ~_1061_;
	assign _1063_ = (_0864_ ? _1055_ : _1053_);
	assign _1064_ = _0863_ & ~_1063_;
	assign _1065_ = _1064_ | _1062_;
	assign _1066_ = _1060_ & ~_1065_;
	assign _1067_ = (_0842_ ? _1055_ : _1053_);
	assign _1068_ = _0869_ & ~_1067_;
	assign _1069_ = (_0842_ ? _1053_ : _1055_);
	assign _1070_ = _0872_ & ~_1069_;
	assign _1071_ = _1070_ | _1068_;
	assign _1072_ = _1066_ & ~_1071_;
	assign _1073_ = (_0881_ ? _1053_ : _1072_);
	assign _1074_ = _0759_ & ~_1073_;
	assign _1075_ = _1046_ & ~_1739_;
	assign _1076_ = _1075_ ^ _1789_;
	assign _1077_ = _1462_ & ~_1076_;
	assign _1078_ = _1077_ | _1074_;
	assign \mchip.cpu.pc_reg.prll_in [6] = (_0885_ ? _1052_ : _1078_);
	assign _1079_ = _1051_ & ~_1789_;
	assign _1080_ = _1079_ ^ \mchip.cpu.pc_reg.prll_out [7];
	assign _1081_ = ~_1080_;
	assign _1082_ = _1054_ & ~_1789_;
	assign _1083_ = _1082_ ^ _1770_;
	assign _1084_ = (_0843_ ? _1083_ : _1081_);
	assign _1085_ = _1084_ | _0850_;
	assign _1086_ = (_0837_ ? _1083_ : _1081_);
	assign _1087_ = _0853_ & ~_1086_;
	assign _1088_ = _1085_ & ~_1087_;
	assign _1089_ = (_0859_ ? _1083_ : _1081_);
	assign _1090_ = _0858_ & ~_1089_;
	assign _1091_ = (_0864_ ? _1083_ : _1081_);
	assign _1092_ = _0863_ & ~_1091_;
	assign _1093_ = _1092_ | _1090_;
	assign _1094_ = _1088_ & ~_1093_;
	assign _1095_ = (_0842_ ? _1083_ : _1081_);
	assign _1096_ = _0869_ & ~_1095_;
	assign _1097_ = (_0842_ ? _1081_ : _1083_);
	assign _1098_ = _0872_ & ~_1097_;
	assign _1099_ = _1098_ | _1096_;
	assign _1100_ = _1094_ & ~_1099_;
	assign _1101_ = (_0881_ ? _1081_ : _1100_);
	assign _1102_ = _0759_ & ~_1101_;
	assign _1103_ = ~(\mchip.cpu.pc_reg.prll_out [6] & \mchip.cpu.pc_reg.prll_out [5]);
	assign _1104_ = _1046_ & ~_1103_;
	assign _1105_ = _1104_ ^ _1770_;
	assign _1106_ = _1462_ & ~_1105_;
	assign _1107_ = _1106_ | _1102_;
	assign \mchip.cpu.pc_reg.prll_in [7] = (_0885_ ? _1080_ : _1107_);
	assign _1108_ = ~(\mchip.cpu.pc_reg.prll_out [7] & \mchip.cpu.pc_reg.prll_out [6]);
	assign _1109_ = _1108_ | _1050_;
	assign _1110_ = _0988_ & ~_1109_;
	assign _1111_ = _1110_ ^ \mchip.cpu.pc_reg.prll_out [8];
	assign _1112_ = ~_1111_;
	assign _1113_ = ~(_1109_ | _0996_);
	assign _1114_ = _1113_ ^ _1830_;
	assign _1115_ = (_0843_ ? _1114_ : _1112_);
	assign _1116_ = _1115_ | _0850_;
	assign _1117_ = (_0837_ ? _1114_ : _1112_);
	assign _1118_ = _0853_ & ~_1117_;
	assign _1119_ = _1116_ & ~_1118_;
	assign _1120_ = (_0859_ ? _1114_ : _1112_);
	assign _1121_ = _0858_ & ~_1120_;
	assign _1122_ = (_0864_ ? _1114_ : _1112_);
	assign _1123_ = _0863_ & ~_1122_;
	assign _1124_ = _1123_ | _1121_;
	assign _1125_ = _1119_ & ~_1124_;
	assign _1126_ = (_0842_ ? _1114_ : _1112_);
	assign _1127_ = _0869_ & ~_1126_;
	assign _1128_ = (_0842_ ? _1112_ : _1114_);
	assign _1129_ = _0872_ & ~_1128_;
	assign _1130_ = _1129_ | _1127_;
	assign _1131_ = _1125_ & ~_1130_;
	assign _1132_ = (_0881_ ? _1112_ : _1131_);
	assign _1133_ = _0759_ & ~_1132_;
	assign _1134_ = _1104_ & ~_1770_;
	assign _1135_ = _1134_ ^ _1830_;
	assign _1136_ = _1462_ & ~_1135_;
	assign _1137_ = _1136_ | _1133_;
	assign \mchip.cpu.pc_reg.prll_in [8] = (_0885_ ? _1111_ : _1137_);
	assign _1138_ = _1110_ & ~_1830_;
	assign _1139_ = _1138_ ^ \mchip.cpu.pc_reg.prll_out [9];
	assign _1140_ = ~_1139_;
	assign _1141_ = _1113_ & ~_1830_;
	assign _1142_ = _1141_ ^ _1811_;
	assign _1143_ = (_0843_ ? _1142_ : _1140_);
	assign _1144_ = _1143_ | _0850_;
	assign _1145_ = (_0837_ ? _1142_ : _1140_);
	assign _1146_ = _0853_ & ~_1145_;
	assign _1147_ = _1144_ & ~_1146_;
	assign _1148_ = (_0859_ ? _1142_ : _1140_);
	assign _1149_ = _0858_ & ~_1148_;
	assign _1150_ = (_0864_ ? _1142_ : _1140_);
	assign _1151_ = _0863_ & ~_1150_;
	assign _1152_ = _1151_ | _1149_;
	assign _1153_ = _1147_ & ~_1152_;
	assign _1154_ = (_0842_ ? _1142_ : _1140_);
	assign _1155_ = _0869_ & ~_1154_;
	assign _1156_ = (_0842_ ? _1140_ : _1142_);
	assign _1157_ = _0872_ & ~_1156_;
	assign _1158_ = _1157_ | _1155_;
	assign _1159_ = _1153_ & ~_1158_;
	assign _1160_ = (_0881_ ? _1140_ : _1159_);
	assign _1161_ = _0759_ & ~_1160_;
	assign _1162_ = ~(\mchip.cpu.pc_reg.prll_out [8] & \mchip.cpu.pc_reg.prll_out [7]);
	assign _1163_ = _1162_ | _1103_;
	assign _1164_ = _1046_ & ~_1163_;
	assign _1165_ = _1164_ ^ _1811_;
	assign _1166_ = _1462_ & ~_1165_;
	assign _1167_ = _1166_ | _1161_;
	assign \mchip.cpu.pc_reg.prll_in [9] = (_0885_ ? _1139_ : _1167_);
	assign _1168_ = ~(\mchip.cpu.pc_reg.prll_out [9] & \mchip.cpu.pc_reg.prll_out [8]);
	assign _1169_ = _1110_ & ~_1168_;
	assign _1170_ = _1169_ ^ \mchip.cpu.pc_reg.prll_out [10];
	assign _1171_ = ~_1170_;
	assign _1172_ = _1113_ & ~_1168_;
	assign _1173_ = _1172_ ^ _1868_;
	assign _1174_ = (_0843_ ? _1173_ : _1171_);
	assign _1175_ = _1174_ | _0850_;
	assign _1176_ = (_0837_ ? _1173_ : _1171_);
	assign _1177_ = _0853_ & ~_1176_;
	assign _1178_ = _1175_ & ~_1177_;
	assign _1179_ = (_0859_ ? _1173_ : _1171_);
	assign _1180_ = _0858_ & ~_1179_;
	assign _1181_ = (_0864_ ? _1173_ : _1171_);
	assign _1182_ = _0863_ & ~_1181_;
	assign _1183_ = _1182_ | _1180_;
	assign _1184_ = _1178_ & ~_1183_;
	assign _1185_ = (_0842_ ? _1173_ : _1171_);
	assign _1186_ = _0869_ & ~_1185_;
	assign _1187_ = (_0842_ ? _1171_ : _1173_);
	assign _1188_ = _0872_ & ~_1187_;
	assign _1189_ = _1188_ | _1186_;
	assign _1190_ = _1184_ & ~_1189_;
	assign _1191_ = (_0881_ ? _1171_ : _1190_);
	assign _1192_ = _0759_ & ~_1191_;
	assign _1193_ = _1164_ & ~_1811_;
	assign _1194_ = _1193_ ^ _1868_;
	assign _1195_ = _1462_ & ~_1194_;
	assign _1196_ = _1195_ | _1192_;
	assign \mchip.cpu.pc_reg.prll_in [10] = (_0885_ ? _1170_ : _1196_);
	assign _1197_ = _1169_ & ~_1868_;
	assign _1198_ = _1197_ ^ \mchip.cpu.pc_reg.prll_out [11];
	assign _1199_ = ~_1198_;
	assign _1200_ = _1172_ & ~_1868_;
	assign _1201_ = _1200_ ^ _1850_;
	assign _1202_ = (_0843_ ? _1201_ : _1199_);
	assign _1203_ = _1202_ | _0850_;
	assign _1204_ = (_0837_ ? _1201_ : _1199_);
	assign _1205_ = _0853_ & ~_1204_;
	assign _1206_ = _1203_ & ~_1205_;
	assign _1207_ = (_0859_ ? _1201_ : _1199_);
	assign _1208_ = _0858_ & ~_1207_;
	assign _1209_ = (_0864_ ? _1201_ : _1199_);
	assign _1210_ = _0863_ & ~_1209_;
	assign _1211_ = _1210_ | _1208_;
	assign _1212_ = _1206_ & ~_1211_;
	assign _1213_ = (_0842_ ? _1201_ : _1199_);
	assign _1214_ = _0869_ & ~_1213_;
	assign _1215_ = (_0842_ ? _1199_ : _1201_);
	assign _1216_ = _0872_ & ~_1215_;
	assign _1217_ = _1216_ | _1214_;
	assign _1218_ = _1212_ & ~_1217_;
	assign _1219_ = (_0881_ ? _1199_ : _1218_);
	assign _1220_ = _0759_ & ~_1219_;
	assign _1221_ = ~(\mchip.cpu.pc_reg.prll_out [10] & \mchip.cpu.pc_reg.prll_out [9]);
	assign _1222_ = _1164_ & ~_1221_;
	assign _1223_ = _1222_ ^ _1850_;
	assign _1224_ = _1462_ & ~_1223_;
	assign _1225_ = _1224_ | _1220_;
	assign \mchip.cpu.pc_reg.prll_in [11] = (_0885_ ? _1198_ : _1225_);
	assign _1226_ = ~(\mchip.cpu.pc_reg.prll_out [11] & \mchip.cpu.pc_reg.prll_out [10]);
	assign _1227_ = _1226_ | _1168_;
	assign _1228_ = _1110_ & ~_1227_;
	assign _1229_ = _1228_ ^ \mchip.cpu.pc_reg.prll_out [12];
	assign _1230_ = ~_1229_;
	assign _1231_ = _1113_ & ~_1227_;
	assign _1232_ = _1231_ ^ _1907_;
	assign _1233_ = (_0843_ ? _1232_ : _1230_);
	assign _1234_ = _1233_ | _0850_;
	assign _1235_ = (_0837_ ? _1232_ : _1230_);
	assign _1236_ = _0853_ & ~_1235_;
	assign _1237_ = _1234_ & ~_1236_;
	assign _1238_ = (_0859_ ? _1232_ : _1230_);
	assign _1239_ = _0858_ & ~_1238_;
	assign _1240_ = (_0864_ ? _1232_ : _1230_);
	assign _1241_ = _0863_ & ~_1240_;
	assign _1242_ = _1241_ | _1239_;
	assign _1243_ = _1237_ & ~_1242_;
	assign _1244_ = (_0842_ ? _1232_ : _1230_);
	assign _1245_ = _0869_ & ~_1244_;
	assign _1246_ = (_0842_ ? _1230_ : _1232_);
	assign _1247_ = _0872_ & ~_1246_;
	assign _1248_ = _1247_ | _1245_;
	assign _1249_ = _1243_ & ~_1248_;
	assign _1250_ = (_0881_ ? _1230_ : _1249_);
	assign _1251_ = _0759_ & ~_1250_;
	assign _1252_ = _1222_ & ~_1850_;
	assign _1253_ = _1252_ ^ _1907_;
	assign _1254_ = _1462_ & ~_1253_;
	assign _1255_ = _1254_ | _1251_;
	assign \mchip.cpu.pc_reg.prll_in [12] = (_0885_ ? _1229_ : _1255_);
	assign _1256_ = _1228_ & ~_1907_;
	assign _1257_ = _1256_ ^ \mchip.cpu.pc_reg.prll_out [13];
	assign _1258_ = ~_1257_;
	assign _1259_ = _1231_ & ~_1907_;
	assign _1260_ = _1259_ ^ _1889_;
	assign _1261_ = (_0843_ ? _1260_ : _1258_);
	assign _1262_ = _1261_ | _0850_;
	assign _1263_ = (_0837_ ? _1260_ : _1258_);
	assign _1264_ = _0853_ & ~_1263_;
	assign _1265_ = _1262_ & ~_1264_;
	assign _1266_ = (_0859_ ? _1260_ : _1258_);
	assign _1267_ = _0858_ & ~_1266_;
	assign _1268_ = (_0864_ ? _1260_ : _1258_);
	assign _1269_ = _0863_ & ~_1268_;
	assign _1270_ = _1269_ | _1267_;
	assign _1271_ = _1265_ & ~_1270_;
	assign _1272_ = (_0842_ ? _1260_ : _1258_);
	assign _1273_ = _0869_ & ~_1272_;
	assign _1274_ = (_0842_ ? _1258_ : _1260_);
	assign _1275_ = _0872_ & ~_1274_;
	assign _1276_ = _1275_ | _1273_;
	assign _1277_ = _1271_ & ~_1276_;
	assign _1278_ = (_0881_ ? _1258_ : _1277_);
	assign _1279_ = _0759_ & ~_1278_;
	assign _1280_ = ~(\mchip.cpu.pc_reg.prll_out [12] & \mchip.cpu.pc_reg.prll_out [11]);
	assign _1281_ = _1280_ | _1221_;
	assign _1282_ = _1164_ & ~_1281_;
	assign _1283_ = _1282_ ^ _1889_;
	assign _1284_ = _1462_ & ~_1283_;
	assign _1285_ = _1284_ | _1279_;
	assign \mchip.cpu.pc_reg.prll_in [13] = (_0885_ ? _1257_ : _1285_);
	assign _1286_ = ~(\mchip.cpu.pc_reg.prll_out [13] & \mchip.cpu.pc_reg.prll_out [12]);
	assign _1287_ = _1228_ & ~_1286_;
	assign _1288_ = _1287_ ^ \mchip.cpu.pc_reg.prll_out [14];
	assign _1289_ = ~_1288_;
	assign _1290_ = _1231_ & ~_1286_;
	assign _1291_ = _1290_ ^ _1946_;
	assign _1292_ = (_0843_ ? _1291_ : _1289_);
	assign _1293_ = _1292_ | _0850_;
	assign _1294_ = (_0837_ ? _1291_ : _1289_);
	assign _1295_ = _0853_ & ~_1294_;
	assign _1296_ = _1293_ & ~_1295_;
	assign _1297_ = (_0859_ ? _1291_ : _1289_);
	assign _1298_ = _0858_ & ~_1297_;
	assign _1299_ = (_0864_ ? _1291_ : _1289_);
	assign _1300_ = _0863_ & ~_1299_;
	assign _1301_ = _1300_ | _1298_;
	assign _1302_ = _1296_ & ~_1301_;
	assign _1303_ = (_0842_ ? _1291_ : _1289_);
	assign _1304_ = _0869_ & ~_1303_;
	assign _1305_ = (_0842_ ? _1289_ : _1291_);
	assign _1306_ = _0872_ & ~_1305_;
	assign _1307_ = _1306_ | _1304_;
	assign _1308_ = _1302_ & ~_1307_;
	assign _1309_ = (_0881_ ? _1289_ : _1308_);
	assign _1310_ = _0759_ & ~_1309_;
	assign _1311_ = _1282_ & ~_1889_;
	assign _1312_ = _1311_ ^ _1946_;
	assign _1313_ = _1462_ & ~_1312_;
	assign _1314_ = _1313_ | _1310_;
	assign \mchip.cpu.pc_reg.prll_in [14] = (_0885_ ? _1288_ : _1314_);
	assign _1315_ = _1287_ & ~_1946_;
	assign _1316_ = _1315_ ^ \mchip.cpu.pc_reg.prll_out [15];
	assign _1317_ = ~_1316_;
	assign _1318_ = _1290_ & ~_1946_;
	assign _1319_ = _1318_ ^ _1927_;
	assign _1320_ = (_0843_ ? _1319_ : _1317_);
	assign _1321_ = _1320_ | _0850_;
	assign _1322_ = (_0837_ ? _1319_ : _1317_);
	assign _1323_ = _0853_ & ~_1322_;
	assign _1324_ = _1321_ & ~_1323_;
	assign _1325_ = (_0859_ ? _1319_ : _1317_);
	assign _1326_ = _0858_ & ~_1325_;
	assign _1327_ = (_0864_ ? _1319_ : _1317_);
	assign _1328_ = _0863_ & ~_1327_;
	assign _1329_ = _1328_ | _1326_;
	assign _1330_ = _1324_ & ~_1329_;
	assign _1331_ = (_0842_ ? _1319_ : _1317_);
	assign _1332_ = _0869_ & ~_1331_;
	assign _1333_ = (_0842_ ? _1317_ : _1319_);
	assign _1334_ = _0872_ & ~_1333_;
	assign _1335_ = _1334_ | _1332_;
	assign _1336_ = _1330_ & ~_1335_;
	assign _1337_ = (_0881_ ? _1317_ : _1336_);
	assign _1338_ = _0759_ & ~_1337_;
	assign _1339_ = ~(\mchip.cpu.pc_reg.prll_out [14] & \mchip.cpu.pc_reg.prll_out [13]);
	assign _1340_ = _1282_ & ~_1339_;
	assign _1341_ = _1340_ ^ _1927_;
	assign _1342_ = _1462_ & ~_1341_;
	assign _1343_ = _1342_ | _1338_;
	assign \mchip.cpu.pc_reg.prll_in [15] = (_0885_ ? _1316_ : _1343_);
	assign _1344_ = ~(\mchip.cpu.bus_pc  | _1454_);
	assign _1345_ = _1454_ & ~\mchip.cpu.bus_pc ;
	assign _1346_ = (\mchip.cpu.bus_mar  ? _1345_ : _1344_);
	assign _1347_ = \mchip.cpu.bus_pc  & _1454_;
	assign _1348_ = _1347_ & ~\mchip.cpu.bus_mar ;
	assign _1349_ = _1348_ | _1346_;
	assign _1350_ = (\mchip.cpu.pc_reg.low_b  ? _0758_ : _1830_);
	assign _1351_ = _1350_ | ~_1348_;
	assign _1352_ = _1344_ & ~\mchip.cpu.bus_mar ;
	assign _1353_ = (\mchip.cpu.mdr_shift_reg.low_b  ? \mchip.cpu.mdr_shift_reg.prll_out [0] : \mchip.cpu.mdr_shift_reg.prll_out [8]);
	assign _1354_ = _1353_ & _1352_;
	assign _1355_ = ~(_1345_ & \mchip.cpu.bus_mar );
	assign _1356_ = (\mchip.cpu.mar_shift_reg.low_b  ? \mchip.cpu.mar_shift_reg.prll_out [0] : \mchip.cpu.mar_shift_reg.prll_out [8]);
	assign _1357_ = _1356_ & ~_1355_;
	assign _1358_ = _1357_ | _1354_;
	assign _1359_ = _1351_ & ~_1358_;
	assign io_out[0] = _1349_ & ~_1359_;
	assign _0047_ = ~\mchip.cpu.pc_reg.low_b ;
	assign _1360_ = (\mchip.cpu.mar_shift_reg.low_b  ? \mchip.cpu.mar_shift_reg.prll_out [1] : \mchip.cpu.mar_shift_reg.prll_out [9]);
	assign _1361_ = _1355_ | ~_1360_;
	assign _1362_ = (\mchip.cpu.mdr_shift_reg.low_b  ? \mchip.cpu.mdr_shift_reg.prll_out [1] : \mchip.cpu.mdr_shift_reg.prll_out [9]);
	assign _1363_ = _1362_ & _1352_;
	assign _1364_ = _1361_ & ~_1363_;
	assign _1365_ = (\mchip.cpu.pc_reg.low_b  ? _0920_ : _1811_);
	assign _1366_ = _1348_ & ~_1365_;
	assign _1367_ = _1364_ & ~_1366_;
	assign io_out[1] = _1349_ & ~_1367_;
	assign _1368_ = (\mchip.cpu.mar_shift_reg.low_b  ? \mchip.cpu.mar_shift_reg.prll_out [2] : \mchip.cpu.mar_shift_reg.prll_out [10]);
	assign _1369_ = _1355_ | ~_1368_;
	assign _1370_ = (\mchip.cpu.mdr_shift_reg.low_b  ? \mchip.cpu.mdr_shift_reg.prll_out [2] : \mchip.cpu.mdr_shift_reg.prll_out [10]);
	assign _1371_ = _1370_ & _1352_;
	assign _1372_ = _1369_ & ~_1371_;
	assign _1373_ = (\mchip.cpu.pc_reg.low_b  ? _1726_ : _1868_);
	assign _1374_ = _1348_ & ~_1373_;
	assign _1375_ = _1372_ & ~_1374_;
	assign io_out[2] = _1349_ & ~_1375_;
	assign _1376_ = (\mchip.cpu.mar_shift_reg.low_b  ? \mchip.cpu.mar_shift_reg.prll_out [3] : \mchip.cpu.mar_shift_reg.prll_out [11]);
	assign _1377_ = _1355_ | ~_1376_;
	assign _1378_ = (\mchip.cpu.mdr_shift_reg.low_b  ? \mchip.cpu.mdr_shift_reg.prll_out [3] : \mchip.cpu.mdr_shift_reg.prll_out [11]);
	assign _1379_ = _1378_ & _1352_;
	assign _1380_ = _1377_ & ~_1379_;
	assign _1381_ = (\mchip.cpu.pc_reg.low_b  ? _1715_ : _1850_);
	assign _1382_ = _1348_ & ~_1381_;
	assign _1383_ = _1380_ & ~_1382_;
	assign io_out[3] = _1349_ & ~_1383_;
	assign _1384_ = (\mchip.cpu.mar_shift_reg.low_b  ? \mchip.cpu.mar_shift_reg.prll_out [4] : \mchip.cpu.mar_shift_reg.prll_out [12]);
	assign _1385_ = _1355_ | ~_1384_;
	assign _1386_ = (\mchip.cpu.mdr_shift_reg.low_b  ? \mchip.cpu.mdr_shift_reg.prll_out [4] : \mchip.cpu.mdr_shift_reg.prll_out [12]);
	assign _1387_ = _1386_ & _1352_;
	assign _1388_ = _1385_ & ~_1387_;
	assign _1389_ = (\mchip.cpu.pc_reg.low_b  ? _1758_ : _1907_);
	assign _1390_ = _1348_ & ~_1389_;
	assign _1391_ = _1388_ & ~_1390_;
	assign io_out[4] = _1349_ & ~_1391_;
	assign _1392_ = (\mchip.cpu.mar_shift_reg.low_b  ? \mchip.cpu.mar_shift_reg.prll_out [5] : \mchip.cpu.mar_shift_reg.prll_out [13]);
	assign _1393_ = _1355_ | ~_1392_;
	assign _1394_ = (\mchip.cpu.mdr_shift_reg.low_b  ? \mchip.cpu.mdr_shift_reg.prll_out [5] : \mchip.cpu.mdr_shift_reg.prll_out [13]);
	assign _1395_ = _1394_ & _1352_;
	assign _1396_ = _1393_ & ~_1395_;
	assign _1397_ = (\mchip.cpu.pc_reg.low_b  ? _1739_ : _1889_);
	assign _1398_ = _1348_ & ~_1397_;
	assign _1399_ = _1396_ & ~_1398_;
	assign io_out[5] = _1349_ & ~_1399_;
	assign _1400_ = (\mchip.cpu.mar_shift_reg.low_b  ? \mchip.cpu.mar_shift_reg.prll_out [6] : \mchip.cpu.mar_shift_reg.prll_out [14]);
	assign _1401_ = _1355_ | ~_1400_;
	assign _1402_ = (\mchip.cpu.mdr_shift_reg.low_b  ? \mchip.cpu.mdr_shift_reg.prll_out [6] : \mchip.cpu.mdr_shift_reg.prll_out [14]);
	assign _1403_ = _1402_ & _1352_;
	assign _1404_ = _1401_ & ~_1403_;
	assign _1405_ = (\mchip.cpu.pc_reg.low_b  ? _1789_ : _1946_);
	assign _1406_ = _1348_ & ~_1405_;
	assign _1407_ = _1404_ & ~_1406_;
	assign io_out[6] = _1349_ & ~_1407_;
	assign _1408_ = (\mchip.cpu.mar_shift_reg.low_b  ? \mchip.cpu.mar_shift_reg.prll_out [7] : \mchip.cpu.mar_shift_reg.prll_out [15]);
	assign _1409_ = _1355_ | ~_1408_;
	assign _1410_ = (\mchip.cpu.mdr_shift_reg.low_b  ? \mchip.cpu.mdr_shift_reg.prll_out [7] : \mchip.cpu.mdr_shift_reg.prll_out [15]);
	assign _1411_ = _1410_ & _1352_;
	assign _1412_ = _1409_ & ~_1411_;
	assign _1413_ = (\mchip.cpu.pc_reg.low_b  ? _1770_ : _1927_);
	assign _1414_ = _1348_ & ~_1413_;
	assign _1415_ = _1412_ & ~_1414_;
	assign io_out[7] = _1349_ & ~_1415_;
	assign _0030_ = ~\mchip.cpu.mdr_shift_reg.low_b ;
	assign _0029_ = ~\mchip.cpu.mar_shift_reg.low_b ;
	assign _2028_[0] = ~\mchip.cpu.instr_shift.count [0];
	assign _1416_ = \mchip.cpu.ctrl_fsm.halt  | io_in[13];
	assign _1417_ = _1416_ | ~_1467_;
	assign _0002_ = \mchip.cpu.ctrl_fsm.cs [7] & ~_1417_;
	assign _0006_ = \mchip.cpu.ctrl_fsm.cs [10] & ~io_in[13];
	assign _1418_ = io_in[13] | ~io_in[8];
	assign _0007_ = \mchip.cpu.ctrl_fsm.cs [13] & ~_1418_;
	assign _0008_ = \mchip.cpu.ctrl_fsm.cs [4] & ~io_in[13];
	assign _1419_ = _1536_ | _1490_;
	assign _0048_ = _1488_ & ~_1419_;
	assign _1420_ = io_in[13] | ~_1449_;
	assign _1421_ = _1420_ | _1442_;
	assign _0000_ = \mchip.cpu.ctrl_fsm.cs [6] & ~_1421_;
	assign _0001_ = \mchip.cpu.ctrl_fsm.cs [5] & ~io_in[13];
	assign _0005_ = \mchip.cpu.ctrl_fsm.cs [2] & ~_0028_;
	assign _0004_ = \mchip.cpu.ctrl_fsm.cs [0] & ~_1418_;
	assign _0003_ = \mchip.cpu.ctrl_fsm.cs [11] & ~io_in[13];
	assign _2029_[1] = \mchip.cpu.instr_shift.count [1] ^ \mchip.cpu.instr_shift.count [0];
	assign _2029_[2] = _1496_ ^ \mchip.cpu.instr_shift.count [2];
	assign _1422_ = _1496_ & \mchip.cpu.instr_shift.count [2];
	assign _2029_[3] = _1422_ ^ \mchip.cpu.instr_shift.count [3];
	assign _1423_ = ~(\mchip.cpu.instr_shift.count [2] & \mchip.cpu.instr_shift.count [3]);
	assign _1424_ = _1496_ & ~_1423_;
	assign _2029_[4] = _1424_ ^ \mchip.cpu.instr_shift.count [4];
	assign _1425_ = ~\mchip.cpu.instr_shift.instruction [2];
	assign _1426_ = \mchip.cpu.instr_shift.instruction [0] | \mchip.cpu.instr_shift.instruction [1];
	assign _1427_ = _1426_ | _1425_;
	assign _1428_ = \mchip.cpu.instr_shift.instruction [12] & ~_1427_;
	assign _1429_ = \mchip.cpu.instr_shift.instruction [13] & ~_1427_;
	assign _1430_ = _1428_ & ~_1429_;
	assign _1431_ = \mchip.cpu.instr_shift.instruction [15] & ~_1427_;
	assign _1432_ = ~\mchip.cpu.instr_shift.instruction [14];
	assign _1433_ = _1427_ | _1432_;
	assign _1434_ = _1433_ & ~_1431_;
	assign _1435_ = _1434_ & _1430_;
	assign _1436_ = ~(_1429_ | _1428_);
	assign _1437_ = _1436_ & _1434_;
	assign _1438_ = _1429_ & ~_1428_;
	assign _1439_ = _1438_ & _1434_;
	assign _1440_ = _1439_ | _1437_;
	assign _1441_ = _1440_ | _1435_;
	assign _1442_ = _1441_ & ~_1427_;
	assign _1443_ = _1433_ | _1431_;
	assign _1444_ = _1430_ & ~_1443_;
	assign _1445_ = _1436_ & ~_1443_;
	assign _1446_ = _1438_ & ~_1443_;
	assign _1447_ = _1446_ | _1445_;
	assign _1448_ = _1447_ | _1444_;
	assign _1449_ = _1448_ & ~_1427_;
	assign _1450_ = ~(_1449_ | _1442_);
	assign _1451_ = \mchip.cpu.ctrl_fsm.cs [6] & ~_1450_;
	assign _1452_ = ~(_1451_ | \mchip.cpu.ctrl_fsm.cs [9]);
	assign _1453_ = ~(\mchip.cpu.ctrl_fsm.cs [9] | \mchip.cpu.ctrl_fsm.cs [6]);
	assign \mchip.cpu.bus_mar  = ~(_1453_ | _1452_);
	assign _1454_ = ~(\mchip.cpu.ctrl_fsm.cs [3] | \mchip.cpu.ctrl_fsm.cs [11]);
	assign \mchip.cpu.bus_mdr  = ~_1454_;
	assign \mchip.cpu.bus_pc  = \mchip.cpu.ctrl_fsm.cs [4] | \mchip.cpu.ctrl_fsm.cs [10];
	assign _1455_ = ~\mchip.cpu.instr_shift.count [4];
	assign _1456_ = \mchip.cpu.instr_shift.count [2] | \mchip.cpu.instr_shift.count [3];
	assign _1457_ = \mchip.cpu.instr_shift.count [0] | ~\mchip.cpu.instr_shift.count [1];
	assign _1458_ = _1457_ | _1456_;
	assign _1459_ = _1455_ & ~_1458_;
	assign _1460_ = \mchip.cpu.instr_shift.instruction [1] | ~\mchip.cpu.instr_shift.instruction [0];
	assign _1461_ = _1460_ | \mchip.cpu.instr_shift.instruction [2];
	assign _1462_ = ~(_1461_ & _1427_);
	assign _1463_ = \mchip.cpu.instr_shift.count [1] | \mchip.cpu.instr_shift.count [0];
	assign _1464_ = \mchip.cpu.instr_shift.count [3] | ~\mchip.cpu.instr_shift.count [2];
	assign _1465_ = _1464_ | _1463_;
	assign _1466_ = _1455_ & ~_1465_;
	assign _1467_ = (_1462_ ? _1466_ : _1459_);
	assign _1468_ = \mchip.cpu.instr_shift.instruction [1] & ~\mchip.cpu.instr_shift.instruction [0];
	assign _1469_ = ~(_1468_ & \mchip.cpu.instr_shift.instruction [2]);
	assign \mchip.cpu.ctrl_fsm.halt  = _1467_ & ~_1469_;
	assign _0028_ = io_in[13] | ~io_in[9];
	assign _1470_ = _1467_ | io_in[13];
	assign _1471_ = \mchip.cpu.ctrl_fsm.cs [7] & ~_1470_;
	assign _1472_ = \mchip.cpu.ctrl_fsm.cs [8] & ~_0028_;
	assign _0013_ = _1472_ | _1471_;
	assign _1473_ = \mchip.cpu.instr_shift.instruction [1] | \mchip.cpu.instr_shift.instruction [2];
	assign _1474_ = _1473_ & _1427_;
	assign _1475_ = ~(\mchip.cpu.instr_shift.instruction [15] | \mchip.cpu.instr_shift.instruction [14]);
	assign _1476_ = \mchip.cpu.instr_shift.instruction [13] & ~\mchip.cpu.instr_shift.instruction [12];
	assign _1477_ = ~(_1476_ & _1475_);
	assign _1478_ = \mchip.cpu.instr_shift.instruction [13] | \mchip.cpu.instr_shift.instruction [12];
	assign _1479_ = _1475_ & ~_1478_;
	assign _1480_ = _1477_ & ~_1479_;
	assign _1481_ = \mchip.cpu.instr_shift.instruction [13] | ~\mchip.cpu.instr_shift.instruction [12];
	assign _1482_ = _1475_ & ~_1481_;
	assign _1483_ = _1482_ | ~_1480_;
	assign _1484_ = _1483_ & ~_1427_;
	assign _1485_ = _1473_ & ~_1484_;
	assign _1486_ = ~(_1485_ | _1474_);
	assign _1487_ = _1486_ & _1467_;
	assign _1488_ = _1487_ & ~io_in[13];
	assign _1489_ = (\mchip.cpu.instr_shift.instruction [0] ? \mchip.cpu.instr_shift.instruction [2] : \mchip.cpu.instr_shift.instruction [1]);
	assign _1490_ = \mchip.cpu.instr_shift.instruction [9] & ~_1489_;
	assign _1491_ = ~_1490_;
	assign _1492_ = \mchip.cpu.instr_shift.instruction [11] & ~_1489_;
	assign _1493_ = \mchip.cpu.instr_shift.instruction [10] & ~_1489_;
	assign _1494_ = _1492_ | ~_1493_;
	assign _1495_ = _1494_ | _1491_;
	assign _0051_ = _1488_ & ~_1495_;
	assign _0019_ = _0051_ | io_in[13];
	assign _1496_ = \mchip.cpu.instr_shift.count [1] & \mchip.cpu.instr_shift.count [0];
	assign _1497_ = _1496_ | _1456_;
	assign _1498_ = _1497_ | \mchip.cpu.instr_shift.count [4];
	assign _1499_ = ~(_1498_ | _1459_);
	assign _1500_ = io_in[9] & ~_1499_;
	assign _1501_ = _1465_ & _1456_;
	assign _1502_ = _1501_ | \mchip.cpu.instr_shift.count [4];
	assign _1503_ = _1502_ | _1466_;
	assign _1504_ = ~(_1503_ | _1461_);
	assign _1505_ = _1427_ & ~_1504_;
	assign _0026_ = _1500_ & ~_1505_;
	assign _1506_ = ~io_in[9];
	assign _0025_ = _1499_ & ~_1506_;
	assign \mchip.cpu.mar_shift_reg.load  = \mchip.cpu.ctrl_fsm.cs [1] & ~_1427_;
	assign _0024_ = \mchip.cpu.bus_mar  & ~\mchip.cpu.mar_shift_reg.load ;
	assign _1507_ = ~(\mchip.cpu.ctrl_fsm.cs [12] | \mchip.cpu.ctrl_fsm.cs [5]);
	assign _0014_ = \mchip.cpu.mar_shift_reg.load  | ~_1507_;
	assign _1508_ = io_in[8] | io_in[13];
	assign _1509_ = \mchip.cpu.ctrl_fsm.cs [0] & ~_1508_;
	assign _1510_ = io_in[9] | io_in[13];
	assign _1511_ = \mchip.cpu.ctrl_fsm.cs [8] & ~_1510_;
	assign _1512_ = _1511_ | _1509_;
	assign _1513_ = io_in[13] | ~_1427_;
	assign _1514_ = \mchip.cpu.ctrl_fsm.cs [1] & ~_1513_;
	assign _1515_ = _1514_ | \mchip.cpu.ctrl_fsm.cs [12];
	assign _1516_ = io_in[13] | \mchip.cpu.ctrl_fsm.cs [3];
	assign _1517_ = _1516_ | _1515_;
	assign _0009_ = _1517_ | _1512_;
	assign _1518_ = _1427_ | io_in[13];
	assign _1519_ = \mchip.cpu.ctrl_fsm.cs [1] & ~_1518_;
	assign _1520_ = \mchip.cpu.ctrl_fsm.cs [13] & ~_1508_;
	assign _0010_ = _1520_ | _1519_;
	assign _1521_ = _1493_ | ~_1492_;
	assign _1522_ = _1521_ | _1491_;
	assign _0053_ = _1488_ & ~_1522_;
	assign _0017_ = _0053_ | io_in[13];
	assign _1523_ = _1521_ | _1490_;
	assign _0052_ = _1488_ & ~_1523_;
	assign _0018_ = _0052_ | io_in[13];
	assign _1524_ = ~(_1493_ & _1492_);
	assign _1525_ = _1524_ | _1490_;
	assign _0054_ = _1488_ & ~_1525_;
	assign _0016_ = _0054_ | io_in[13];
	assign _1526_ = \mchip.cpu.mar_shift_reg.load  | _1454_;
	assign _0023_ = _1507_ & ~_1526_;
	assign _1527_ = _1449_ | io_in[13];
	assign _1528_ = _1527_ | _1442_;
	assign _1529_ = \mchip.cpu.ctrl_fsm.cs [6] & ~_1528_;
	assign _1530_ = \mchip.cpu.ctrl_fsm.cs [9] & ~io_in[13];
	assign _0012_ = _1530_ | _1529_;
	assign _0022_ = \mchip.cpu.bus_pc  & ~\mchip.cpu.ctrl_fsm.cs [1];
	assign _1531_ = io_in[13] | ~_1442_;
	assign _1532_ = \mchip.cpu.ctrl_fsm.cs [6] & ~_1531_;
	assign _1533_ = \mchip.cpu.ctrl_fsm.cs [2] & ~_1510_;
	assign _0011_ = _1533_ | _1532_;
	assign _1534_ = _1524_ | _1491_;
	assign _0055_ = _1488_ & ~_1534_;
	assign _0015_ = _0055_ | io_in[13];
	assign _0027_ = \mchip.cpu.ctrl_fsm.cs [1] & ~_1462_;
	assign _1535_ = _1494_ | _1490_;
	assign _0050_ = _1488_ & ~_1535_;
	assign _0020_ = _0050_ | io_in[13];
	assign _1536_ = _1493_ | _1492_;
	assign _1537_ = _1536_ | _1491_;
	assign _0049_ = _1488_ & ~_1537_;
	assign _0021_ = _0049_ | io_in[13];
	assign _1538_ = ~(\mchip.cpu.instr_shift.instruction [0] | \mchip.cpu.instr_shift.instruction [1]);
	assign _1539_ = (\mchip.cpu.instr_shift.instruction [2] ? _1538_ : _1468_);
	assign _1540_ = _1473_ & ~_1539_;
	assign _1541_ = \mchip.cpu.instr_shift.instruction [5] & ~_1540_;
	assign _1542_ = \mchip.cpu.instr_shift.instruction [4] & ~_1540_;
	assign _1543_ = \mchip.cpu.instr_shift.instruction [3] & ~_1540_;
	assign _1544_ = _1543_ | _1542_;
	assign _1545_ = ~(_1544_ | _1541_);
	assign _1546_ = ~_1545_;
	assign _1547_ = ~\mchip.cpu.rf.reg_file[6] [0];
	assign _1548_ = ~\mchip.cpu.rf.reg_file[7] [0];
	assign _1549_ = (_1543_ ? _1548_ : _1547_);
	assign _1550_ = ~\mchip.cpu.rf.reg_file[4] [0];
	assign _1551_ = ~\mchip.cpu.rf.reg_file[5] [0];
	assign _1552_ = (_1543_ ? _1551_ : _1550_);
	assign _1553_ = (_1542_ ? _1549_ : _1552_);
	assign _1554_ = ~\mchip.cpu.rf.reg_file[2] [0];
	assign _1555_ = ~\mchip.cpu.rf.reg_file[3] [0];
	assign _1556_ = (_1543_ ? _1555_ : _1554_);
	assign _1557_ = ~\mchip.cpu.rf.reg_file[0] [0];
	assign _1558_ = ~\mchip.cpu.rf.reg_file[1] [0];
	assign _1559_ = (_1543_ ? _1558_ : _1557_);
	assign _1560_ = (_1542_ ? _1556_ : _1559_);
	assign _1561_ = (_1541_ ? _1553_ : _1560_);
	assign _1562_ = _1546_ & ~_1561_;
	assign _1563_ = \mchip.cpu.instr_shift.instruction [0] & \mchip.cpu.instr_shift.instruction [1];
	assign _1564_ = _1563_ & ~\mchip.cpu.instr_shift.instruction [2];
	assign _1565_ = (_1564_ ? \mchip.cpu.pc_reg.prll_out [0] : _1562_);
	assign _1566_ = (\mchip.cpu.instr_shift.instruction [2] ? _1538_ : _1563_);
	assign _1567_ = _1461_ & ~_1566_;
	assign _1568_ = _1426_ | \mchip.cpu.instr_shift.instruction [2];
	assign _1569_ = _1568_ & ~_1539_;
	assign _1570_ = \mchip.cpu.instr_shift.instruction [8] & ~_1569_;
	assign _1571_ = _1569_ | ~\mchip.cpu.instr_shift.instruction [6];
	assign _1572_ = \mchip.cpu.instr_shift.instruction [7] & ~_1569_;
	assign _1573_ = _1572_ | ~_1571_;
	assign _1574_ = ~(_1573_ | _1570_);
	assign _1575_ = (_1571_ ? _1547_ : _1548_);
	assign _1576_ = (_1571_ ? _1550_ : _1551_);
	assign _1577_ = (_1572_ ? _1575_ : _1576_);
	assign _1578_ = (_1571_ ? _1554_ : _1555_);
	assign _1579_ = (_1571_ ? _1557_ : _1558_);
	assign _1580_ = (_1572_ ? _1578_ : _1579_);
	assign _1581_ = (_1570_ ? _1577_ : _1580_);
	assign _1582_ = _1581_ | _1574_;
	assign _1583_ = ~_1582_;
	assign _1584_ = (_1448_ ? \mchip.cpu.instr_shift.imm [0] : _1583_);
	assign _1585_ = (_1441_ ? \mchip.cpu.instr_shift.imm [0] : _1584_);
	assign _1586_ = _1585_ & ~_1427_;
	assign _1587_ = \mchip.cpu.instr_shift.imm [0] & ~_1461_;
	assign _1588_ = _1587_ | _1586_;
	assign _1589_ = (_1567_ ? _1583_ : _1588_);
	assign _1590_ = _1589_ | _1565_;
	assign _1591_ = _1589_ & _1565_;
	assign _1592_ = _1590_ & ~_1591_;
	assign _1593_ = \mchip.cpu.instr_shift.instruction [14] & ~_1473_;
	assign _1594_ = \mchip.cpu.instr_shift.instruction [15] & ~_1473_;
	assign _1595_ = _1593_ & ~_1594_;
	assign _1596_ = \mchip.cpu.instr_shift.instruction [13] & ~_1473_;
	assign _1597_ = \mchip.cpu.instr_shift.instruction [12] & ~_1473_;
	assign _1598_ = _1597_ | _1596_;
	assign _1599_ = _1595_ & ~_1598_;
	assign _1600_ = ~\mchip.cpu.rf.reg_file[6] [1];
	assign _1601_ = ~\mchip.cpu.rf.reg_file[7] [1];
	assign _1602_ = (_1571_ ? _1600_ : _1601_);
	assign _1603_ = ~\mchip.cpu.rf.reg_file[4] [1];
	assign _1604_ = ~\mchip.cpu.rf.reg_file[5] [1];
	assign _1605_ = (_1571_ ? _1603_ : _1604_);
	assign _1606_ = (_1572_ ? _1602_ : _1605_);
	assign _1607_ = ~\mchip.cpu.rf.reg_file[2] [1];
	assign _1608_ = ~\mchip.cpu.rf.reg_file[3] [1];
	assign _1609_ = (_1571_ ? _1607_ : _1608_);
	assign _1610_ = ~\mchip.cpu.rf.reg_file[0] [1];
	assign _1611_ = ~\mchip.cpu.rf.reg_file[1] [1];
	assign _1612_ = (_1571_ ? _1610_ : _1611_);
	assign _1613_ = (_1572_ ? _1609_ : _1612_);
	assign _1614_ = (_1570_ ? _1606_ : _1613_);
	assign _1615_ = _1574_ | _1614_;
	assign _1616_ = \mchip.cpu.instr_shift.imm [1] & ~_1461_;
	assign _1617_ = ~_1615_;
	assign _1618_ = (_1448_ ? \mchip.cpu.instr_shift.imm [1] : _1617_);
	assign _1619_ = (_1441_ ? \mchip.cpu.instr_shift.imm [1] : _1618_);
	assign _1620_ = _1619_ & ~_1427_;
	assign _1621_ = ~(_1620_ | _1616_);
	assign _1622_ = (_1567_ ? _1615_ : _1621_);
	assign _1623_ = ~_1622_;
	assign _1624_ = _1589_ | ~_1565_;
	assign _1625_ = _1624_ | _1623_;
	assign _1626_ = ~\mchip.cpu.rf.reg_file[6] [2];
	assign _1627_ = ~\mchip.cpu.rf.reg_file[7] [2];
	assign _1628_ = (_1571_ ? _1626_ : _1627_);
	assign _1629_ = ~\mchip.cpu.rf.reg_file[4] [2];
	assign _1630_ = ~\mchip.cpu.rf.reg_file[5] [2];
	assign _1631_ = (_1571_ ? _1629_ : _1630_);
	assign _1632_ = (_1572_ ? _1628_ : _1631_);
	assign _1633_ = ~\mchip.cpu.rf.reg_file[2] [2];
	assign _1634_ = ~\mchip.cpu.rf.reg_file[3] [2];
	assign _1635_ = (_1571_ ? _1633_ : _1634_);
	assign _1636_ = ~\mchip.cpu.rf.reg_file[0] [2];
	assign _1637_ = ~\mchip.cpu.rf.reg_file[1] [2];
	assign _1638_ = (_1571_ ? _1636_ : _1637_);
	assign _1639_ = (_1572_ ? _1635_ : _1638_);
	assign _1640_ = (_1570_ ? _1632_ : _1639_);
	assign _1641_ = _1640_ | _1574_;
	assign _1642_ = ~_1641_;
	assign _1643_ = \mchip.cpu.instr_shift.imm [2] & ~_1461_;
	assign _1644_ = ~\mchip.cpu.instr_shift.imm [2];
	assign _1645_ = (_1448_ ? _1644_ : _1641_);
	assign _1646_ = (_1441_ ? _1644_ : _1645_);
	assign _1647_ = ~(_1646_ | _1427_);
	assign _1648_ = _1647_ | _1564_;
	assign _1649_ = _1648_ | _1643_;
	assign _1650_ = (_1567_ ? _1642_ : _1649_);
	assign _1651_ = _1650_ | _1625_;
	assign _1652_ = ~\mchip.cpu.rf.reg_file[6] [3];
	assign _1653_ = ~\mchip.cpu.rf.reg_file[7] [3];
	assign _1654_ = (_1571_ ? _1652_ : _1653_);
	assign _1655_ = ~\mchip.cpu.rf.reg_file[4] [3];
	assign _1656_ = ~\mchip.cpu.rf.reg_file[5] [3];
	assign _1657_ = (_1571_ ? _1655_ : _1656_);
	assign _1658_ = (_1572_ ? _1654_ : _1657_);
	assign _1659_ = ~\mchip.cpu.rf.reg_file[2] [3];
	assign _1660_ = ~\mchip.cpu.rf.reg_file[3] [3];
	assign _1661_ = (_1571_ ? _1659_ : _1660_);
	assign _1662_ = ~\mchip.cpu.rf.reg_file[0] [3];
	assign _1663_ = ~\mchip.cpu.rf.reg_file[1] [3];
	assign _1664_ = (_1571_ ? _1662_ : _1663_);
	assign _1665_ = (_1572_ ? _1661_ : _1664_);
	assign _1666_ = (_1570_ ? _1658_ : _1665_);
	assign _1667_ = _1666_ | _1574_;
	assign _1668_ = ~_1667_;
	assign _1669_ = \mchip.cpu.instr_shift.imm [3] & ~_1461_;
	assign _1670_ = (_1448_ ? \mchip.cpu.instr_shift.imm [3] : _1668_);
	assign _1671_ = (_1441_ ? \mchip.cpu.instr_shift.imm [3] : _1670_);
	assign _1672_ = _1671_ & ~_1427_;
	assign _1673_ = _1672_ | _1669_;
	assign _1674_ = (_1567_ ? _1668_ : _1673_);
	assign _1675_ = _1674_ | _1651_;
	assign _1676_ = ~\mchip.cpu.rf.reg_file[6] [4];
	assign _1677_ = ~\mchip.cpu.rf.reg_file[7] [4];
	assign _1678_ = (_1571_ ? _1676_ : _1677_);
	assign _1679_ = ~\mchip.cpu.rf.reg_file[4] [4];
	assign _1680_ = ~\mchip.cpu.rf.reg_file[5] [4];
	assign _1681_ = (_1571_ ? _1679_ : _1680_);
	assign _1682_ = (_1572_ ? _1678_ : _1681_);
	assign _1683_ = ~\mchip.cpu.rf.reg_file[2] [4];
	assign _1684_ = ~\mchip.cpu.rf.reg_file[3] [4];
	assign _1685_ = (_1571_ ? _1683_ : _1684_);
	assign _1686_ = ~\mchip.cpu.rf.reg_file[0] [4];
	assign _1687_ = ~\mchip.cpu.rf.reg_file[1] [4];
	assign _1688_ = (_1571_ ? _1686_ : _1687_);
	assign _1689_ = (_1572_ ? _1685_ : _1688_);
	assign _1690_ = (_1570_ ? _1682_ : _1689_);
	assign _1691_ = _1690_ | _1574_;
	assign _1692_ = ~_1691_;
	assign _1693_ = \mchip.cpu.instr_shift.imm [4] & ~_1461_;
	assign _1694_ = (_1448_ ? \mchip.cpu.instr_shift.imm [4] : _1692_);
	assign _1695_ = (_1441_ ? \mchip.cpu.instr_shift.imm [4] : _1694_);
	assign _1696_ = _1695_ & ~_1427_;
	assign _1697_ = _1696_ | _1693_;
	assign _1698_ = (_1567_ ? _1692_ : _1697_);
	assign _1699_ = _1698_ | _1675_;
	assign _1700_ = _1599_ & ~_1699_;
	assign _1701_ = _1597_ & ~_1596_;
	assign _1702_ = _1701_ & _1595_;
	assign _1703_ = ~_1565_;
	assign _1704_ = (_1543_ ? _1601_ : _1600_);
	assign _1705_ = (_1543_ ? _1604_ : _1603_);
	assign _1706_ = (_1542_ ? _1704_ : _1705_);
	assign _1707_ = (_1543_ ? _1608_ : _1607_);
	assign _1708_ = (_1543_ ? _1611_ : _1610_);
	assign _1709_ = (_1542_ ? _1707_ : _1708_);
	assign _1710_ = (_1541_ ? _1706_ : _1709_);
	assign _1711_ = _1546_ & ~_1710_;
	assign _1712_ = (_1564_ ? \mchip.cpu.pc_reg.prll_out [1] : _1711_);
	assign _1713_ = ~_1712_;
	assign _1714_ = (_1589_ ? _1713_ : _1703_);
	assign _1715_ = ~\mchip.cpu.pc_reg.prll_out [3];
	assign _1716_ = (_1543_ ? _1653_ : _1652_);
	assign _1717_ = (_1543_ ? _1656_ : _1655_);
	assign _1718_ = (_1542_ ? _1716_ : _1717_);
	assign _1719_ = (_1543_ ? _1660_ : _1659_);
	assign _1720_ = (_1543_ ? _1663_ : _1662_);
	assign _1721_ = (_1542_ ? _1719_ : _1720_);
	assign _1722_ = (_1541_ ? _1718_ : _1721_);
	assign _1723_ = _1546_ & ~_1722_;
	assign _1724_ = ~_1723_;
	assign _1725_ = (_1564_ ? _1715_ : _1724_);
	assign _1726_ = ~\mchip.cpu.pc_reg.prll_out [2];
	assign _1727_ = (_1543_ ? _1627_ : _1626_);
	assign _1728_ = (_1543_ ? _1630_ : _1629_);
	assign _1729_ = (_1542_ ? _1727_ : _1728_);
	assign _1730_ = (_1543_ ? _1634_ : _1633_);
	assign _1731_ = (_1543_ ? _1637_ : _1636_);
	assign _1732_ = (_1542_ ? _1730_ : _1731_);
	assign _1733_ = (_1541_ ? _1729_ : _1732_);
	assign _1734_ = _1546_ & ~_1733_;
	assign _1735_ = ~_1734_;
	assign _1736_ = (_1564_ ? _1726_ : _1735_);
	assign _1737_ = (_1589_ ? _1725_ : _1736_);
	assign _1738_ = (_1622_ ? _1714_ : _1737_);
	assign _1739_ = ~\mchip.cpu.pc_reg.prll_out [5];
	assign _1740_ = ~\mchip.cpu.rf.reg_file[6] [5];
	assign _1741_ = ~\mchip.cpu.rf.reg_file[7] [5];
	assign _1742_ = (_1543_ ? _1741_ : _1740_);
	assign _1743_ = ~\mchip.cpu.rf.reg_file[4] [5];
	assign _1744_ = ~\mchip.cpu.rf.reg_file[5] [5];
	assign _1745_ = (_1543_ ? _1744_ : _1743_);
	assign _1746_ = (_1542_ ? _1742_ : _1745_);
	assign _1747_ = ~\mchip.cpu.rf.reg_file[2] [5];
	assign _1748_ = ~\mchip.cpu.rf.reg_file[3] [5];
	assign _1749_ = (_1543_ ? _1748_ : _1747_);
	assign _1750_ = ~\mchip.cpu.rf.reg_file[0] [5];
	assign _1751_ = ~\mchip.cpu.rf.reg_file[1] [5];
	assign _1752_ = (_1543_ ? _1751_ : _1750_);
	assign _1753_ = (_1542_ ? _1749_ : _1752_);
	assign _1754_ = (_1541_ ? _1746_ : _1753_);
	assign _1755_ = _1546_ & ~_1754_;
	assign _1756_ = ~_1755_;
	assign _1757_ = (_1564_ ? _1739_ : _1756_);
	assign _1758_ = ~\mchip.cpu.pc_reg.prll_out [4];
	assign _1759_ = (_1543_ ? _1677_ : _1676_);
	assign _1760_ = (_1543_ ? _1680_ : _1679_);
	assign _1761_ = (_1542_ ? _1759_ : _1760_);
	assign _1762_ = (_1543_ ? _1684_ : _1683_);
	assign _1763_ = (_1543_ ? _1687_ : _1686_);
	assign _1764_ = (_1542_ ? _1762_ : _1763_);
	assign _1765_ = (_1541_ ? _1761_ : _1764_);
	assign _1766_ = _1546_ & ~_1765_;
	assign _1767_ = ~_1766_;
	assign _1768_ = (_1564_ ? _1758_ : _1767_);
	assign _1769_ = (_1589_ ? _1757_ : _1768_);
	assign _1770_ = ~\mchip.cpu.pc_reg.prll_out [7];
	assign _1771_ = ~\mchip.cpu.rf.reg_file[6] [7];
	assign _1772_ = ~\mchip.cpu.rf.reg_file[7] [7];
	assign _1773_ = (_1543_ ? _1772_ : _1771_);
	assign _1774_ = ~\mchip.cpu.rf.reg_file[4] [7];
	assign _1775_ = ~\mchip.cpu.rf.reg_file[5] [7];
	assign _1776_ = (_1543_ ? _1775_ : _1774_);
	assign _1777_ = (_1542_ ? _1773_ : _1776_);
	assign _1778_ = ~\mchip.cpu.rf.reg_file[2] [7];
	assign _1779_ = ~\mchip.cpu.rf.reg_file[3] [7];
	assign _1780_ = (_1543_ ? _1779_ : _1778_);
	assign _1781_ = ~\mchip.cpu.rf.reg_file[0] [7];
	assign _1782_ = ~\mchip.cpu.rf.reg_file[1] [7];
	assign _1783_ = (_1543_ ? _1782_ : _1781_);
	assign _1784_ = (_1542_ ? _1780_ : _1783_);
	assign _1785_ = (_1541_ ? _1777_ : _1784_);
	assign _1786_ = _1546_ & ~_1785_;
	assign _1787_ = ~_1786_;
	assign _1788_ = (_1564_ ? _1770_ : _1787_);
	assign _1789_ = ~\mchip.cpu.pc_reg.prll_out [6];
	assign _1790_ = ~\mchip.cpu.rf.reg_file[6] [6];
	assign _1791_ = ~\mchip.cpu.rf.reg_file[7] [6];
	assign _1792_ = (_1543_ ? _1791_ : _1790_);
	assign _1793_ = ~\mchip.cpu.rf.reg_file[4] [6];
	assign _1794_ = ~\mchip.cpu.rf.reg_file[5] [6];
	assign _1795_ = (_1543_ ? _1794_ : _1793_);
	assign _1796_ = (_1542_ ? _1792_ : _1795_);
	assign _1797_ = ~\mchip.cpu.rf.reg_file[2] [6];
	assign _1798_ = ~\mchip.cpu.rf.reg_file[3] [6];
	assign _1799_ = (_1543_ ? _1798_ : _1797_);
	assign _1800_ = ~\mchip.cpu.rf.reg_file[0] [6];
	assign _1801_ = ~\mchip.cpu.rf.reg_file[1] [6];
	assign _1802_ = (_1543_ ? _1801_ : _1800_);
	assign _1803_ = (_1542_ ? _1799_ : _1802_);
	assign _1804_ = (_1541_ ? _1796_ : _1803_);
	assign _1805_ = _1546_ & ~_1804_;
	assign _1806_ = ~_1805_;
	assign _1807_ = (_1564_ ? _1789_ : _1806_);
	assign _1808_ = (_1589_ ? _1788_ : _1807_);
	assign _1809_ = (_1622_ ? _1769_ : _1808_);
	assign _1810_ = (_1650_ ? _1809_ : _1738_);
	assign _1811_ = ~\mchip.cpu.pc_reg.prll_out [9];
	assign _1812_ = ~\mchip.cpu.rf.reg_file[6] [9];
	assign _1813_ = ~\mchip.cpu.rf.reg_file[7] [9];
	assign _1814_ = (_1543_ ? _1813_ : _1812_);
	assign _1815_ = ~\mchip.cpu.rf.reg_file[4] [9];
	assign _1816_ = ~\mchip.cpu.rf.reg_file[5] [9];
	assign _1817_ = (_1543_ ? _1816_ : _1815_);
	assign _1818_ = (_1542_ ? _1814_ : _1817_);
	assign _1819_ = ~\mchip.cpu.rf.reg_file[2] [9];
	assign _1820_ = ~\mchip.cpu.rf.reg_file[3] [9];
	assign _1821_ = (_1543_ ? _1820_ : _1819_);
	assign _1822_ = ~\mchip.cpu.rf.reg_file[0] [9];
	assign _1823_ = ~\mchip.cpu.rf.reg_file[1] [9];
	assign _1824_ = (_1543_ ? _1823_ : _1822_);
	assign _1825_ = (_1542_ ? _1821_ : _1824_);
	assign _1826_ = (_1541_ ? _1818_ : _1825_);
	assign _1827_ = _1546_ & ~_1826_;
	assign _1828_ = ~_1827_;
	assign _1829_ = (_1564_ ? _1811_ : _1828_);
	assign _1830_ = ~\mchip.cpu.pc_reg.prll_out [8];
	assign _1831_ = ~\mchip.cpu.rf.reg_file[6] [8];
	assign _1832_ = ~\mchip.cpu.rf.reg_file[7] [8];
	assign _1833_ = (_1543_ ? _1832_ : _1831_);
	assign _1834_ = ~\mchip.cpu.rf.reg_file[4] [8];
	assign _1835_ = ~\mchip.cpu.rf.reg_file[5] [8];
	assign _1836_ = (_1543_ ? _1835_ : _1834_);
	assign _1837_ = (_1542_ ? _1833_ : _1836_);
	assign _1838_ = ~\mchip.cpu.rf.reg_file[2] [8];
	assign _1839_ = ~\mchip.cpu.rf.reg_file[3] [8];
	assign _1840_ = (_1543_ ? _1839_ : _1838_);
	assign _1841_ = ~\mchip.cpu.rf.reg_file[0] [8];
	assign _1842_ = ~\mchip.cpu.rf.reg_file[1] [8];
	assign _1843_ = (_1543_ ? _1842_ : _1841_);
	assign _1844_ = (_1542_ ? _1840_ : _1843_);
	assign _1845_ = (_1541_ ? _1837_ : _1844_);
	assign _1846_ = _1546_ & ~_1845_;
	assign _1847_ = ~_1846_;
	assign _1848_ = (_1564_ ? _1830_ : _1847_);
	assign _1849_ = (_1589_ ? _1829_ : _1848_);
	assign _1850_ = ~\mchip.cpu.pc_reg.prll_out [11];
	assign _1851_ = ~\mchip.cpu.rf.reg_file[6] [11];
	assign _1852_ = ~\mchip.cpu.rf.reg_file[7] [11];
	assign _1853_ = (_1543_ ? _1852_ : _1851_);
	assign _1854_ = ~\mchip.cpu.rf.reg_file[4] [11];
	assign _1855_ = ~\mchip.cpu.rf.reg_file[5] [11];
	assign _1856_ = (_1543_ ? _1855_ : _1854_);
	assign _1857_ = (_1542_ ? _1853_ : _1856_);
	assign _1858_ = ~\mchip.cpu.rf.reg_file[2] [11];
	assign _1859_ = ~\mchip.cpu.rf.reg_file[3] [11];
	assign _1860_ = (_1543_ ? _1859_ : _1858_);
	assign _1861_ = ~\mchip.cpu.rf.reg_file[0] [11];
	assign _1862_ = ~\mchip.cpu.rf.reg_file[1] [11];
	assign _1863_ = (_1543_ ? _1862_ : _1861_);
	assign _1864_ = (_1542_ ? _1860_ : _1863_);
	assign _1865_ = (_1541_ ? _1857_ : _1864_);
	assign _1866_ = _1865_ | _1545_;
	assign _1867_ = (_1564_ ? _1850_ : _1866_);
	assign _1868_ = ~\mchip.cpu.pc_reg.prll_out [10];
	assign _1869_ = ~\mchip.cpu.rf.reg_file[6] [10];
	assign _1870_ = ~\mchip.cpu.rf.reg_file[7] [10];
	assign _1871_ = (_1543_ ? _1870_ : _1869_);
	assign _1872_ = ~\mchip.cpu.rf.reg_file[4] [10];
	assign _1873_ = ~\mchip.cpu.rf.reg_file[5] [10];
	assign _1874_ = (_1543_ ? _1873_ : _1872_);
	assign _1875_ = (_1542_ ? _1871_ : _1874_);
	assign _1876_ = ~\mchip.cpu.rf.reg_file[2] [10];
	assign _1877_ = ~\mchip.cpu.rf.reg_file[3] [10];
	assign _1878_ = (_1543_ ? _1877_ : _1876_);
	assign _1879_ = ~\mchip.cpu.rf.reg_file[0] [10];
	assign _1880_ = ~\mchip.cpu.rf.reg_file[1] [10];
	assign _1881_ = (_1543_ ? _1880_ : _1879_);
	assign _1882_ = (_1542_ ? _1878_ : _1881_);
	assign _1883_ = (_1541_ ? _1875_ : _1882_);
	assign _1884_ = _1546_ & ~_1883_;
	assign _1885_ = ~_1884_;
	assign _1886_ = (_1564_ ? _1868_ : _1885_);
	assign _1887_ = (_1589_ ? _1867_ : _1886_);
	assign _1888_ = (_1622_ ? _1849_ : _1887_);
	assign _1889_ = ~\mchip.cpu.pc_reg.prll_out [13];
	assign _1890_ = ~\mchip.cpu.rf.reg_file[6] [13];
	assign _1891_ = ~\mchip.cpu.rf.reg_file[7] [13];
	assign _1892_ = (_1543_ ? _1891_ : _1890_);
	assign _1893_ = ~\mchip.cpu.rf.reg_file[4] [13];
	assign _1894_ = ~\mchip.cpu.rf.reg_file[5] [13];
	assign _1895_ = (_1543_ ? _1894_ : _1893_);
	assign _1896_ = (_1542_ ? _1892_ : _1895_);
	assign _1897_ = ~\mchip.cpu.rf.reg_file[2] [13];
	assign _1898_ = ~\mchip.cpu.rf.reg_file[3] [13];
	assign _1899_ = (_1543_ ? _1898_ : _1897_);
	assign _1900_ = ~\mchip.cpu.rf.reg_file[0] [13];
	assign _1901_ = ~\mchip.cpu.rf.reg_file[1] [13];
	assign _1902_ = (_1543_ ? _1901_ : _1900_);
	assign _1903_ = (_1542_ ? _1899_ : _1902_);
	assign _1904_ = (_1541_ ? _1896_ : _1903_);
	assign _1905_ = _1904_ | _1545_;
	assign _1906_ = (_1564_ ? _1889_ : _1905_);
	assign _1907_ = ~\mchip.cpu.pc_reg.prll_out [12];
	assign _1908_ = ~\mchip.cpu.rf.reg_file[6] [12];
	assign _1909_ = ~\mchip.cpu.rf.reg_file[7] [12];
	assign _1910_ = (_1543_ ? _1909_ : _1908_);
	assign _1911_ = ~\mchip.cpu.rf.reg_file[4] [12];
	assign _1912_ = ~\mchip.cpu.rf.reg_file[5] [12];
	assign _1913_ = (_1543_ ? _1912_ : _1911_);
	assign _1914_ = (_1542_ ? _1910_ : _1913_);
	assign _1915_ = ~\mchip.cpu.rf.reg_file[2] [12];
	assign _1916_ = ~\mchip.cpu.rf.reg_file[3] [12];
	assign _1917_ = (_1543_ ? _1916_ : _1915_);
	assign _1918_ = ~\mchip.cpu.rf.reg_file[0] [12];
	assign _1919_ = ~\mchip.cpu.rf.reg_file[1] [12];
	assign _1920_ = (_1543_ ? _1919_ : _1918_);
	assign _1921_ = (_1542_ ? _1917_ : _1920_);
	assign _1922_ = (_1541_ ? _1914_ : _1921_);
	assign _1923_ = _1546_ & ~_1922_;
	assign _1924_ = ~_1923_;
	assign _1925_ = (_1564_ ? _1907_ : _1924_);
	assign _1926_ = (_1589_ ? _1906_ : _1925_);
	assign _1927_ = ~\mchip.cpu.pc_reg.prll_out [15];
	assign _1928_ = ~\mchip.cpu.rf.reg_file[6] [15];
	assign _1929_ = ~\mchip.cpu.rf.reg_file[7] [15];
	assign _1930_ = (_1543_ ? _1929_ : _1928_);
	assign _1931_ = ~\mchip.cpu.rf.reg_file[4] [15];
	assign _1932_ = ~\mchip.cpu.rf.reg_file[5] [15];
	assign _1933_ = (_1543_ ? _1932_ : _1931_);
	assign _1934_ = (_1542_ ? _1930_ : _1933_);
	assign _1935_ = ~\mchip.cpu.rf.reg_file[2] [15];
	assign _1936_ = ~\mchip.cpu.rf.reg_file[3] [15];
	assign _1937_ = (_1543_ ? _1936_ : _1935_);
	assign _1938_ = ~\mchip.cpu.rf.reg_file[0] [15];
	assign _1939_ = ~\mchip.cpu.rf.reg_file[1] [15];
	assign _1940_ = (_1543_ ? _1939_ : _1938_);
	assign _1941_ = (_1542_ ? _1937_ : _1940_);
	assign _1942_ = (_1541_ ? _1934_ : _1941_);
	assign _1943_ = _1546_ & ~_1942_;
	assign _1944_ = ~_1943_;
	assign _1945_ = (_1564_ ? _1927_ : _1944_);
	assign _1946_ = ~\mchip.cpu.pc_reg.prll_out [14];
	assign _1947_ = ~\mchip.cpu.rf.reg_file[6] [14];
	assign _1948_ = ~\mchip.cpu.rf.reg_file[7] [14];
	assign _1949_ = (_1543_ ? _1948_ : _1947_);
	assign _1950_ = ~\mchip.cpu.rf.reg_file[4] [14];
	assign _1951_ = ~\mchip.cpu.rf.reg_file[5] [14];
	assign _1952_ = (_1543_ ? _1951_ : _1950_);
	assign _1953_ = (_1542_ ? _1949_ : _1952_);
	assign _1954_ = ~\mchip.cpu.rf.reg_file[2] [14];
	assign _1955_ = ~\mchip.cpu.rf.reg_file[3] [14];
	assign _1956_ = (_1543_ ? _1955_ : _1954_);
	assign _1957_ = ~\mchip.cpu.rf.reg_file[0] [14];
	assign _1958_ = ~\mchip.cpu.rf.reg_file[1] [14];
	assign _1959_ = (_1543_ ? _1958_ : _1957_);
	assign _1960_ = (_1542_ ? _1956_ : _1959_);
	assign _1961_ = (_1541_ ? _1953_ : _1960_);
	assign _1962_ = _1546_ & ~_1961_;
	assign _1963_ = ~_1962_;
	assign _1964_ = (_1564_ ? _1946_ : _1963_);
	assign _1965_ = (_1589_ ? _1945_ : _1964_);
	assign _1966_ = (_1622_ ? _1926_ : _1965_);
	assign _1967_ = (_1650_ ? _1966_ : _1888_);
	assign _1968_ = (_1674_ ? _1967_ : _1810_);
	assign _1969_ = _1968_ | _1698_;
	assign _1970_ = _1702_ & ~_1969_;
	assign _1971_ = _1970_ | _1700_;
	assign _1972_ = _1597_ | ~_1596_;
	assign _1973_ = _1595_ & ~_1972_;
	assign _1974_ = (_1698_ ? _1945_ : _1968_);
	assign _1975_ = _1973_ & ~_1974_;
	assign _1976_ = ~(_1597_ & _1596_);
	assign _1977_ = _1594_ | _1593_;
	assign _1978_ = ~(_1977_ | _1976_);
	assign _1979_ = _1592_ & _1978_;
	assign _1980_ = _1979_ | _1975_;
	assign _1981_ = ~(_1977_ | _1972_);
	assign _1982_ = _1981_ & _1590_;
	assign _1983_ = _1595_ & ~_1976_;
	assign _1984_ = _1983_ & _1591_;
	assign _1985_ = _1984_ | _1982_;
	assign _1986_ = _1985_ | _1980_;
	assign _1987_ = _1986_ | _1971_;
	assign _1988_ = _1983_ | _1981_;
	assign _1989_ = _1978_ | _1973_;
	assign _1990_ = _1989_ | _1988_;
	assign _1991_ = _1595_ & ~_1596_;
	assign _1992_ = _1991_ | _1990_;
	assign \mchip.cpu.alu_result [0] = (_1992_ ? _1987_ : _1592_);
	assign _1993_ = (_1589_ ? _1703_ : _1713_);
	assign _1994_ = _1993_ | _1623_;
	assign _1995_ = _1994_ | _1650_;
	assign _1996_ = _1995_ | _1674_;
	assign _1997_ = _1996_ | _1698_;
	assign _1998_ = _1599_ & ~_1997_;
	assign _1999_ = (_1589_ ? _1736_ : _1713_);
	assign _2000_ = (_1589_ ? _1768_ : _1725_);
	assign _2001_ = (_1622_ ? _1999_ : _2000_);
	assign _2002_ = (_1589_ ? _1807_ : _1757_);
	assign _2003_ = (_1589_ ? _1848_ : _1788_);
	assign _2004_ = (_1622_ ? _2002_ : _2003_);
	assign _2005_ = (_1650_ ? _2004_ : _2001_);
	assign _2006_ = (_1589_ ? _1886_ : _1829_);
	assign _2007_ = (_1589_ ? _1925_ : _1867_);
	assign _2008_ = (_1622_ ? _2006_ : _2007_);
	assign _2009_ = (_1589_ ? _1964_ : _1906_);
	assign _2010_ = _1945_ | _1589_;
	assign _2011_ = (_1622_ ? _2009_ : _2010_);
	assign _2012_ = (_1650_ ? _2011_ : _2008_);
	assign _2013_ = (_1674_ ? _2012_ : _2005_);
	assign _2014_ = _2013_ | _1698_;
	assign _2015_ = _1702_ & ~_2014_;
	assign _2016_ = _2015_ | _1998_;
	assign _2017_ = (_1622_ ? _2009_ : _1945_);
	assign _2018_ = (_1650_ ? _2017_ : _2008_);
	assign _2019_ = (_1674_ ? _2018_ : _2005_);
	assign _2020_ = (_1698_ ? _1945_ : _2019_);
	assign _2021_ = _1973_ & ~_2020_;
	assign _2022_ = _1713_ | _1622_;
	assign _2023_ = _1622_ & ~_1712_;
	assign _2024_ = _2023_ | ~_2022_;
	assign _2025_ = _1978_ & ~_2024_;
	assign _2026_ = _2025_ | _2021_;
	assign _2027_ = _1981_ & ~_2023_;
	assign _0056_ = _1983_ & ~_2022_;
	assign _0057_ = _0056_ | _2027_;
	assign _0058_ = _0057_ | _2026_;
	assign _0059_ = _0058_ | _2016_;
	assign _0060_ = _1565_ | ~_1589_;
	assign _0061_ = ~(_1589_ ^ _1622_);
	assign _0062_ = _1701_ & ~_1977_;
	assign _0063_ = (_0062_ ? _1623_ : _0061_);
	assign _0064_ = _0063_ ^ _1712_;
	assign _0065_ = ~(_0064_ ^ _0060_);
	assign \mchip.cpu.alu_result [1] = (_1992_ ? _0059_ : _0065_);
	assign _0066_ = (_1589_ ? _1713_ : _1736_);
	assign _0067_ = (_1622_ ? _0066_ : _1624_);
	assign _0068_ = _0067_ | _1650_;
	assign _0069_ = _0068_ | _1674_;
	assign _0070_ = _0069_ | _1698_;
	assign _0071_ = _1599_ & ~_0070_;
	assign _0072_ = (_1622_ ? _1737_ : _1769_);
	assign _0073_ = (_1622_ ? _1808_ : _1849_);
	assign _0074_ = (_1650_ ? _0073_ : _0072_);
	assign _0075_ = (_1622_ ? _1887_ : _1926_);
	assign _0076_ = _1965_ | _1623_;
	assign _0077_ = (_1650_ ? _0076_ : _0075_);
	assign _0078_ = (_1674_ ? _0077_ : _0074_);
	assign _0079_ = _0078_ | _1698_;
	assign _0080_ = _1702_ & ~_0079_;
	assign _0081_ = _0080_ | _0071_;
	assign _0082_ = (_1622_ ? _1965_ : _1945_);
	assign _0083_ = (_1650_ ? _0082_ : _0075_);
	assign _0084_ = (_1674_ ? _0083_ : _0074_);
	assign _0085_ = (_1698_ ? _1945_ : _0084_);
	assign _0086_ = _1973_ & ~_0085_;
	assign _0087_ = _1736_ | ~_1650_;
	assign _0088_ = _1736_ & ~_1650_;
	assign _0089_ = _0088_ | ~_0087_;
	assign _0090_ = _1978_ & ~_0089_;
	assign _0091_ = _0090_ | _0086_;
	assign _0092_ = _1981_ & ~_0088_;
	assign _0093_ = _1983_ & ~_0087_;
	assign _0094_ = _0093_ | _0092_;
	assign _0095_ = _0094_ | _0091_;
	assign _0096_ = _0095_ | _0081_;
	assign _0097_ = _0060_ & ~_0064_;
	assign _0098_ = _1712_ & ~_0063_;
	assign _0099_ = _0098_ | _0097_;
	assign _0100_ = ~_1650_;
	assign _0101_ = _1622_ & ~_1589_;
	assign _0102_ = _0101_ ^ _1650_;
	assign _0103_ = (_0062_ ? _0100_ : _0102_);
	assign _0104_ = _0103_ ^ _1736_;
	assign _0105_ = ~(_0104_ ^ _0099_);
	assign \mchip.cpu.alu_result [2] = (_1992_ ? _0096_ : _0105_);
	assign _0106_ = (_1589_ ? _1736_ : _1725_);
	assign _0107_ = (_1622_ ? _0106_ : _1993_);
	assign _0108_ = _0107_ | _1650_;
	assign _0109_ = _0108_ | _1674_;
	assign _0110_ = _0109_ | _1698_;
	assign _0111_ = _1599_ & ~_0110_;
	assign _0112_ = (_1622_ ? _2000_ : _2002_);
	assign _0113_ = (_1622_ ? _2003_ : _2006_);
	assign _0114_ = (_1650_ ? _0113_ : _0112_);
	assign _0115_ = (_1622_ ? _2007_ : _2009_);
	assign _0116_ = _2010_ | _1623_;
	assign _0117_ = (_1650_ ? _0116_ : _0115_);
	assign _0118_ = (_1674_ ? _0117_ : _0114_);
	assign _0119_ = _0118_ | _1698_;
	assign _0120_ = _1702_ & ~_0119_;
	assign _0121_ = _0120_ | _0111_;
	assign _0122_ = (_1650_ ? _1945_ : _0115_);
	assign _0123_ = (_1674_ ? _0122_ : _0114_);
	assign _0124_ = (_1698_ ? _1945_ : _0123_);
	assign _0125_ = _1973_ & ~_0124_;
	assign _0126_ = _1725_ | ~_1674_;
	assign _0127_ = _1725_ & ~_1674_;
	assign _0128_ = _0127_ | ~_0126_;
	assign _0129_ = _1978_ & ~_0128_;
	assign _0130_ = _0129_ | _0125_;
	assign _0131_ = _1981_ & ~_0127_;
	assign _0132_ = _1983_ & ~_0126_;
	assign _0133_ = _0132_ | _0131_;
	assign _0134_ = _0133_ | _0130_;
	assign _0135_ = _0134_ | _0121_;
	assign _0136_ = _0103_ & ~_1736_;
	assign _0137_ = _0099_ & ~_0104_;
	assign _0138_ = ~(_0137_ | _0136_);
	assign _0139_ = _0101_ & ~_1650_;
	assign _0140_ = ~(_0139_ ^ _1674_);
	assign _0141_ = (_0062_ ? _1674_ : _0140_);
	assign _0142_ = ~(_0141_ ^ _1725_);
	assign _0143_ = _0142_ ^ _0138_;
	assign \mchip.cpu.alu_result [3] = (_1992_ ? _0135_ : _0143_);
	assign _0144_ = (_1589_ ? _1725_ : _1768_);
	assign _0145_ = (_1622_ ? _0144_ : _0066_);
	assign _0146_ = (_1650_ ? _1625_ : _0145_);
	assign _0147_ = _0146_ | _1674_;
	assign _0148_ = _0147_ | _1698_;
	assign _0149_ = _1599_ & ~_0148_;
	assign _0150_ = (_1650_ ? _1888_ : _1809_);
	assign _0151_ = _1966_ | _1650_;
	assign _0152_ = (_1674_ ? _0151_ : _0150_);
	assign _0153_ = _0152_ | _1698_;
	assign _0154_ = _1702_ & ~_0153_;
	assign _0155_ = _0154_ | _0149_;
	assign _0156_ = (_1650_ ? _1945_ : _1966_);
	assign _0157_ = (_1674_ ? _0156_ : _0150_);
	assign _0158_ = (_1698_ ? _1945_ : _0157_);
	assign _0159_ = _1973_ & ~_0158_;
	assign _0160_ = _1768_ | ~_1698_;
	assign _0161_ = _1768_ & ~_1698_;
	assign _0162_ = _0161_ | ~_0160_;
	assign _0163_ = _1978_ & ~_0162_;
	assign _0164_ = _0163_ | _0159_;
	assign _0165_ = _1981_ & ~_0161_;
	assign _0166_ = _1983_ & ~_0160_;
	assign _0167_ = _0166_ | _0165_;
	assign _0168_ = _0167_ | _0164_;
	assign _0169_ = _0168_ | _0155_;
	assign _0170_ = _0142_ | _0104_;
	assign _0171_ = _0099_ & ~_0170_;
	assign _0172_ = ~(_0141_ | _1725_);
	assign _0173_ = _0136_ & ~_0142_;
	assign _0174_ = _0173_ | _0172_;
	assign _0175_ = _0174_ | _0171_;
	assign _0176_ = ~_1698_;
	assign _0177_ = _1674_ | _1650_;
	assign _0178_ = _0101_ & ~_0177_;
	assign _0179_ = _0178_ ^ _1698_;
	assign _0180_ = (_0062_ ? _0176_ : _0179_);
	assign _0181_ = _0180_ ^ _1768_;
	assign _0182_ = ~(_0181_ ^ _0175_);
	assign \mchip.cpu.alu_result [4] = (_1992_ ? _0169_ : _0182_);
	assign _0183_ = (_1589_ ? _1768_ : _1757_);
	assign _0184_ = (_1622_ ? _0183_ : _0106_);
	assign _0185_ = (_1650_ ? _1994_ : _0184_);
	assign _0186_ = _0185_ | _1674_;
	assign _0187_ = _0186_ | _1698_;
	assign _0188_ = _1599_ & ~_0187_;
	assign _0189_ = (_1650_ ? _2008_ : _2004_);
	assign _0190_ = _2011_ | _1650_;
	assign _0191_ = (_1674_ ? _0190_ : _0189_);
	assign _0192_ = _0191_ | _1698_;
	assign _0193_ = _1702_ & ~_0192_;
	assign _0194_ = _0193_ | _0188_;
	assign _0195_ = (_1650_ ? _1945_ : _2017_);
	assign _0196_ = (_1674_ ? _0195_ : _0189_);
	assign _0197_ = (_1698_ ? _1945_ : _0196_);
	assign _0198_ = _1973_ & ~_0197_;
	assign _0199_ = (_1571_ ? _1740_ : _1741_);
	assign _0200_ = (_1571_ ? _1743_ : _1744_);
	assign _0201_ = (_1572_ ? _0199_ : _0200_);
	assign _0202_ = (_1571_ ? _1747_ : _1748_);
	assign _0203_ = (_1571_ ? _1750_ : _1751_);
	assign _0204_ = (_1572_ ? _0202_ : _0203_);
	assign _0205_ = (_1570_ ? _0201_ : _0204_);
	assign _0206_ = _0205_ | _1574_;
	assign _0207_ = ~_0206_;
	assign _0208_ = \mchip.cpu.instr_shift.imm [5] & ~_1461_;
	assign _0209_ = (_1448_ ? \mchip.cpu.instr_shift.imm [5] : _0207_);
	assign _0210_ = (_1441_ ? \mchip.cpu.instr_shift.imm [5] : _0209_);
	assign _0211_ = _0210_ & ~_1427_;
	assign _0212_ = _0211_ | _0208_;
	assign _0213_ = (_1567_ ? _0207_ : _0212_);
	assign _0214_ = _1757_ | ~_0213_;
	assign _0215_ = _1757_ & ~_0213_;
	assign _0216_ = _0215_ | ~_0214_;
	assign _0217_ = _1978_ & ~_0216_;
	assign _0218_ = _0217_ | _0198_;
	assign _0219_ = _1981_ & ~_0215_;
	assign _0220_ = _1983_ & ~_0214_;
	assign _0221_ = _0220_ | _0219_;
	assign _0222_ = _0221_ | _0218_;
	assign _0223_ = _0222_ | _0194_;
	assign _0224_ = _0180_ & ~_1768_;
	assign _0225_ = _0175_ & ~_0181_;
	assign _0226_ = ~(_0225_ | _0224_);
	assign _0227_ = ~_0213_;
	assign _0228_ = _0178_ & ~_1698_;
	assign _0229_ = _0228_ ^ _0213_;
	assign _0230_ = (_0062_ ? _0227_ : _0229_);
	assign _0231_ = _0230_ ^ _1757_;
	assign _0232_ = _0231_ ^ _0226_;
	assign \mchip.cpu.alu_result [5] = (_1992_ ? _0223_ : _0232_);
	assign _0233_ = (_1589_ ? _1757_ : _1807_);
	assign _0234_ = (_1622_ ? _0233_ : _0144_);
	assign _0235_ = (_1650_ ? _0067_ : _0234_);
	assign _0236_ = _0235_ | _1674_;
	assign _0237_ = _0236_ | _1698_;
	assign _0238_ = _1599_ & ~_0237_;
	assign _0239_ = (_1650_ ? _0075_ : _0073_);
	assign _0240_ = _0076_ | _1650_;
	assign _0241_ = (_1674_ ? _0240_ : _0239_);
	assign _0242_ = _0241_ | _1698_;
	assign _0243_ = _1702_ & ~_0242_;
	assign _0244_ = _0243_ | _0238_;
	assign _0245_ = (_1650_ ? _1945_ : _0082_);
	assign _0246_ = (_1674_ ? _0245_ : _0239_);
	assign _0247_ = (_1698_ ? _1945_ : _0246_);
	assign _0248_ = _1973_ & ~_0247_;
	assign _0249_ = (_1571_ ? _1790_ : _1791_);
	assign _0250_ = (_1571_ ? _1793_ : _1794_);
	assign _0251_ = (_1572_ ? _0249_ : _0250_);
	assign _0252_ = (_1571_ ? _1797_ : _1798_);
	assign _0253_ = (_1571_ ? _1800_ : _1801_);
	assign _0254_ = (_1572_ ? _0252_ : _0253_);
	assign _0255_ = (_1570_ ? _0251_ : _0254_);
	assign _0256_ = _0255_ | _1574_;
	assign _0257_ = ~_0256_;
	assign _0258_ = (_1448_ ? \mchip.cpu.instr_shift.imm [6] : _0257_);
	assign _0259_ = (_1441_ ? \mchip.cpu.instr_shift.imm [6] : _0258_);
	assign _0260_ = _0259_ & ~_1427_;
	assign _0261_ = \mchip.cpu.instr_shift.imm [6] & ~_1461_;
	assign _0262_ = _0261_ | _0260_;
	assign _0263_ = (_1567_ ? _0257_ : _0262_);
	assign _0264_ = _1807_ | ~_0263_;
	assign _0265_ = _1807_ & ~_0263_;
	assign _0266_ = _0265_ | ~_0264_;
	assign _0267_ = _1978_ & ~_0266_;
	assign _0268_ = _0267_ | _0248_;
	assign _0269_ = _1981_ & ~_0265_;
	assign _0270_ = _1983_ & ~_0264_;
	assign _0271_ = _0270_ | _0269_;
	assign _0272_ = _0271_ | _0268_;
	assign _0273_ = _0272_ | _0244_;
	assign _0274_ = _0231_ | _0181_;
	assign _0275_ = _0175_ & ~_0274_;
	assign _0276_ = _0230_ & ~_1757_;
	assign _0277_ = _0224_ & ~_0231_;
	assign _0278_ = _0277_ | _0276_;
	assign _0279_ = _0278_ | _0275_;
	assign _0280_ = ~_0263_;
	assign _0281_ = _0213_ | _1698_;
	assign _0282_ = _0178_ & ~_0281_;
	assign _0283_ = _0282_ ^ _0263_;
	assign _0284_ = (_0062_ ? _0280_ : _0283_);
	assign _0285_ = _0284_ ^ _1807_;
	assign _0286_ = ~(_0285_ ^ _0279_);
	assign \mchip.cpu.alu_result [6] = (_1992_ ? _0273_ : _0286_);
	assign _0287_ = (_1589_ ? _1807_ : _1788_);
	assign _0288_ = (_1622_ ? _0287_ : _0183_);
	assign _0289_ = (_1650_ ? _0107_ : _0288_);
	assign _0290_ = _0289_ | _1674_;
	assign _0291_ = _0290_ | _1698_;
	assign _0292_ = _1599_ & ~_0291_;
	assign _0293_ = (_1650_ ? _0115_ : _0113_);
	assign _0294_ = _0116_ | _1650_;
	assign _0295_ = (_1674_ ? _0294_ : _0293_);
	assign _0296_ = _0295_ | _1698_;
	assign _0297_ = _1702_ & ~_0296_;
	assign _0298_ = _0297_ | _0292_;
	assign _0299_ = (_1674_ ? _1945_ : _0293_);
	assign _0300_ = (_1698_ ? _1945_ : _0299_);
	assign _0301_ = _1973_ & ~_0300_;
	assign _0302_ = (_1571_ ? _1771_ : _1772_);
	assign _0303_ = (_1571_ ? _1774_ : _1775_);
	assign _0304_ = (_1572_ ? _0302_ : _0303_);
	assign _0305_ = (_1571_ ? _1778_ : _1779_);
	assign _0306_ = (_1571_ ? _1781_ : _1782_);
	assign _0307_ = (_1572_ ? _0305_ : _0306_);
	assign _0308_ = (_1570_ ? _0304_ : _0307_);
	assign _0309_ = _0308_ | _1574_;
	assign _0310_ = ~_0309_;
	assign _0311_ = \mchip.cpu.instr_shift.imm [7] & ~_1461_;
	assign _0312_ = (_1448_ ? \mchip.cpu.instr_shift.imm [7] : _0310_);
	assign _0313_ = (_1441_ ? \mchip.cpu.instr_shift.imm [7] : _0312_);
	assign _0314_ = _0313_ & ~_1427_;
	assign _0315_ = _0314_ | _0311_;
	assign _0316_ = (_1567_ ? _0310_ : _0315_);
	assign _0317_ = _1788_ | ~_0316_;
	assign _0318_ = _1788_ & ~_0316_;
	assign _0319_ = _0318_ | ~_0317_;
	assign _0320_ = _1978_ & ~_0319_;
	assign _0321_ = _0320_ | _0301_;
	assign _0322_ = _1981_ & ~_0318_;
	assign _0323_ = _1983_ & ~_0317_;
	assign _0324_ = _0323_ | _0322_;
	assign _0325_ = _0324_ | _0321_;
	assign _0326_ = _0325_ | _0298_;
	assign _0327_ = _0284_ & ~_1807_;
	assign _0328_ = _0279_ & ~_0285_;
	assign _0329_ = ~(_0328_ | _0327_);
	assign _0330_ = ~_0316_;
	assign _0331_ = _0282_ & ~_0263_;
	assign _0332_ = _0331_ ^ _0316_;
	assign _0333_ = (_0062_ ? _0330_ : _0332_);
	assign _0334_ = _0333_ ^ _1788_;
	assign _0335_ = _0334_ ^ _0329_;
	assign \mchip.cpu.alu_result [7] = (_1992_ ? _0326_ : _0335_);
	assign _0336_ = (_1589_ ? _1788_ : _1848_);
	assign _0337_ = (_1622_ ? _0336_ : _0233_);
	assign _0338_ = (_1650_ ? _0145_ : _0337_);
	assign _0339_ = (_1674_ ? _1651_ : _0338_);
	assign _0340_ = _0339_ | _1698_;
	assign _0341_ = _1599_ & ~_0340_;
	assign _0342_ = _1967_ | _1674_;
	assign _0343_ = _0342_ | _1698_;
	assign _0344_ = _1702_ & ~_0343_;
	assign _0345_ = _0344_ | _0341_;
	assign _0346_ = (_1674_ ? _1945_ : _1967_);
	assign _0347_ = (_1698_ ? _1945_ : _0346_);
	assign _0348_ = _1973_ & ~_0347_;
	assign _0349_ = (_1571_ ? _1831_ : _1832_);
	assign _0350_ = (_1571_ ? _1834_ : _1835_);
	assign _0351_ = (_1572_ ? _0349_ : _0350_);
	assign _0352_ = (_1571_ ? _1838_ : _1839_);
	assign _0353_ = (_1571_ ? _1841_ : _1842_);
	assign _0354_ = (_1572_ ? _0352_ : _0353_);
	assign _0355_ = (_1570_ ? _0351_ : _0354_);
	assign _0356_ = _0355_ | _1574_;
	assign _0357_ = ~_0356_;
	assign _0358_ = (_1448_ ? \mchip.cpu.instr_shift.imm [8] : _0357_);
	assign _0359_ = (_1441_ ? \mchip.cpu.instr_shift.imm [8] : _0358_);
	assign _0360_ = _0359_ & ~_1427_;
	assign _0361_ = \mchip.cpu.instr_shift.imm [8] & ~_1461_;
	assign _0362_ = _0361_ | _0360_;
	assign _0363_ = (_1567_ ? _0357_ : _0362_);
	assign _0364_ = _1848_ | ~_0363_;
	assign _0365_ = _1848_ & ~_0363_;
	assign _0366_ = _0365_ | ~_0364_;
	assign _0367_ = _1978_ & ~_0366_;
	assign _0368_ = _0367_ | _0348_;
	assign _0369_ = _1981_ & ~_0365_;
	assign _0370_ = _1983_ & ~_0364_;
	assign _0371_ = _0370_ | _0369_;
	assign _0372_ = _0371_ | _0368_;
	assign _0373_ = _0372_ | _0345_;
	assign _0374_ = _0334_ | _0285_;
	assign _0375_ = _0374_ | _0274_;
	assign _0376_ = _0175_ & ~_0375_;
	assign _0377_ = _0333_ & ~_1788_;
	assign _0378_ = _0327_ & ~_0334_;
	assign _0379_ = _0378_ | _0377_;
	assign _0380_ = _0278_ & ~_0374_;
	assign _0381_ = _0380_ | _0379_;
	assign _0382_ = _0381_ | _0376_;
	assign _0383_ = ~_0363_;
	assign _0384_ = _0316_ | _0263_;
	assign _0385_ = _0384_ | _0281_;
	assign _0386_ = _0178_ & ~_0385_;
	assign _0387_ = _0386_ ^ _0363_;
	assign _0388_ = (_0062_ ? _0383_ : _0387_);
	assign _0389_ = _0388_ ^ _1848_;
	assign _0390_ = ~(_0389_ ^ _0382_);
	assign \mchip.cpu.alu_result [8] = (_1992_ ? _0373_ : _0390_);
	assign _0391_ = (_1589_ ? _1848_ : _1829_);
	assign _0392_ = (_1622_ ? _0391_ : _0287_);
	assign _0393_ = (_1650_ ? _0184_ : _0392_);
	assign _0394_ = (_1674_ ? _1995_ : _0393_);
	assign _0395_ = _0394_ | _1698_;
	assign _0396_ = _1599_ & ~_0395_;
	assign _0397_ = _2012_ | _1674_;
	assign _0398_ = _0397_ | _1698_;
	assign _0399_ = _1702_ & ~_0398_;
	assign _0400_ = _0399_ | _0396_;
	assign _0401_ = (_1674_ ? _1945_ : _2018_);
	assign _0402_ = (_1698_ ? _1945_ : _0401_);
	assign _0403_ = _1973_ & ~_0402_;
	assign _0404_ = (_1571_ ? _1812_ : _1813_);
	assign _0405_ = (_1571_ ? _1815_ : _1816_);
	assign _0406_ = (_1572_ ? _0404_ : _0405_);
	assign _0407_ = (_1571_ ? _1819_ : _1820_);
	assign _0408_ = (_1571_ ? _1822_ : _1823_);
	assign _0409_ = (_1572_ ? _0407_ : _0408_);
	assign _0410_ = (_1570_ ? _0406_ : _0409_);
	assign _0411_ = _0410_ | _1574_;
	assign _0412_ = ~_0411_;
	assign _0413_ = \mchip.cpu.instr_shift.imm [9] & ~_1461_;
	assign _0414_ = (_1448_ ? \mchip.cpu.instr_shift.imm [9] : _0412_);
	assign _0415_ = (_1441_ ? \mchip.cpu.instr_shift.imm [9] : _0414_);
	assign _0416_ = _0415_ & ~_1427_;
	assign _0417_ = _0416_ | _0413_;
	assign _0418_ = (_1567_ ? _0412_ : _0417_);
	assign _0419_ = _1829_ | ~_0418_;
	assign _0420_ = _1829_ & ~_0418_;
	assign _0421_ = _0420_ | ~_0419_;
	assign _0422_ = _1978_ & ~_0421_;
	assign _0423_ = _0422_ | _0403_;
	assign _0424_ = _1981_ & ~_0420_;
	assign _0425_ = _1983_ & ~_0419_;
	assign _0426_ = _0425_ | _0424_;
	assign _0427_ = _0426_ | _0423_;
	assign _0428_ = _0427_ | _0400_;
	assign _0429_ = _0388_ & ~_1848_;
	assign _0430_ = _0382_ & ~_0389_;
	assign _0431_ = ~(_0430_ | _0429_);
	assign _0432_ = _0363_ | ~_0386_;
	assign _0433_ = _0432_ ^ _0418_;
	assign _0434_ = (_0062_ ? _0418_ : _0433_);
	assign _0435_ = ~(_0434_ ^ _1829_);
	assign _0436_ = _0435_ ^ _0431_;
	assign \mchip.cpu.alu_result [9] = (_1992_ ? _0428_ : _0436_);
	assign _0437_ = (_1589_ ? _1829_ : _1886_);
	assign _0438_ = (_1622_ ? _0437_ : _0336_);
	assign _0439_ = (_1650_ ? _0234_ : _0438_);
	assign _0440_ = (_1674_ ? _0068_ : _0439_);
	assign _0441_ = _0440_ | _1698_;
	assign _0442_ = _1599_ & ~_0441_;
	assign _0443_ = _0077_ | _1674_;
	assign _0444_ = _0443_ | _1698_;
	assign _0445_ = _1702_ & ~_0444_;
	assign _0446_ = _0445_ | _0442_;
	assign _0447_ = (_1674_ ? _1945_ : _0083_);
	assign _0448_ = (_1698_ ? _1945_ : _0447_);
	assign _0449_ = _1973_ & ~_0448_;
	assign _0450_ = (_1571_ ? _1869_ : _1870_);
	assign _0451_ = (_1571_ ? _1872_ : _1873_);
	assign _0452_ = (_1572_ ? _0450_ : _0451_);
	assign _0453_ = (_1571_ ? _1876_ : _1877_);
	assign _0454_ = (_1571_ ? _1879_ : _1880_);
	assign _0455_ = (_1572_ ? _0453_ : _0454_);
	assign _0456_ = (_1570_ ? _0452_ : _0455_);
	assign _0457_ = ~(_0456_ | _1574_);
	assign _0458_ = ~_0457_;
	assign _0459_ = \mchip.cpu.instr_shift.imm [10] & ~_1461_;
	assign _0460_ = (_1448_ ? \mchip.cpu.instr_shift.imm [10] : _0457_);
	assign _0461_ = (_1441_ ? \mchip.cpu.instr_shift.imm [10] : _0460_);
	assign _0462_ = _0461_ & ~_1427_;
	assign _0463_ = ~(_0462_ | _0459_);
	assign _0464_ = (_1567_ ? _0458_ : _0463_);
	assign _0465_ = _0464_ | _1886_;
	assign _0466_ = _0464_ & _1886_;
	assign _0467_ = _0466_ | ~_0465_;
	assign _0468_ = _1978_ & ~_0467_;
	assign _0469_ = _0468_ | _0449_;
	assign _0470_ = _1981_ & ~_0466_;
	assign _0471_ = _1983_ & ~_0465_;
	assign _0472_ = _0471_ | _0470_;
	assign _0473_ = _0472_ | _0469_;
	assign _0474_ = _0473_ | _0446_;
	assign _0475_ = _0435_ | _0389_;
	assign _0476_ = _0382_ & ~_0475_;
	assign _0477_ = ~(_0434_ | _1829_);
	assign _0478_ = _0429_ & ~_0435_;
	assign _0479_ = _0478_ | _0477_;
	assign _0480_ = _0479_ | _0476_;
	assign _0481_ = ~_0464_;
	assign _0482_ = _0418_ | _0363_;
	assign _0483_ = _0386_ & ~_0482_;
	assign _0484_ = _0483_ ^ _0481_;
	assign _0485_ = (_0062_ ? _0464_ : _0484_);
	assign _0486_ = _0485_ ^ _1886_;
	assign _0487_ = ~(_0486_ ^ _0480_);
	assign \mchip.cpu.alu_result [10] = (_1992_ ? _0474_ : _0487_);
	assign _0488_ = (_1589_ ? _1886_ : _1867_);
	assign _0489_ = (_1622_ ? _0488_ : _0391_);
	assign _0490_ = (_1650_ ? _0288_ : _0489_);
	assign _0491_ = (_1674_ ? _0108_ : _0490_);
	assign _0492_ = _0491_ | _1698_;
	assign _0493_ = _1599_ & ~_0492_;
	assign _0494_ = _0117_ | _1674_;
	assign _0495_ = _0494_ | _1698_;
	assign _0496_ = _1702_ & ~_0495_;
	assign _0497_ = _0496_ | _0493_;
	assign _0498_ = (_1674_ ? _1945_ : _0122_);
	assign _0499_ = (_1698_ ? _1945_ : _0498_);
	assign _0500_ = _1973_ & ~_0499_;
	assign _0501_ = (_1571_ ? _1851_ : _1852_);
	assign _0502_ = (_1571_ ? _1854_ : _1855_);
	assign _0503_ = (_1572_ ? _0501_ : _0502_);
	assign _0504_ = (_1571_ ? _1858_ : _1859_);
	assign _0505_ = (_1571_ ? _1861_ : _1862_);
	assign _0506_ = (_1572_ ? _0504_ : _0505_);
	assign _0507_ = (_1570_ ? _0503_ : _0506_);
	assign _0508_ = ~(_0507_ | _1574_);
	assign _0509_ = \mchip.cpu.instr_shift.imm [11] & ~_1461_;
	assign _0510_ = (_1448_ ? \mchip.cpu.instr_shift.imm [11] : _0508_);
	assign _0511_ = (_1441_ ? \mchip.cpu.instr_shift.imm [11] : _0510_);
	assign _0512_ = _0511_ & ~_1427_;
	assign _0513_ = ~(_0512_ | _0509_);
	assign _0514_ = ~_0513_;
	assign _0515_ = (_1567_ ? _0508_ : _0514_);
	assign _0516_ = _1867_ | ~_0515_;
	assign _0517_ = _1867_ & ~_0515_;
	assign _0518_ = _0517_ | ~_0516_;
	assign _0519_ = _1978_ & ~_0518_;
	assign _0520_ = _0519_ | _0500_;
	assign _0521_ = _1981_ & ~_0517_;
	assign _0522_ = _1983_ & ~_0516_;
	assign _0523_ = _0522_ | _0521_;
	assign _0524_ = _0523_ | _0520_;
	assign _0525_ = _0524_ | _0497_;
	assign _0526_ = _0485_ & ~_1886_;
	assign _0527_ = _0480_ & ~_0486_;
	assign _0528_ = ~(_0527_ | _0526_);
	assign _0529_ = ~_0515_;
	assign _0530_ = _0483_ & ~_0481_;
	assign _0531_ = _0530_ ^ _0515_;
	assign _0532_ = (_0062_ ? _0529_ : _0531_);
	assign _0533_ = _0532_ ^ _1867_;
	assign _0534_ = _0533_ ^ _0528_;
	assign \mchip.cpu.alu_result [11] = (_1992_ ? _0525_ : _0534_);
	assign _0535_ = (_1589_ ? _1867_ : _1925_);
	assign _0536_ = (_1622_ ? _0535_ : _0437_);
	assign _0537_ = (_1650_ ? _0337_ : _0536_);
	assign _0538_ = (_1674_ ? _0146_ : _0537_);
	assign _0539_ = _0538_ | _1698_;
	assign _0540_ = _1599_ & ~_0539_;
	assign _0541_ = _0151_ | _1674_;
	assign _0542_ = _0541_ | _1698_;
	assign _0543_ = _1702_ & ~_0542_;
	assign _0544_ = _0543_ | _0540_;
	assign _0545_ = (_1674_ ? _1945_ : _0156_);
	assign _0546_ = (_1698_ ? _1945_ : _0545_);
	assign _0547_ = _1973_ & ~_0546_;
	assign _0548_ = (_1571_ ? _1908_ : _1909_);
	assign _0549_ = (_1571_ ? _1911_ : _1912_);
	assign _0550_ = (_1572_ ? _0548_ : _0549_);
	assign _0551_ = (_1571_ ? _1915_ : _1916_);
	assign _0552_ = (_1571_ ? _1918_ : _1919_);
	assign _0553_ = (_1572_ ? _0551_ : _0552_);
	assign _0554_ = (_1570_ ? _0550_ : _0553_);
	assign _0555_ = ~(_0554_ | _1574_);
	assign _0556_ = \mchip.cpu.instr_shift.imm [12] & ~_1461_;
	assign _0557_ = (_1448_ ? \mchip.cpu.instr_shift.imm [12] : _0555_);
	assign _0558_ = (_1441_ ? \mchip.cpu.instr_shift.imm [12] : _0557_);
	assign _0559_ = _0558_ & ~_1427_;
	assign _0560_ = _0559_ | _0556_;
	assign _0561_ = (_1567_ ? _0555_ : _0560_);
	assign _0562_ = _1925_ | ~_0561_;
	assign _0563_ = _1925_ & ~_0561_;
	assign _0564_ = _0563_ | ~_0562_;
	assign _0565_ = _1978_ & ~_0564_;
	assign _0566_ = _0565_ | _0547_;
	assign _0567_ = _1981_ & ~_0563_;
	assign _0568_ = _1983_ & ~_0562_;
	assign _0569_ = _0568_ | _0567_;
	assign _0570_ = _0569_ | _0566_;
	assign _0571_ = _0570_ | _0544_;
	assign _0572_ = _0532_ & ~_1867_;
	assign _0573_ = _0526_ & ~_0533_;
	assign _0574_ = _0573_ | _0572_;
	assign _0575_ = _0533_ | _0486_;
	assign _0576_ = _0479_ & ~_0575_;
	assign _0577_ = _0576_ | _0574_;
	assign _0578_ = _0575_ | _0475_;
	assign _0579_ = _0382_ & ~_0578_;
	assign _0580_ = _0579_ | _0577_;
	assign _0581_ = _0515_ | _0481_;
	assign _0582_ = _0581_ | _0482_;
	assign _0583_ = _0582_ | ~_0386_;
	assign _0584_ = _0583_ ^ _0561_;
	assign _0585_ = (_0062_ ? _0561_ : _0584_);
	assign _0586_ = _0585_ ^ _1925_;
	assign _0587_ = _0586_ ^ _0580_;
	assign \mchip.cpu.alu_result [12] = (_1992_ ? _0571_ : _0587_);
	assign _0588_ = (_1589_ ? _1925_ : _1906_);
	assign _0589_ = (_1622_ ? _0588_ : _0488_);
	assign _0590_ = (_1650_ ? _0392_ : _0589_);
	assign _0591_ = (_1674_ ? _0185_ : _0590_);
	assign _0592_ = _0591_ | _1698_;
	assign _0593_ = _1599_ & ~_0592_;
	assign _0594_ = _0190_ | _1674_;
	assign _0595_ = _0594_ | _1698_;
	assign _0596_ = _1702_ & ~_0595_;
	assign _0597_ = _0596_ | _0593_;
	assign _0598_ = (_1674_ ? _1945_ : _0195_);
	assign _0599_ = (_1698_ ? _1945_ : _0598_);
	assign _0600_ = _1973_ & ~_0599_;
	assign _0601_ = (_1571_ ? _1890_ : _1891_);
	assign _0602_ = (_1571_ ? _1893_ : _1894_);
	assign _0603_ = (_1572_ ? _0601_ : _0602_);
	assign _0604_ = (_1571_ ? _1897_ : _1898_);
	assign _0605_ = (_1571_ ? _1900_ : _1901_);
	assign _0606_ = (_1572_ ? _0604_ : _0605_);
	assign _0607_ = (_1570_ ? _0603_ : _0606_);
	assign _0608_ = ~(_0607_ | _1574_);
	assign _0609_ = \mchip.cpu.instr_shift.imm [13] & ~_1461_;
	assign _0610_ = (_1448_ ? \mchip.cpu.instr_shift.imm [13] : _0608_);
	assign _0611_ = (_1441_ ? \mchip.cpu.instr_shift.imm [13] : _0610_);
	assign _0612_ = _0611_ & ~_1427_;
	assign _0613_ = _0612_ | _0609_;
	assign _0614_ = (_1567_ ? _0608_ : _0613_);
	assign _0615_ = _1906_ | ~_0614_;
	assign _0616_ = _1906_ & ~_0614_;
	assign _0617_ = _0616_ | ~_0615_;
	assign _0618_ = _1978_ & ~_0617_;
	assign _0619_ = _0618_ | _0600_;
	assign _0620_ = _1981_ & ~_0616_;
	assign _0621_ = _1983_ & ~_0615_;
	assign _0622_ = _0621_ | _0620_;
	assign _0623_ = _0622_ | _0619_;
	assign _0624_ = _0623_ | _0597_;
	assign _0625_ = ~(_0585_ | _1925_);
	assign _0626_ = ~_0586_;
	assign _0627_ = _0580_ & ~_0626_;
	assign _0628_ = ~(_0627_ | _0625_);
	assign _0629_ = _0583_ | _0561_;
	assign _0630_ = _0614_ ^ _0629_;
	assign _0631_ = (_0062_ ? _0614_ : _0630_);
	assign _0632_ = ~(_0631_ ^ _1906_);
	assign _0633_ = _0632_ ^ _0628_;
	assign \mchip.cpu.alu_result [13] = (_1992_ ? _0624_ : _0633_);
	assign _0634_ = (_1589_ ? _1906_ : _1964_);
	assign _0635_ = (_1622_ ? _0634_ : _0535_);
	assign _0636_ = (_1650_ ? _0438_ : _0635_);
	assign _0637_ = (_1674_ ? _0235_ : _0636_);
	assign _0638_ = _0637_ | _1698_;
	assign _0639_ = _1599_ & ~_0638_;
	assign _0640_ = _0240_ | _1674_;
	assign _0641_ = _0640_ | _1698_;
	assign _0642_ = _1702_ & ~_0641_;
	assign _0643_ = _0642_ | _0639_;
	assign _0644_ = (_1674_ ? _1945_ : _0245_);
	assign _0645_ = (_1698_ ? _1945_ : _0644_);
	assign _0646_ = _1973_ & ~_0645_;
	assign _0647_ = (_1571_ ? _1947_ : _1948_);
	assign _0648_ = (_1571_ ? _1950_ : _1951_);
	assign _0649_ = (_1572_ ? _0647_ : _0648_);
	assign _0650_ = (_1571_ ? _1954_ : _1955_);
	assign _0651_ = (_1571_ ? _1957_ : _1958_);
	assign _0652_ = (_1572_ ? _0650_ : _0651_);
	assign _0653_ = (_1570_ ? _0649_ : _0652_);
	assign _0654_ = ~(_0653_ | _1574_);
	assign _0655_ = \mchip.cpu.instr_shift.imm [14] & ~_1461_;
	assign _0656_ = (_1448_ ? \mchip.cpu.instr_shift.imm [14] : _0654_);
	assign _0657_ = (_1441_ ? \mchip.cpu.instr_shift.imm [14] : _0656_);
	assign _0658_ = _0657_ & ~_1427_;
	assign _0659_ = _0658_ | _0655_;
	assign _0660_ = (_1567_ ? _0654_ : _0659_);
	assign _0661_ = _1964_ | ~_0660_;
	assign _0662_ = _1964_ & ~_0660_;
	assign _0663_ = _0662_ | ~_0661_;
	assign _0664_ = _1978_ & ~_0663_;
	assign _0665_ = _0664_ | _0646_;
	assign _0666_ = _1981_ & ~_0662_;
	assign _0667_ = _1983_ & ~_0661_;
	assign _0668_ = _0667_ | _0666_;
	assign _0669_ = _0668_ | _0665_;
	assign _0670_ = _0669_ | _0643_;
	assign _0671_ = ~(_0631_ | _1906_);
	assign _0672_ = _0625_ & ~_0632_;
	assign _0673_ = _0672_ | _0671_;
	assign _0674_ = _0632_ | _0626_;
	assign _0675_ = _0580_ & ~_0674_;
	assign _0676_ = _0675_ | _0673_;
	assign _0677_ = _0614_ | _0561_;
	assign _0678_ = _0677_ | _0583_;
	assign _0679_ = _0678_ ^ _0660_;
	assign _0680_ = (_0062_ ? _0660_ : _0679_);
	assign _0681_ = _0680_ ^ _1964_;
	assign _0682_ = _0681_ ^ _0676_;
	assign \mchip.cpu.alu_result [14] = (_1992_ ? _0670_ : _0682_);
	assign _0683_ = (_1589_ ? _1964_ : _1945_);
	assign _0684_ = (_1622_ ? _0683_ : _0588_);
	assign _0685_ = (_1650_ ? _0489_ : _0684_);
	assign _0686_ = (_1674_ ? _0289_ : _0685_);
	assign _0687_ = _0686_ | _1698_;
	assign _0688_ = _1599_ & ~_0687_;
	assign _0689_ = _0294_ | _1674_;
	assign _0690_ = _0689_ | _1698_;
	assign _0691_ = _1702_ & ~_0690_;
	assign _0692_ = _0691_ | _0688_;
	assign _0693_ = _1973_ & ~_1945_;
	assign _0694_ = (_1571_ ? _1928_ : _1929_);
	assign _0695_ = (_1571_ ? _1931_ : _1932_);
	assign _0696_ = (_1572_ ? _0694_ : _0695_);
	assign _0697_ = (_1571_ ? _1935_ : _1936_);
	assign _0698_ = (_1571_ ? _1938_ : _1939_);
	assign _0699_ = (_1572_ ? _0697_ : _0698_);
	assign _0700_ = (_1570_ ? _0696_ : _0699_);
	assign _0701_ = ~(_0700_ | _1574_);
	assign _0702_ = \mchip.cpu.instr_shift.imm [15] & ~_1461_;
	assign _0703_ = (_1448_ ? \mchip.cpu.instr_shift.imm [15] : _0701_);
	assign _0704_ = (_1441_ ? \mchip.cpu.instr_shift.imm [15] : _0703_);
	assign _0705_ = _0704_ & ~_1427_;
	assign _0706_ = _0705_ | _0702_;
	assign _0707_ = (_1567_ ? _0701_ : _0706_);
	assign _0708_ = _1945_ | ~_0707_;
	assign _0709_ = _1945_ & ~_0707_;
	assign _0710_ = _0709_ | ~_0708_;
	assign _0711_ = _1978_ & ~_0710_;
	assign _0712_ = _0711_ | _0693_;
	assign _0713_ = _1981_ & ~_0709_;
	assign _0714_ = _1983_ & ~_0708_;
	assign _0715_ = _0714_ | _0713_;
	assign _0716_ = _0715_ | _0712_;
	assign _0717_ = _0716_ | _0692_;
	assign _0718_ = ~(_0680_ | _1964_);
	assign _0719_ = _0681_ & _0676_;
	assign _0720_ = _0719_ | _0718_;
	assign _0721_ = _0678_ | _0660_;
	assign _0722_ = _0707_ ^ _0721_;
	assign _0723_ = (_0062_ ? _0707_ : _0722_);
	assign _0724_ = _0723_ ^ _1945_;
	assign _0725_ = _0724_ ^ _0720_;
	assign \mchip.cpu.alu_result [15] = (_1992_ ? _0717_ : _0725_);
	assign _0726_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [0] : \mchip.cpu.alu_result [0]);
	assign \mchip.cpu.rf.rd_data [0] = (_1427_ ? \mchip.cpu.alu_result [0] : _0726_);
	assign _0727_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [1] : \mchip.cpu.alu_result [1]);
	assign \mchip.cpu.rf.rd_data [1] = (_1427_ ? \mchip.cpu.alu_result [1] : _0727_);
	assign _0728_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [2] : \mchip.cpu.alu_result [2]);
	assign \mchip.cpu.rf.rd_data [2] = (_1427_ ? \mchip.cpu.alu_result [2] : _0728_);
	assign _0729_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [3] : \mchip.cpu.alu_result [3]);
	assign \mchip.cpu.rf.rd_data [3] = (_1427_ ? \mchip.cpu.alu_result [3] : _0729_);
	assign _0730_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [4] : \mchip.cpu.alu_result [4]);
	assign \mchip.cpu.rf.rd_data [4] = (_1427_ ? \mchip.cpu.alu_result [4] : _0730_);
	assign _0731_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [5] : \mchip.cpu.alu_result [5]);
	assign \mchip.cpu.rf.rd_data [5] = (_1427_ ? \mchip.cpu.alu_result [5] : _0731_);
	assign _0732_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [6] : \mchip.cpu.alu_result [6]);
	assign \mchip.cpu.rf.rd_data [6] = (_1427_ ? \mchip.cpu.alu_result [6] : _0732_);
	assign _0733_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [7] : \mchip.cpu.alu_result [7]);
	assign \mchip.cpu.rf.rd_data [7] = (_1427_ ? \mchip.cpu.alu_result [7] : _0733_);
	assign _0734_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [8] : \mchip.cpu.alu_result [8]);
	assign \mchip.cpu.rf.rd_data [8] = (_1427_ ? \mchip.cpu.alu_result [8] : _0734_);
	assign _0735_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [9] : \mchip.cpu.alu_result [9]);
	assign \mchip.cpu.rf.rd_data [9] = (_1427_ ? \mchip.cpu.alu_result [9] : _0735_);
	assign _0736_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [10] : \mchip.cpu.alu_result [10]);
	assign \mchip.cpu.rf.rd_data [10] = (_1427_ ? \mchip.cpu.alu_result [10] : _0736_);
	assign _0737_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [11] : \mchip.cpu.alu_result [11]);
	assign \mchip.cpu.rf.rd_data [11] = (_1427_ ? \mchip.cpu.alu_result [11] : _0737_);
	assign _0738_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [12] : \mchip.cpu.alu_result [12]);
	assign \mchip.cpu.rf.rd_data [12] = (_1427_ ? \mchip.cpu.alu_result [12] : _0738_);
	assign _0739_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [13] : \mchip.cpu.alu_result [13]);
	assign \mchip.cpu.rf.rd_data [13] = (_1427_ ? \mchip.cpu.alu_result [13] : _0739_);
	assign _0740_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [14] : \mchip.cpu.alu_result [14]);
	assign \mchip.cpu.rf.rd_data [14] = (_1427_ ? \mchip.cpu.alu_result [14] : _0740_);
	assign _0741_ = (_1441_ ? \mchip.cpu.mdr_shift_reg.prll_out [15] : \mchip.cpu.alu_result [15]);
	assign \mchip.cpu.rf.rd_data [15] = (_1427_ ? \mchip.cpu.alu_result [15] : _0741_);
	assign _0742_ = (io_in[9] ? io_in[0] : _1583_);
	assign _0031_ = (\mchip.cpu.mar_shift_reg.load  ? _0742_ : io_in[0]);
	assign _0743_ = (io_in[9] ? io_in[1] : _1617_);
	assign _0038_ = (\mchip.cpu.mar_shift_reg.load  ? _0743_ : io_in[1]);
	assign _0744_ = (io_in[9] ? io_in[2] : _1642_);
	assign _0039_ = (\mchip.cpu.mar_shift_reg.load  ? _0744_ : io_in[2]);
	assign _0745_ = (io_in[9] ? io_in[3] : _1668_);
	assign _0040_ = (\mchip.cpu.mar_shift_reg.load  ? _0745_ : io_in[3]);
	assign _0746_ = (io_in[9] ? io_in[4] : _1692_);
	assign _0041_ = (\mchip.cpu.mar_shift_reg.load  ? _0746_ : io_in[4]);
	assign _0747_ = (io_in[9] ? io_in[5] : _0207_);
	assign _0042_ = (\mchip.cpu.mar_shift_reg.load  ? _0747_ : io_in[5]);
	assign _0748_ = (io_in[9] ? io_in[6] : _0257_);
	assign _0043_ = (\mchip.cpu.mar_shift_reg.load  ? _0748_ : io_in[6]);
	assign _0749_ = (io_in[9] ? io_in[7] : _0310_);
	assign _0044_ = (\mchip.cpu.mar_shift_reg.load  ? _0749_ : io_in[7]);
	assign _0750_ = _1506_ & ~_0356_;
	assign _0045_ = (\mchip.cpu.mar_shift_reg.load  ? _0750_ : \mchip.cpu.mdr_shift_reg.prll_out [0]);
	assign _0751_ = _1506_ & ~_0411_;
	assign _0046_ = (\mchip.cpu.mar_shift_reg.load  ? _0751_ : \mchip.cpu.mdr_shift_reg.prll_out [1]);
	assign _0752_ = _0457_ & ~io_in[9];
	assign _0032_ = (\mchip.cpu.mar_shift_reg.load  ? _0752_ : \mchip.cpu.mdr_shift_reg.prll_out [2]);
	assign _0753_ = _0508_ & ~io_in[9];
	assign _0033_ = (\mchip.cpu.mar_shift_reg.load  ? _0753_ : \mchip.cpu.mdr_shift_reg.prll_out [3]);
	assign _0754_ = _0555_ & ~io_in[9];
	assign _0034_ = (\mchip.cpu.mar_shift_reg.load  ? _0754_ : \mchip.cpu.mdr_shift_reg.prll_out [4]);
	assign _0755_ = _0608_ & ~io_in[9];
	assign _0035_ = (\mchip.cpu.mar_shift_reg.load  ? _0755_ : \mchip.cpu.mdr_shift_reg.prll_out [5]);
	assign _0756_ = _0654_ & ~io_in[9];
	assign _0036_ = (\mchip.cpu.mar_shift_reg.load  ? _0756_ : \mchip.cpu.mdr_shift_reg.prll_out [6]);
	assign _0757_ = _0701_ & ~io_in[9];
	assign _0037_ = (\mchip.cpu.mar_shift_reg.load  ? _0757_ : \mchip.cpu.mdr_shift_reg.prll_out [7]);
	assign _0758_ = ~\mchip.cpu.pc_reg.prll_out [0];
	assign _0759_ = _1468_ & ~\mchip.cpu.instr_shift.instruction [2];
	assign _0760_ = \mchip.cpu.instr_shift.instruction [2] | ~\mchip.cpu.instr_shift.instruction [1];
	assign _0761_ = ~(_0759_ & \mchip.cpu.instr_shift.instruction [9]);
	assign _0762_ = _1564_ & \mchip.cpu.instr_shift.instruction [4];
	assign _0763_ = _0761_ & ~_0762_;
	assign _0764_ = _0763_ | _0760_;
	assign _0765_ = _0764_ ^ \mchip.cpu.pc_reg.prll_out [0];
	assign _0766_ = _0701_ ^ _1943_;
	assign _0767_ = _0654_ | ~_1962_;
	assign _0768_ = _0767_ | _0766_;
	assign _0769_ = _1943_ & ~_0701_;
	assign _0770_ = _0768_ & ~_0769_;
	assign _0771_ = ~(_0654_ ^ _1962_);
	assign _0772_ = _0771_ & ~_0766_;
	assign _0773_ = _0608_ | _1905_;
	assign _0774_ = ~(_0608_ ^ _1905_);
	assign _0775_ = _1923_ & ~_0555_;
	assign _0776_ = _0775_ & ~_0774_;
	assign _0777_ = _0773_ & ~_0776_;
	assign _0778_ = _0772_ & ~_0777_;
	assign _0779_ = _0770_ & ~_0778_;
	assign _0780_ = _0555_ ^ _1923_;
	assign _0781_ = _0780_ | _0774_;
	assign _0782_ = _0772_ & ~_0781_;
	assign _0783_ = _0508_ | _1866_;
	assign _0784_ = _0508_ ^ _1866_;
	assign _0785_ = _0457_ | ~_1884_;
	assign _0786_ = _0784_ & ~_0785_;
	assign _0787_ = _0783_ & ~_0786_;
	assign _0788_ = _0457_ ^ _1884_;
	assign _0789_ = _0784_ & ~_0788_;
	assign _0790_ = ~(_0411_ & _1827_);
	assign _0791_ = _0356_ & _1846_;
	assign _0792_ = ~(_0411_ ^ _1827_);
	assign _0793_ = _0791_ & ~_0792_;
	assign _0794_ = _0790_ & ~_0793_;
	assign _0795_ = _0789_ & ~_0794_;
	assign _0796_ = _0787_ & ~_0795_;
	assign _0797_ = _0782_ & ~_0796_;
	assign _0798_ = _0779_ & ~_0797_;
	assign _0799_ = _0309_ & _1786_;
	assign _0800_ = _0309_ ^ _1786_;
	assign _0801_ = ~(_0256_ & _1805_);
	assign _0802_ = _0800_ & ~_0801_;
	assign _0803_ = _0802_ | _0799_;
	assign _0804_ = ~(_0256_ ^ _1805_);
	assign _0805_ = _0800_ & ~_0804_;
	assign _0806_ = ~(_0206_ & _1755_);
	assign _0807_ = _1766_ & _1691_;
	assign _0808_ = ~(_0206_ ^ _1755_);
	assign _0809_ = _0807_ & ~_0808_;
	assign _0810_ = _0806_ & ~_0809_;
	assign _0811_ = _0805_ & ~_0810_;
	assign _0812_ = _0811_ | _0803_;
	assign _0813_ = _1723_ & _1667_;
	assign _0814_ = ~(_1723_ ^ _1667_);
	assign _0815_ = _1734_ & _1641_;
	assign _0816_ = _0815_ & ~_0814_;
	assign _0817_ = _0816_ | _0813_;
	assign _0818_ = _1711_ & _1615_;
	assign _0819_ = _1582_ | _1562_;
	assign _0820_ = ~(_1711_ ^ _1615_);
	assign _0821_ = _0819_ & ~_0820_;
	assign _0822_ = _0821_ | _0818_;
	assign _0823_ = ~(_1734_ ^ _1641_);
	assign _0824_ = _0823_ | _0814_;
	assign _0825_ = _0822_ & ~_0824_;
	assign _0826_ = _0825_ | _0817_;
	assign _0827_ = ~(_1766_ ^ _1691_);
	assign _0828_ = ~(_0827_ | _0808_);
	assign _0829_ = ~(_0828_ & _0805_);
	assign _0830_ = _0826_ & ~_0829_;
	assign _0831_ = _0830_ | _0812_;
	assign _0832_ = ~(_0356_ ^ _1846_);
	assign _0833_ = ~(_0832_ | _0792_);
	assign _0834_ = ~(_0833_ & _0789_);
	assign _0835_ = _0834_ | ~_0782_;
	assign _0836_ = _0831_ & ~_0835_;
	assign _0837_ = _0798_ & ~_0836_;
	assign _0838_ = ~(_1582_ ^ _1562_);
	assign _0839_ = _0838_ | _0820_;
	assign _0840_ = _0839_ | _0824_;
	assign _0841_ = _0840_ | _0829_;
	assign _0842_ = ~(_0841_ | _0835_);
	assign _0843_ = _0842_ | ~_0837_;
	assign _0844_ = (_0843_ ? _0765_ : \mchip.cpu.pc_reg.prll_out [0]);
	assign _0845_ = _0759_ & \mchip.cpu.instr_shift.instruction [15];
	assign _0846_ = ~_0845_;
	assign _0847_ = _0759_ & \mchip.cpu.instr_shift.instruction [13];
	assign _0848_ = _0759_ & ~_1432_;
	assign _0849_ = _0848_ | ~_0847_;
	assign _0850_ = _0849_ | _0846_;
	assign _0851_ = _0850_ | _0844_;
	assign _0852_ = _0848_ | _0847_;
	assign _0853_ = _0845_ & ~_0852_;
	assign _0854_ = (_0837_ ? _0765_ : \mchip.cpu.pc_reg.prll_out [0]);
	assign _0855_ = _0853_ & ~_0854_;
	assign _0856_ = _0851_ & ~_0855_;
	assign _0857_ = _0847_ | ~_0848_;
	assign _0858_ = _0846_ & ~_0857_;
	assign _0859_ = _0837_ ^ _0766_;
	assign _0860_ = (_0859_ ? _0765_ : \mchip.cpu.pc_reg.prll_out [0]);
	assign _0861_ = _0858_ & ~_0860_;
	assign _0862_ = ~(_0848_ & _0847_);
	assign _0863_ = _0846_ & ~_0862_;
	assign _0864_ = _0842_ | ~_0859_;
	assign _0865_ = (_0864_ ? _0765_ : \mchip.cpu.pc_reg.prll_out [0]);
	assign _0866_ = _0863_ & ~_0865_;
	assign _0867_ = _0866_ | _0861_;
	assign _0868_ = _0856_ & ~_0867_;
	assign _0869_ = _0846_ & ~_0852_;
	assign _0870_ = (_0842_ ? _0765_ : \mchip.cpu.pc_reg.prll_out [0]);
	assign _0871_ = _0869_ & ~_0870_;
	assign _0872_ = _0846_ & ~_0849_;
	assign _0873_ = (_0842_ ? \mchip.cpu.pc_reg.prll_out [0] : _0765_);
	assign _0874_ = _0872_ & ~_0873_;
	assign _0875_ = _0874_ | _0871_;
	assign _0876_ = _0868_ & ~_0875_;
	assign _0877_ = _0850_ & ~_0853_;
	assign _0878_ = _0863_ | _0858_;
	assign _0879_ = _0877_ & ~_0878_;
	assign _0880_ = _0872_ | _0869_;
	assign _0881_ = _0879_ & ~_0880_;
	assign _0882_ = (_0881_ ? \mchip.cpu.pc_reg.prll_out [0] : _0876_);
	assign _0883_ = _0759_ & ~_0882_;
	assign _0884_ = _0759_ | _1462_;
	assign _0885_ = ~(_0884_ | _1564_);
	assign \mchip.cpu.pc_reg.prll_in [0] = (_0885_ ? _0758_ : _0883_);
	assign _0886_ = \mchip.cpu.pc_reg.prll_out [1] ^ \mchip.cpu.pc_reg.prll_out [0];
	assign _0887_ = ~_0886_;
	assign _0888_ = \mchip.cpu.pc_reg.prll_out [0] & ~_0764_;
	assign _0889_ = ~_0760_;
	assign _0890_ = ~(_1564_ & \mchip.cpu.instr_shift.instruction [5]);
	assign _0891_ = _0759_ & \mchip.cpu.instr_shift.instruction [10];
	assign _0892_ = _0890_ & ~_0891_;
	assign _0893_ = _0889_ & ~_0892_;
	assign _0894_ = _0893_ ^ \mchip.cpu.pc_reg.prll_out [1];
	assign _0895_ = ~(_0894_ ^ _0888_);
	assign _0896_ = (_0843_ ? _0895_ : _0887_);
	assign _0897_ = _0896_ | _0850_;
	assign _0898_ = (_0837_ ? _0895_ : _0887_);
	assign _0899_ = _0853_ & ~_0898_;
	assign _0900_ = _0897_ & ~_0899_;
	assign _0901_ = (_0859_ ? _0895_ : _0887_);
	assign _0902_ = _0858_ & ~_0901_;
	assign _0903_ = (_0864_ ? _0895_ : _0887_);
	assign _0904_ = _0863_ & ~_0903_;
	assign _0905_ = _0904_ | _0902_;
	assign _0906_ = _0900_ & ~_0905_;
	assign _0907_ = (_0842_ ? _0895_ : _0887_);
	assign _0908_ = _0869_ & ~_0907_;
	assign _0909_ = (_0842_ ? _0887_ : _0895_);
	assign _0910_ = _0872_ & ~_0909_;
	assign _0911_ = _0910_ | _0908_;
	assign _0912_ = _0906_ & ~_0911_;
	assign _0913_ = (_0881_ ? _0887_ : _0912_);
	assign _0914_ = _0759_ & ~_0913_;
	assign _0915_ = _1462_ & ~\mchip.cpu.pc_reg.prll_out [1];
	assign _0916_ = _0915_ | _0914_;
	assign \mchip.cpu.pc_reg.prll_in [1] = (_0885_ ? _0886_ : _0916_);
	assign _0917_ = \mchip.cpu.pc_reg.prll_out [1] & \mchip.cpu.pc_reg.prll_out [0];
	assign _0918_ = _0917_ ^ \mchip.cpu.pc_reg.prll_out [2];
	assign _0919_ = ~_0918_;
	assign _0920_ = ~\mchip.cpu.pc_reg.prll_out [1];
	assign _0921_ = _0893_ & ~_0920_;
	assign _0922_ = _0894_ & _0888_;
	assign _0923_ = ~(_0922_ | _0921_);
	assign _0924_ = ~(_1564_ & \mchip.cpu.instr_shift.instruction [6]);
	assign _0925_ = _0759_ & \mchip.cpu.instr_shift.instruction [11];
	assign _0926_ = _0924_ & ~_0925_;
	assign _0927_ = _0889_ & ~_0926_;
	assign _0928_ = _0927_ ^ \mchip.cpu.pc_reg.prll_out [2];
	assign _0929_ = _0928_ ^ _0923_;
	assign _0930_ = (_0843_ ? _0929_ : _0919_);
	assign _0931_ = _0930_ | _0850_;
	assign _0932_ = (_0837_ ? _0929_ : _0919_);
	assign _0933_ = _0853_ & ~_0932_;
	assign _0934_ = _0931_ & ~_0933_;
	assign _0935_ = (_0859_ ? _0929_ : _0919_);
	assign _0936_ = _0858_ & ~_0935_;
	assign _0937_ = (_0864_ ? _0929_ : _0919_);
	assign _0938_ = _0863_ & ~_0937_;
	assign _0939_ = _0938_ | _0936_;
	assign _0940_ = _0934_ & ~_0939_;
	assign _0941_ = (_0842_ ? _0929_ : _0919_);
	assign _0942_ = _0869_ & ~_0941_;
	assign _0943_ = (_0842_ ? _0919_ : _0929_);
	assign _0944_ = _0872_ & ~_0943_;
	assign _0945_ = _0944_ | _0942_;
	assign _0946_ = _0940_ & ~_0945_;
	assign _0947_ = (_0881_ ? _0919_ : _0946_);
	assign _0948_ = _0759_ & ~_0947_;
	assign _0949_ = ~(\mchip.cpu.pc_reg.prll_out [2] ^ \mchip.cpu.pc_reg.prll_out [1]);
	assign _0950_ = _1462_ & ~_0949_;
	assign _0951_ = _0950_ | _0948_;
	assign \mchip.cpu.pc_reg.prll_in [2] = (_0885_ ? _0918_ : _0951_);
	assign _0952_ = _0917_ & ~_1726_;
	assign _0953_ = _0952_ ^ \mchip.cpu.pc_reg.prll_out [3];
	assign _0954_ = ~_0953_;
	assign _0955_ = _0927_ & ~_1726_;
	assign _0956_ = _0923_ | ~_0928_;
	assign _0957_ = _0956_ & ~_0955_;
	assign _0958_ = ~(_1564_ & \mchip.cpu.instr_shift.instruction [7]);
	assign _0959_ = _0759_ & \mchip.cpu.instr_shift.instruction [12];
	assign _0960_ = _0958_ & ~_0959_;
	assign _0961_ = _0889_ & ~_0960_;
	assign _0962_ = _0961_ ^ \mchip.cpu.pc_reg.prll_out [3];
	assign _0963_ = _0962_ ^ _0957_;
	assign _0964_ = (_0843_ ? _0963_ : _0954_);
	assign _0965_ = _0964_ | _0850_;
	assign _0966_ = (_0837_ ? _0963_ : _0954_);
	assign _0967_ = _0853_ & ~_0966_;
	assign _0968_ = _0965_ & ~_0967_;
	assign _0969_ = (_0859_ ? _0963_ : _0954_);
	assign _0970_ = _0858_ & ~_0969_;
	assign _0971_ = (_0864_ ? _0963_ : _0954_);
	assign _0972_ = _0863_ & ~_0971_;
	assign _0973_ = _0972_ | _0970_;
	assign _0974_ = _0968_ & ~_0973_;
	assign _0975_ = (_0842_ ? _0963_ : _0954_);
	assign _0976_ = _0869_ & ~_0975_;
	assign _0977_ = (_0842_ ? _0954_ : _0963_);
	assign _0978_ = _0872_ & ~_0977_;
	assign _0979_ = _0978_ | _0976_;
	assign _0980_ = _0974_ & ~_0979_;
	assign _0981_ = (_0881_ ? _0954_ : _0980_);
	assign _0982_ = _0759_ & ~_0981_;
	assign _0983_ = \mchip.cpu.pc_reg.prll_out [2] & \mchip.cpu.pc_reg.prll_out [1];
	assign _0984_ = _0983_ ^ _1715_;
	assign _0985_ = _1462_ & ~_0984_;
	assign _0986_ = _0985_ | _0982_;
	assign \mchip.cpu.pc_reg.prll_in [3] = (_0885_ ? _0953_ : _0986_);
	assign _0987_ = ~(\mchip.cpu.pc_reg.prll_out [3] & \mchip.cpu.pc_reg.prll_out [2]);
	assign _0988_ = _0917_ & ~_0987_;
	assign _0989_ = _0988_ ^ \mchip.cpu.pc_reg.prll_out [4];
	assign _0990_ = ~_0989_;
	assign _0991_ = ~(_0961_ & \mchip.cpu.pc_reg.prll_out [3]);
	assign _0992_ = _0962_ & _0955_;
	assign _0993_ = _0991_ & ~_0992_;
	assign _0994_ = _0962_ & _0928_;
	assign _0995_ = _0994_ & ~_0923_;
	assign _0996_ = _0993_ & ~_0995_;
	assign _0997_ = _0996_ ^ \mchip.cpu.pc_reg.prll_out [4];
	assign _0998_ = (_0843_ ? _0997_ : _0990_);
	assign _0999_ = _0998_ | _0850_;
	assign _1000_ = (_0837_ ? _0997_ : _0990_);
	assign _1001_ = _0853_ & ~_1000_;
	assign _1002_ = _0999_ & ~_1001_;
	assign _1003_ = (_0859_ ? _0997_ : _0990_);
	assign _1004_ = _0858_ & ~_1003_;
	assign _1005_ = (_0864_ ? _0997_ : _0990_);
	assign _1006_ = _0863_ & ~_1005_;
	assign _1007_ = _1006_ | _1004_;
	assign _1008_ = _1002_ & ~_1007_;
	assign _1009_ = (_0842_ ? _0997_ : _0990_);
	assign _1010_ = _0869_ & ~_1009_;
	assign _1011_ = (_0842_ ? _0990_ : _0997_);
	assign _1012_ = _0872_ & ~_1011_;
	assign _1013_ = _1012_ | _1010_;
	assign _1014_ = _1008_ & ~_1013_;
	assign _1015_ = (_0881_ ? _0990_ : _1014_);
	assign _1016_ = _0759_ & ~_1015_;
	assign _1017_ = _0983_ & ~_1715_;
	assign _1018_ = _1017_ ^ _1758_;
	assign _1019_ = _1462_ & ~_1018_;
	assign _1020_ = _1019_ | _1016_;
	assign \mchip.cpu.pc_reg.prll_in [4] = (_0885_ ? _0989_ : _1020_);
	assign _1021_ = _0988_ & ~_1758_;
	assign _1022_ = _1021_ ^ \mchip.cpu.pc_reg.prll_out [5];
	assign _1023_ = ~_1022_;
	assign _1024_ = \mchip.cpu.pc_reg.prll_out [4] & ~_0996_;
	assign _1025_ = _1024_ ^ _1739_;
	assign _1026_ = (_0843_ ? _1025_ : _1023_);
	assign _1027_ = _1026_ | _0850_;
	assign _1028_ = (_0837_ ? _1025_ : _1023_);
	assign _1029_ = _0853_ & ~_1028_;
	assign _1030_ = _1027_ & ~_1029_;
	assign _1031_ = (_0859_ ? _1025_ : _1023_);
	assign _1032_ = _0858_ & ~_1031_;
	assign _1033_ = (_0864_ ? _1025_ : _1023_);
	assign _1034_ = _0863_ & ~_1033_;
	assign _1035_ = _1034_ | _1032_;
	assign _1036_ = _1030_ & ~_1035_;
	assign _1037_ = (_0842_ ? _1025_ : _1023_);
	assign _1038_ = _0869_ & ~_1037_;
	always @(posedge io_in[10])
		if (_0028_)
			\mchip.cpu.instr_shift.count [0] <= 1'h0;
		else
			\mchip.cpu.instr_shift.count [0] <= _2028_[0];
	always @(posedge io_in[10])
		if (_0028_)
			\mchip.cpu.instr_shift.count [1] <= 1'h0;
		else
			\mchip.cpu.instr_shift.count [1] <= _2029_[1];
	always @(posedge io_in[10])
		if (_0028_)
			\mchip.cpu.instr_shift.count [2] <= 1'h0;
		else
			\mchip.cpu.instr_shift.count [2] <= _2029_[2];
	always @(posedge io_in[10])
		if (_0028_)
			\mchip.cpu.instr_shift.count [3] <= 1'h0;
		else
			\mchip.cpu.instr_shift.count [3] <= _2029_[3];
	always @(posedge io_in[10])
		if (_0028_)
			\mchip.cpu.instr_shift.count [4] <= 1'h0;
		else
			\mchip.cpu.instr_shift.count [4] <= _2029_[4];
	reg \mchip.cpu.ctrl_fsm.cs_reg[0] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[0]  <= _0009_;
	assign \mchip.cpu.ctrl_fsm.cs [0] = \mchip.cpu.ctrl_fsm.cs_reg[0] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[1] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[1]  <= _0002_;
	assign \mchip.cpu.ctrl_fsm.cs [1] = \mchip.cpu.ctrl_fsm.cs_reg[1] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[2] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[2]  <= _0011_;
	assign \mchip.cpu.ctrl_fsm.cs [2] = \mchip.cpu.ctrl_fsm.cs_reg[2] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[3] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[3]  <= _0003_;
	assign \mchip.cpu.ctrl_fsm.cs [3] = \mchip.cpu.ctrl_fsm.cs_reg[3] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[4] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[4]  <= _0004_;
	assign \mchip.cpu.ctrl_fsm.cs [4] = \mchip.cpu.ctrl_fsm.cs_reg[4] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[5] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[5]  <= _0005_;
	assign \mchip.cpu.ctrl_fsm.cs [5] = \mchip.cpu.ctrl_fsm.cs_reg[5] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[6] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[6]  <= _0012_;
	assign \mchip.cpu.ctrl_fsm.cs [6] = \mchip.cpu.ctrl_fsm.cs_reg[6] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[7] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[7]  <= _0013_;
	assign \mchip.cpu.ctrl_fsm.cs [7] = \mchip.cpu.ctrl_fsm.cs_reg[7] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[8] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[8]  <= _0006_;
	assign \mchip.cpu.ctrl_fsm.cs [8] = \mchip.cpu.ctrl_fsm.cs_reg[8] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[9] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[9]  <= _0007_;
	assign \mchip.cpu.ctrl_fsm.cs [9] = \mchip.cpu.ctrl_fsm.cs_reg[9] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[10] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[10]  <= _0008_;
	assign \mchip.cpu.ctrl_fsm.cs [10] = \mchip.cpu.ctrl_fsm.cs_reg[10] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[11] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[11]  <= _0000_;
	assign \mchip.cpu.ctrl_fsm.cs [11] = \mchip.cpu.ctrl_fsm.cs_reg[11] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[12] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[12]  <= _0001_;
	assign \mchip.cpu.ctrl_fsm.cs [12] = \mchip.cpu.ctrl_fsm.cs_reg[12] ;
	reg \mchip.cpu.ctrl_fsm.cs_reg[13] ;
	always @(posedge io_in[10]) \mchip.cpu.ctrl_fsm.cs_reg[13]  <= _0010_;
	assign \mchip.cpu.ctrl_fsm.cs [13] = \mchip.cpu.ctrl_fsm.cs_reg[13] ;
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [0] <= \mchip.cpu.rf.rd_data [0];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [1] <= \mchip.cpu.rf.rd_data [1];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [2] <= \mchip.cpu.rf.rd_data [2];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [3] <= \mchip.cpu.rf.rd_data [3];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [4] <= \mchip.cpu.rf.rd_data [4];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [5] <= \mchip.cpu.rf.rd_data [5];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [6] <= \mchip.cpu.rf.rd_data [6];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [7] <= \mchip.cpu.rf.rd_data [7];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [8] <= \mchip.cpu.rf.rd_data [8];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [9] <= \mchip.cpu.rf.rd_data [9];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [10] <= \mchip.cpu.rf.rd_data [10];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [11] <= \mchip.cpu.rf.rd_data [11];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [12] <= \mchip.cpu.rf.rd_data [12];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [13] <= \mchip.cpu.rf.rd_data [13];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [14] <= \mchip.cpu.rf.rd_data [14];
	always @(posedge io_in[10])
		if (_0048_)
			\mchip.cpu.rf.reg_file[0] [15] <= \mchip.cpu.rf.rd_data [15];
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [0] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [0] <= \mchip.cpu.rf.rd_data [0];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [1] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [1] <= \mchip.cpu.rf.rd_data [1];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [2] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [2] <= \mchip.cpu.rf.rd_data [2];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [3] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [3] <= \mchip.cpu.rf.rd_data [3];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [4] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [4] <= \mchip.cpu.rf.rd_data [4];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [5] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [5] <= \mchip.cpu.rf.rd_data [5];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [6] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [6] <= \mchip.cpu.rf.rd_data [6];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [7] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [7] <= \mchip.cpu.rf.rd_data [7];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [8] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [8] <= \mchip.cpu.rf.rd_data [8];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [9] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [9] <= \mchip.cpu.rf.rd_data [9];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [10] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [10] <= \mchip.cpu.rf.rd_data [10];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [11] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [11] <= \mchip.cpu.rf.rd_data [11];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [12] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [12] <= \mchip.cpu.rf.rd_data [12];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [13] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [13] <= \mchip.cpu.rf.rd_data [13];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [14] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [14] <= \mchip.cpu.rf.rd_data [14];
		end
	always @(posedge io_in[10])
		if (_0020_) begin
			if (!_0050_)
				\mchip.cpu.rf.reg_file[2] [15] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[2] [15] <= \mchip.cpu.rf.rd_data [15];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [0] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [0] <= \mchip.cpu.rf.rd_data [0];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [1] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [1] <= \mchip.cpu.rf.rd_data [1];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [2] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [2] <= \mchip.cpu.rf.rd_data [2];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [3] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [3] <= \mchip.cpu.rf.rd_data [3];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [4] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [4] <= \mchip.cpu.rf.rd_data [4];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [5] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [5] <= \mchip.cpu.rf.rd_data [5];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [6] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [6] <= \mchip.cpu.rf.rd_data [6];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [7] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [7] <= \mchip.cpu.rf.rd_data [7];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [8] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [8] <= \mchip.cpu.rf.rd_data [8];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [9] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [9] <= \mchip.cpu.rf.rd_data [9];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [10] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [10] <= \mchip.cpu.rf.rd_data [10];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [11] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [11] <= \mchip.cpu.rf.rd_data [11];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [12] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [12] <= \mchip.cpu.rf.rd_data [12];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [13] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [13] <= \mchip.cpu.rf.rd_data [13];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [14] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [14] <= \mchip.cpu.rf.rd_data [14];
		end
	always @(posedge io_in[10])
		if (_0018_) begin
			if (!_0052_)
				\mchip.cpu.rf.reg_file[4] [15] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[4] [15] <= \mchip.cpu.rf.rd_data [15];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [0] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [0] <= \mchip.cpu.rf.rd_data [0];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [1] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [1] <= \mchip.cpu.rf.rd_data [1];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [2] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [2] <= \mchip.cpu.rf.rd_data [2];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [3] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [3] <= \mchip.cpu.rf.rd_data [3];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [4] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [4] <= \mchip.cpu.rf.rd_data [4];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [5] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [5] <= \mchip.cpu.rf.rd_data [5];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [6] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [6] <= \mchip.cpu.rf.rd_data [6];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [7] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [7] <= \mchip.cpu.rf.rd_data [7];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [8] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [8] <= \mchip.cpu.rf.rd_data [8];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [9] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [9] <= \mchip.cpu.rf.rd_data [9];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [10] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [10] <= \mchip.cpu.rf.rd_data [10];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [11] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [11] <= \mchip.cpu.rf.rd_data [11];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [12] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [12] <= \mchip.cpu.rf.rd_data [12];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [13] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [13] <= \mchip.cpu.rf.rd_data [13];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [14] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [14] <= \mchip.cpu.rf.rd_data [14];
		end
	always @(posedge io_in[10])
		if (_0019_) begin
			if (!_0051_)
				\mchip.cpu.rf.reg_file[3] [15] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[3] [15] <= \mchip.cpu.rf.rd_data [15];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [0] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [0] <= \mchip.cpu.rf.rd_data [0];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [1] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [1] <= \mchip.cpu.rf.rd_data [1];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [2] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [2] <= \mchip.cpu.rf.rd_data [2];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [3] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [3] <= \mchip.cpu.rf.rd_data [3];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [4] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [4] <= \mchip.cpu.rf.rd_data [4];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [5] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [5] <= \mchip.cpu.rf.rd_data [5];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [6] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [6] <= \mchip.cpu.rf.rd_data [6];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [7] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [7] <= \mchip.cpu.rf.rd_data [7];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [8] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [8] <= \mchip.cpu.rf.rd_data [8];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [9] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [9] <= \mchip.cpu.rf.rd_data [9];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [10] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [10] <= \mchip.cpu.rf.rd_data [10];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [11] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [11] <= \mchip.cpu.rf.rd_data [11];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [12] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [12] <= \mchip.cpu.rf.rd_data [12];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [13] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [13] <= \mchip.cpu.rf.rd_data [13];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [14] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [14] <= \mchip.cpu.rf.rd_data [14];
		end
	always @(posedge io_in[10])
		if (_0015_) begin
			if (!_0055_)
				\mchip.cpu.rf.reg_file[7] [15] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[7] [15] <= \mchip.cpu.rf.rd_data [15];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [0] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [0] <= \mchip.cpu.rf.rd_data [0];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [1] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [1] <= \mchip.cpu.rf.rd_data [1];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [2] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [2] <= \mchip.cpu.rf.rd_data [2];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [3] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [3] <= \mchip.cpu.rf.rd_data [3];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [4] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [4] <= \mchip.cpu.rf.rd_data [4];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [5] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [5] <= \mchip.cpu.rf.rd_data [5];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [6] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [6] <= \mchip.cpu.rf.rd_data [6];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [7] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [7] <= \mchip.cpu.rf.rd_data [7];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [8] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [8] <= \mchip.cpu.rf.rd_data [8];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [9] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [9] <= \mchip.cpu.rf.rd_data [9];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [10] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [10] <= \mchip.cpu.rf.rd_data [10];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [11] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [11] <= \mchip.cpu.rf.rd_data [11];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [12] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [12] <= \mchip.cpu.rf.rd_data [12];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [13] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [13] <= \mchip.cpu.rf.rd_data [13];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [14] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [14] <= \mchip.cpu.rf.rd_data [14];
		end
	always @(posedge io_in[10])
		if (_0016_) begin
			if (!_0054_)
				\mchip.cpu.rf.reg_file[6] [15] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[6] [15] <= \mchip.cpu.rf.rd_data [15];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [0] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [0] <= \mchip.cpu.rf.rd_data [0];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [1] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [1] <= \mchip.cpu.rf.rd_data [1];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [2] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [2] <= \mchip.cpu.rf.rd_data [2];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [3] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [3] <= \mchip.cpu.rf.rd_data [3];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [4] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [4] <= \mchip.cpu.rf.rd_data [4];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [5] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [5] <= \mchip.cpu.rf.rd_data [5];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [6] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [6] <= \mchip.cpu.rf.rd_data [6];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [7] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [7] <= \mchip.cpu.rf.rd_data [7];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [8] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [8] <= \mchip.cpu.rf.rd_data [8];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [9] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [9] <= \mchip.cpu.rf.rd_data [9];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [10] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [10] <= \mchip.cpu.rf.rd_data [10];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [11] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [11] <= \mchip.cpu.rf.rd_data [11];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [12] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [12] <= \mchip.cpu.rf.rd_data [12];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [13] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [13] <= \mchip.cpu.rf.rd_data [13];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [14] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [14] <= \mchip.cpu.rf.rd_data [14];
		end
	always @(posedge io_in[10])
		if (_0021_) begin
			if (!_0049_)
				\mchip.cpu.rf.reg_file[1] [15] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[1] [15] <= \mchip.cpu.rf.rd_data [15];
		end
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [1] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [1] <= \mchip.cpu.pc_reg.prll_in [1];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [2] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [2] <= \mchip.cpu.pc_reg.prll_in [2];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [3] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [3] <= \mchip.cpu.pc_reg.prll_in [3];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [4] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [4] <= \mchip.cpu.pc_reg.prll_in [4];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [5] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [5] <= \mchip.cpu.pc_reg.prll_in [5];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [6] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [6] <= \mchip.cpu.pc_reg.prll_in [6];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [7] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [7] <= \mchip.cpu.pc_reg.prll_in [7];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [8] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [8] <= \mchip.cpu.pc_reg.prll_in [8];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [9] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [9] <= \mchip.cpu.pc_reg.prll_in [9];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [10] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [10] <= \mchip.cpu.pc_reg.prll_in [10];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [11] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [11] <= \mchip.cpu.pc_reg.prll_in [11];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [12] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [12] <= \mchip.cpu.pc_reg.prll_in [12];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [13] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [13] <= \mchip.cpu.pc_reg.prll_in [13];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [14] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [14] <= \mchip.cpu.pc_reg.prll_in [14];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [15] <= 1'h0;
		else if (\mchip.cpu.ctrl_fsm.cs [1])
			\mchip.cpu.pc_reg.prll_out [15] <= \mchip.cpu.pc_reg.prll_in [15];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [0] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [0] <= \mchip.cpu.instr_shift.instruction [8];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [1] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [1] <= \mchip.cpu.instr_shift.instruction [9];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [2] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [2] <= \mchip.cpu.instr_shift.instruction [10];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [3] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [3] <= \mchip.cpu.instr_shift.instruction [11];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [4] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [4] <= \mchip.cpu.instr_shift.instruction [12];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [5] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [5] <= \mchip.cpu.instr_shift.instruction [13];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [6] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [6] <= \mchip.cpu.instr_shift.instruction [14];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [7] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [7] <= \mchip.cpu.instr_shift.instruction [15];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [8] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [8] <= io_in[0];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [9] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [9] <= io_in[1];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [10] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [10] <= io_in[2];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [11] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [11] <= io_in[3];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [12] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [12] <= io_in[4];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [13] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [13] <= io_in[5];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [14] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [14] <= io_in[6];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.instruction [15] <= 1'h0;
		else if (_0025_)
			\mchip.cpu.instr_shift.instruction [15] <= io_in[7];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [0] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [0] <= \mchip.cpu.instr_shift.imm [8];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [1] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [1] <= \mchip.cpu.instr_shift.imm [9];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [2] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [2] <= \mchip.cpu.instr_shift.imm [10];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [3] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [3] <= \mchip.cpu.instr_shift.imm [11];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [4] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [4] <= \mchip.cpu.instr_shift.imm [12];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [5] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [5] <= \mchip.cpu.instr_shift.imm [13];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [6] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [6] <= \mchip.cpu.instr_shift.imm [14];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [7] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [7] <= \mchip.cpu.instr_shift.imm [15];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [8] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [8] <= io_in[0];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [9] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [9] <= io_in[1];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [10] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [10] <= io_in[2];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [11] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [11] <= io_in[3];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [12] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [12] <= io_in[4];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [13] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [13] <= io_in[5];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [14] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [14] <= io_in[6];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.instr_shift.imm [15] <= 1'h0;
		else if (_0026_)
			\mchip.cpu.instr_shift.imm [15] <= io_in[7];
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [0] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [0] <= \mchip.cpu.rf.rd_data [0];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [1] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [1] <= \mchip.cpu.rf.rd_data [1];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [2] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [2] <= \mchip.cpu.rf.rd_data [2];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [3] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [3] <= \mchip.cpu.rf.rd_data [3];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [4] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [4] <= \mchip.cpu.rf.rd_data [4];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [5] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [5] <= \mchip.cpu.rf.rd_data [5];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [6] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [6] <= \mchip.cpu.rf.rd_data [6];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [7] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [7] <= \mchip.cpu.rf.rd_data [7];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [8] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [8] <= \mchip.cpu.rf.rd_data [8];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [9] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [9] <= \mchip.cpu.rf.rd_data [9];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [10] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [10] <= \mchip.cpu.rf.rd_data [10];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [11] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [11] <= \mchip.cpu.rf.rd_data [11];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [12] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [12] <= \mchip.cpu.rf.rd_data [12];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [13] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [13] <= \mchip.cpu.rf.rd_data [13];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [14] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [14] <= \mchip.cpu.rf.rd_data [14];
		end
	always @(posedge io_in[10])
		if (_0017_) begin
			if (!_0053_)
				\mchip.cpu.rf.reg_file[5] [15] <= 1'h0;
			else
				\mchip.cpu.rf.reg_file[5] [15] <= \mchip.cpu.rf.rd_data [15];
		end
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.low_b  <= 1'h1;
		else if (_0022_)
			\mchip.cpu.pc_reg.low_b  <= _0047_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.low_b  <= 1'h1;
		else if (_0023_)
			\mchip.cpu.mdr_shift_reg.low_b  <= _0030_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [0] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [0] <= _0031_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [1] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [1] <= _0038_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [2] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [2] <= _0039_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [3] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [3] <= _0040_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [4] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [4] <= _0041_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [5] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [5] <= _0042_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [6] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [6] <= _0043_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [7] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [7] <= _0044_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [8] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [8] <= _0045_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [9] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [9] <= _0046_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [10] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [10] <= _0032_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [11] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [11] <= _0033_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [12] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [12] <= _0034_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [13] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [13] <= _0035_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [14] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [14] <= _0036_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mdr_shift_reg.prll_out [15] <= 1'h0;
		else if (_0014_)
			\mchip.cpu.mdr_shift_reg.prll_out [15] <= _0037_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.pc_reg.prll_out [0] <= 1'h0;
		else if (_0027_)
			\mchip.cpu.pc_reg.prll_out [0] <= \mchip.cpu.pc_reg.prll_in [0];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.low_b  <= 1'h1;
		else if (_0024_)
			\mchip.cpu.mar_shift_reg.low_b  <= _0029_;
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [0] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [0] <= \mchip.cpu.alu_result [0];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [1] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [1] <= \mchip.cpu.alu_result [1];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [2] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [2] <= \mchip.cpu.alu_result [2];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [3] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [3] <= \mchip.cpu.alu_result [3];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [4] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [4] <= \mchip.cpu.alu_result [4];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [5] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [5] <= \mchip.cpu.alu_result [5];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [6] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [6] <= \mchip.cpu.alu_result [6];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [7] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [7] <= \mchip.cpu.alu_result [7];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [8] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [8] <= \mchip.cpu.alu_result [8];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [9] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [9] <= \mchip.cpu.alu_result [9];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [10] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [10] <= \mchip.cpu.alu_result [10];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [11] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [11] <= \mchip.cpu.alu_result [11];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [12] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [12] <= \mchip.cpu.alu_result [12];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [13] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [13] <= \mchip.cpu.alu_result [13];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [14] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [14] <= \mchip.cpu.alu_result [14];
	always @(posedge io_in[10])
		if (io_in[13])
			\mchip.cpu.mar_shift_reg.prll_out [15] <= 1'h0;
		else if (\mchip.cpu.mar_shift_reg.load )
			\mchip.cpu.mar_shift_reg.prll_out [15] <= \mchip.cpu.alu_result [15];
	assign _2028_[4:1] = 4'h0;
	assign _2029_[0] = _2028_[0];
	assign io_out[13:8] = {2'h0, \mchip.cpu.ctrl_fsm.halt , \mchip.cpu.bus_mdr , \mchip.cpu.bus_mar , \mchip.cpu.bus_pc };
	assign \mchip.clock  = io_in[12];
	assign \mchip.cpu.alu.result  = \mchip.cpu.alu_result ;
	assign \mchip.cpu.ard_clk  = io_in[10];
	assign \mchip.cpu.ard_data_ready  = io_in[9];
	assign \mchip.cpu.ard_receive_ready  = io_in[8];
	assign \mchip.cpu.clk  = io_in[12];
	assign \mchip.cpu.ctrl  = {2'h0, \mchip.cpu.bus_mdr , \mchip.cpu.bus_mar , 1'h0, \mchip.cpu.bus_pc , 1'h0, \mchip.cpu.mar_shift_reg.load , \mchip.cpu.mar_shift_reg.load , \mchip.cpu.ctrl_fsm.cs [1]};
	assign \mchip.cpu.ctrl_fsm.ard_data_ready  = io_in[9];
	assign \mchip.cpu.ctrl_fsm.ard_receive_ready  = io_in[8];
	assign \mchip.cpu.ctrl_fsm.bus_mar  = \mchip.cpu.bus_mar ;
	assign \mchip.cpu.ctrl_fsm.bus_mdr  = \mchip.cpu.bus_mdr ;
	assign \mchip.cpu.ctrl_fsm.bus_pc  = \mchip.cpu.bus_pc ;
	assign \mchip.cpu.ctrl_fsm.clk  = io_in[10];
	assign \mchip.cpu.ctrl_fsm.cs [14] = 1'h0;
	assign \mchip.cpu.ctrl_fsm.ctrl  = {2'h0, \mchip.cpu.bus_mdr , \mchip.cpu.bus_mar , 1'h0, \mchip.cpu.bus_pc , 1'h0, \mchip.cpu.mar_shift_reg.load , \mchip.cpu.mar_shift_reg.load , \mchip.cpu.ctrl_fsm.cs [1]};
	assign \mchip.cpu.ctrl_fsm.rst  = io_in[13];
	assign \mchip.cpu.ctrl_fsm.signals  = {\mchip.cpu.instr_shift.instruction [2:0], 41'h00000000000};
	assign \mchip.cpu.dec  = {\mchip.cpu.instr_shift.instruction [2:0], 41'h00000000000};
	assign \mchip.cpu.dec_instr.instruction  = \mchip.cpu.instr_shift.instruction ;
	assign \mchip.cpu.dec_instr.signals  = {\mchip.cpu.instr_shift.instruction [2:0], 41'h00000000000};
	assign \mchip.cpu.error_instr  = 1'h0;
	assign \mchip.cpu.halt  = \mchip.cpu.ctrl_fsm.halt ;
	assign \mchip.cpu.imm  = \mchip.cpu.instr_shift.imm ;
	assign \mchip.cpu.in_bus  = io_in[7:0];
	assign \mchip.cpu.instr  = \mchip.cpu.instr_shift.instruction ;
	assign \mchip.cpu.instr_shift.clk  = io_in[10];
	assign \mchip.cpu.instr_shift.data_ready  = io_in[9];
	assign \mchip.cpu.instr_shift.error  = 1'h0;
	assign \mchip.cpu.instr_shift.halt  = \mchip.cpu.ctrl_fsm.halt ;
	assign \mchip.cpu.instr_shift.opcode  = \mchip.cpu.instr_shift.instruction [2:0];
	assign \mchip.cpu.instr_shift.rst  = io_in[13];
	assign \mchip.cpu.instr_shift.serial_in  = io_in[7:0];
	assign \mchip.cpu.mar_in  = \mchip.cpu.alu_result ;
	assign \mchip.cpu.mar_out  = \mchip.cpu.mar_shift_reg.prll_out ;
	assign \mchip.cpu.mar_shift_reg.clk  = io_in[10];
	assign \mchip.cpu.mar_shift_reg.prll_in  = \mchip.cpu.alu_result ;
	assign \mchip.cpu.mar_shift_reg.rst  = io_in[13];
	assign \mchip.cpu.mar_shift_reg.serial_in  = 8'h00;
	assign \mchip.cpu.mar_shift_reg.shift_in  = 1'h0;
	assign \mchip.cpu.mar_shift_reg.shift_out  = \mchip.cpu.bus_mar ;
	assign \mchip.cpu.mdr_out  = \mchip.cpu.mdr_shift_reg.prll_out ;
	assign \mchip.cpu.mdr_shift_reg.clk  = io_in[10];
	assign \mchip.cpu.mdr_shift_reg.load  = \mchip.cpu.mar_shift_reg.load ;
	assign \mchip.cpu.mdr_shift_reg.rst  = io_in[13];
	assign \mchip.cpu.mdr_shift_reg.serial_in  = io_in[7:0];
	assign \mchip.cpu.mdr_shift_reg.shift_in  = 1'h0;
	assign \mchip.cpu.mdr_shift_reg.shift_out  = \mchip.cpu.bus_mdr ;
	assign \mchip.cpu.out_bus  = io_out[7:0];
	assign \mchip.cpu.pc  = \mchip.cpu.pc_reg.prll_out ;
	assign \mchip.cpu.pc_in  = \mchip.cpu.pc_reg.prll_in ;
	assign \mchip.cpu.pc_reg.clk  = io_in[10];
	assign \mchip.cpu.pc_reg.load  = \mchip.cpu.ctrl_fsm.cs [1];
	assign \mchip.cpu.pc_reg.rst  = io_in[13];
	assign \mchip.cpu.pc_reg.shift_out  = \mchip.cpu.bus_pc ;
	assign \mchip.cpu.rd_data  = \mchip.cpu.rf.rd_data ;
	assign \mchip.cpu.rf.clk  = io_in[10];
	assign \mchip.cpu.rf.rd  = 3'h0;
	assign \mchip.cpu.rf.rs1  = 3'h0;
	assign \mchip.cpu.rf.rs2  = 3'h0;
	assign \mchip.cpu.rf.rst  = io_in[13];
	assign \mchip.cpu.rst  = io_in[13];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.cpu.ctrl_fsm.halt , \mchip.cpu.bus_mdr , \mchip.cpu.bus_mar , \mchip.cpu.bus_pc , io_out[7:0]};
	assign \mchip.reset  = io_in[13];
endmodule
module d20_zhehuax_16bit_fpu (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	reg _0016_;
	reg _0017_;
	reg _0018_;
	reg _0019_;
	reg _0020_;
	reg _0021_;
	reg _0022_;
	reg _0023_;
	reg _0024_;
	reg _0025_;
	reg _0026_;
	reg _0027_;
	reg _0028_;
	reg _0029_;
	reg _0030_;
	reg _0031_;
	reg _0032_;
	reg _0033_;
	reg _0034_;
	reg _0035_;
	reg _0036_;
	reg _0037_;
	reg _0038_;
	reg _0039_;
	reg _0040_;
	reg _0041_;
	reg _0042_;
	reg _0043_;
	reg _0044_;
	reg _0045_;
	reg _0046_;
	reg _0047_;
	reg _0048_;
	reg _0049_;
	reg _0050_;
	reg _0051_;
	reg _0052_;
	reg _0053_;
	reg _0054_;
	reg _0055_;
	reg _0056_;
	reg _0057_;
	reg _0058_;
	reg _0059_;
	reg _0060_;
	reg _0061_;
	reg _0062_;
	reg _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire _2025_;
	wire _2026_;
	wire _2027_;
	wire _2028_;
	wire _2029_;
	wire _2030_;
	wire _2031_;
	wire _2032_;
	wire _2033_;
	wire _2034_;
	wire _2035_;
	wire _2036_;
	wire _2037_;
	wire _2038_;
	wire _2039_;
	wire _2040_;
	wire _2041_;
	wire _2042_;
	wire _2043_;
	wire _2044_;
	wire _2045_;
	wire _2046_;
	wire _2047_;
	wire _2048_;
	wire _2049_;
	wire _2050_;
	wire _2051_;
	wire _2052_;
	wire _2053_;
	wire _2054_;
	wire _2055_;
	wire _2056_;
	wire _2057_;
	wire _2058_;
	wire _2059_;
	wire _2060_;
	wire _2061_;
	wire _2062_;
	wire _2063_;
	wire _2064_;
	wire _2065_;
	wire _2066_;
	wire _2067_;
	wire _2068_;
	wire _2069_;
	wire _2070_;
	wire _2071_;
	wire _2072_;
	wire _2073_;
	wire _2074_;
	wire _2075_;
	wire _2076_;
	wire _2077_;
	wire _2078_;
	wire _2079_;
	wire _2080_;
	wire _2081_;
	wire _2082_;
	wire _2083_;
	wire _2084_;
	wire _2085_;
	wire _2086_;
	wire _2087_;
	wire _2088_;
	wire _2089_;
	wire _2090_;
	wire _2091_;
	wire _2092_;
	wire _2093_;
	wire _2094_;
	wire _2095_;
	wire _2096_;
	wire _2097_;
	wire _2098_;
	wire _2099_;
	wire _2100_;
	wire _2101_;
	wire _2102_;
	wire _2103_;
	wire _2104_;
	wire _2105_;
	wire _2106_;
	wire _2107_;
	wire _2108_;
	wire _2109_;
	wire _2110_;
	wire _2111_;
	wire _2112_;
	wire _2113_;
	wire _2114_;
	wire _2115_;
	wire _2116_;
	wire _2117_;
	wire _2118_;
	wire _2119_;
	wire _2120_;
	wire _2121_;
	wire _2122_;
	wire _2123_;
	wire _2124_;
	wire _2125_;
	wire _2126_;
	wire _2127_;
	wire _2128_;
	wire _2129_;
	wire _2130_;
	wire _2131_;
	wire _2132_;
	wire _2133_;
	wire _2134_;
	wire _2135_;
	wire _2136_;
	wire _2137_;
	wire _2138_;
	wire _2139_;
	wire _2140_;
	wire _2141_;
	wire _2142_;
	wire _2143_;
	wire _2144_;
	wire _2145_;
	wire _2146_;
	wire _2147_;
	wire _2148_;
	wire _2149_;
	wire _2150_;
	wire _2151_;
	wire _2152_;
	wire _2153_;
	wire _2154_;
	wire _2155_;
	wire _2156_;
	wire _2157_;
	wire _2158_;
	wire _2159_;
	wire _2160_;
	wire _2161_;
	wire _2162_;
	wire _2163_;
	wire _2164_;
	wire _2165_;
	wire _2166_;
	wire _2167_;
	wire _2168_;
	wire _2169_;
	wire _2170_;
	wire _2171_;
	wire _2172_;
	wire _2173_;
	wire _2174_;
	wire _2175_;
	wire _2176_;
	wire _2177_;
	wire _2178_;
	wire _2179_;
	wire _2180_;
	wire _2181_;
	wire _2182_;
	wire _2183_;
	wire _2184_;
	wire _2185_;
	wire _2186_;
	wire _2187_;
	wire _2188_;
	wire _2189_;
	wire _2190_;
	wire _2191_;
	wire _2192_;
	wire _2193_;
	wire _2194_;
	wire _2195_;
	wire _2196_;
	wire _2197_;
	wire _2198_;
	wire _2199_;
	wire _2200_;
	wire _2201_;
	wire _2202_;
	wire _2203_;
	wire _2204_;
	wire _2205_;
	wire _2206_;
	wire _2207_;
	wire _2208_;
	wire _2209_;
	wire _2210_;
	wire _2211_;
	wire _2212_;
	wire _2213_;
	wire _2214_;
	wire _2215_;
	wire _2216_;
	wire _2217_;
	wire _2218_;
	wire _2219_;
	wire _2220_;
	wire _2221_;
	wire _2222_;
	wire _2223_;
	wire _2224_;
	wire _2225_;
	wire _2226_;
	wire _2227_;
	wire _2228_;
	wire _2229_;
	wire _2230_;
	wire _2231_;
	wire _2232_;
	wire _2233_;
	wire _2234_;
	wire _2235_;
	wire _2236_;
	wire _2237_;
	wire _2238_;
	wire _2239_;
	wire _2240_;
	wire _2241_;
	wire _2242_;
	wire _2243_;
	wire _2244_;
	wire _2245_;
	wire _2246_;
	wire _2247_;
	wire _2248_;
	wire _2249_;
	wire _2250_;
	wire _2251_;
	wire _2252_;
	wire _2253_;
	wire _2254_;
	wire _2255_;
	wire _2256_;
	wire _2257_;
	wire _2258_;
	wire _2259_;
	wire _2260_;
	wire _2261_;
	wire _2262_;
	wire _2263_;
	wire _2264_;
	wire _2265_;
	wire _2266_;
	wire _2267_;
	wire _2268_;
	wire _2269_;
	wire _2270_;
	wire _2271_;
	wire _2272_;
	wire _2273_;
	wire _2274_;
	wire _2275_;
	wire _2276_;
	wire _2277_;
	wire _2278_;
	wire _2279_;
	wire _2280_;
	wire _2281_;
	wire _2282_;
	wire _2283_;
	wire _2284_;
	wire _2285_;
	wire _2286_;
	wire _2287_;
	wire _2288_;
	wire _2289_;
	wire _2290_;
	wire _2291_;
	wire _2292_;
	wire _2293_;
	wire _2294_;
	wire _2295_;
	wire _2296_;
	wire _2297_;
	wire _2298_;
	wire _2299_;
	wire _2300_;
	wire _2301_;
	wire _2302_;
	wire _2303_;
	wire _2304_;
	wire _2305_;
	wire _2306_;
	wire _2307_;
	wire _2308_;
	wire _2309_;
	wire _2310_;
	wire _2311_;
	wire _2312_;
	wire _2313_;
	wire _2314_;
	wire _2315_;
	wire _2316_;
	wire _2317_;
	wire _2318_;
	wire _2319_;
	wire _2320_;
	wire _2321_;
	wire _2322_;
	wire _2323_;
	wire _2324_;
	wire _2325_;
	wire _2326_;
	wire _2327_;
	wire _2328_;
	wire _2329_;
	wire _2330_;
	wire _2331_;
	wire _2332_;
	wire _2333_;
	wire _2334_;
	wire _2335_;
	wire _2336_;
	wire _2337_;
	wire _2338_;
	wire _2339_;
	wire _2340_;
	wire _2341_;
	wire _2342_;
	wire _2343_;
	wire _2344_;
	wire _2345_;
	wire _2346_;
	wire _2347_;
	wire _2348_;
	wire _2349_;
	wire _2350_;
	wire _2351_;
	wire _2352_;
	wire _2353_;
	wire _2354_;
	wire _2355_;
	wire _2356_;
	wire _2357_;
	wire _2358_;
	wire _2359_;
	wire _2360_;
	wire _2361_;
	wire _2362_;
	wire _2363_;
	wire _2364_;
	wire _2365_;
	wire _2366_;
	wire _2367_;
	wire _2368_;
	wire _2369_;
	wire _2370_;
	wire _2371_;
	wire _2372_;
	wire _2373_;
	wire _2374_;
	wire _2375_;
	wire _2376_;
	wire _2377_;
	wire _2378_;
	wire _2379_;
	wire _2380_;
	wire _2381_;
	wire _2382_;
	wire _2383_;
	wire _2384_;
	wire _2385_;
	wire _2386_;
	wire _2387_;
	wire _2388_;
	wire _2389_;
	wire _2390_;
	wire _2391_;
	wire _2392_;
	wire _2393_;
	wire _2394_;
	wire _2395_;
	wire _2396_;
	wire _2397_;
	wire _2398_;
	wire _2399_;
	wire _2400_;
	wire _2401_;
	wire _2402_;
	wire _2403_;
	wire _2404_;
	wire _2405_;
	wire _2406_;
	wire _2407_;
	wire _2408_;
	wire _2409_;
	wire _2410_;
	wire _2411_;
	wire _2412_;
	wire _2413_;
	wire _2414_;
	wire _2415_;
	wire _2416_;
	wire _2417_;
	wire _2418_;
	wire _2419_;
	wire _2420_;
	wire _2421_;
	wire _2422_;
	wire _2423_;
	wire _2424_;
	wire _2425_;
	wire _2426_;
	wire _2427_;
	wire _2428_;
	wire _2429_;
	wire _2430_;
	wire _2431_;
	wire _2432_;
	wire _2433_;
	wire _2434_;
	wire _2435_;
	wire _2436_;
	wire _2437_;
	wire _2438_;
	wire _2439_;
	wire _2440_;
	wire _2441_;
	wire _2442_;
	wire _2443_;
	wire _2444_;
	wire _2445_;
	wire _2446_;
	wire _2447_;
	wire _2448_;
	wire _2449_;
	wire _2450_;
	wire _2451_;
	wire _2452_;
	wire _2453_;
	wire _2454_;
	wire _2455_;
	wire _2456_;
	wire _2457_;
	wire _2458_;
	wire _2459_;
	wire _2460_;
	wire _2461_;
	wire _2462_;
	wire _2463_;
	wire _2464_;
	wire _2465_;
	wire _2466_;
	wire _2467_;
	wire _2468_;
	wire _2469_;
	wire _2470_;
	wire _2471_;
	wire _2472_;
	wire _2473_;
	wire _2474_;
	wire _2475_;
	wire _2476_;
	wire _2477_;
	wire _2478_;
	wire _2479_;
	wire _2480_;
	wire _2481_;
	wire _2482_;
	wire _2483_;
	wire _2484_;
	wire _2485_;
	wire _2486_;
	wire _2487_;
	wire _2488_;
	wire _2489_;
	wire _2490_;
	wire _2491_;
	wire _2492_;
	wire _2493_;
	wire _2494_;
	wire _2495_;
	wire _2496_;
	wire _2497_;
	wire _2498_;
	wire _2499_;
	wire _2500_;
	wire _2501_;
	wire _2502_;
	wire _2503_;
	wire _2504_;
	wire _2505_;
	wire _2506_;
	wire _2507_;
	wire _2508_;
	wire _2509_;
	wire _2510_;
	wire _2511_;
	wire _2512_;
	wire _2513_;
	wire _2514_;
	wire _2515_;
	wire _2516_;
	wire _2517_;
	wire _2518_;
	wire _2519_;
	wire _2520_;
	wire _2521_;
	wire _2522_;
	wire _2523_;
	wire _2524_;
	wire _2525_;
	wire _2526_;
	wire _2527_;
	wire _2528_;
	wire _2529_;
	wire _2530_;
	wire _2531_;
	wire _2532_;
	wire _2533_;
	wire _2534_;
	wire _2535_;
	wire _2536_;
	wire _2537_;
	wire _2538_;
	wire _2539_;
	wire _2540_;
	wire _2541_;
	wire _2542_;
	wire _2543_;
	wire _2544_;
	wire _2545_;
	wire _2546_;
	wire _2547_;
	wire _2548_;
	wire _2549_;
	wire _2550_;
	wire _2551_;
	wire _2552_;
	wire _2553_;
	wire _2554_;
	wire _2555_;
	wire _2556_;
	wire _2557_;
	wire _2558_;
	wire _2559_;
	wire _2560_;
	wire _2561_;
	wire _2562_;
	wire _2563_;
	wire _2564_;
	wire _2565_;
	wire _2566_;
	wire _2567_;
	wire _2568_;
	wire _2569_;
	wire _2570_;
	wire _2571_;
	wire _2572_;
	wire _2573_;
	wire _2574_;
	wire _2575_;
	wire _2576_;
	wire _2577_;
	wire _2578_;
	wire _2579_;
	wire _2580_;
	wire _2581_;
	wire _2582_;
	wire _2583_;
	wire _2584_;
	wire _2585_;
	wire _2586_;
	wire _2587_;
	wire _2588_;
	wire _2589_;
	wire _2590_;
	wire _2591_;
	wire _2592_;
	wire _2593_;
	wire _2594_;
	wire _2595_;
	wire _2596_;
	wire _2597_;
	wire _2598_;
	wire _2599_;
	wire _2600_;
	wire _2601_;
	wire _2602_;
	wire _2603_;
	wire _2604_;
	wire _2605_;
	wire _2606_;
	wire _2607_;
	wire _2608_;
	wire _2609_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [15:0] \mchip.calc.b ;
	wire [4:0] \mchip.calc.max_exp ;
	wire [4:0] \mchip.calc.min_exp ;
	wire \mchip.clock ;
	wire \mchip.in1.clock ;
	wire [9:0] \mchip.in1.data_in ;
	wire \mchip.in1.reset ;
	wire \mchip.in1.start ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.out1.clock ;
	wire [9:0] \mchip.out1.data_out ;
	wire \mchip.out1.done_calc ;
	wire \mchip.out1.reset ;
	wire \mchip.reset ;
	wire \mchip.signal ;
	assign _2378_ = io_in[1] & ~io_in[0];
	assign _2389_ = io_in[0] & ~io_in[1];
	assign _0000_ = ~(_2389_ | _2378_);
	assign _2410_ = _0016_ & ~io_in[13];
	assign _0006_ = ~_2410_;
	assign _2431_ = _2410_ | _2389_;
	assign _0002_ = _2378_ & ~_2431_;
	assign _0001_ = io_in[1] & io_in[0];
	assign _2462_ = _2389_ | ~_2410_;
	assign _0003_ = _2378_ & ~_2462_;
	assign _0004_ = _2389_ & ~_2410_;
	assign _0005_ = _2410_ & _2389_;
	assign \mchip.in1.start  = _0063_ & ~io_in[13];
	assign _2523_ = _0042_ & ~io_in[13];
	assign _2533_ = _0018_ & ~io_in[13];
	assign _2544_ = _0017_ & ~io_in[13];
	assign _2555_ = ~(_2544_ | _2533_);
	assign _2566_ = _0058_ & ~io_in[13];
	assign _2577_ = _0057_ & ~io_in[13];
	assign _2588_ = _2577_ | _2566_;
	assign _2599_ = _0056_ & ~io_in[13];
	assign _0064_ = _0055_ & ~io_in[13];
	assign _0075_ = _0064_ | _2599_;
	assign _0086_ = _0075_ | _2588_;
	assign _0097_ = _0054_ & ~io_in[13];
	assign _0108_ = _0053_ & ~io_in[13];
	assign _0119_ = _0108_ | _0097_;
	assign _0130_ = _0052_ & ~io_in[13];
	assign _0141_ = _0051_ & ~io_in[13];
	assign _0152_ = _0141_ | _0130_;
	assign _0162_ = _0152_ | _0119_;
	assign _0173_ = _0162_ | _0086_;
	assign _0184_ = _2555_ & ~_0173_;
	assign _0195_ = io_in[13] | ~_0023_;
	assign _0206_ = io_in[13] | ~_0020_;
	assign _0217_ = _0019_ & ~io_in[13];
	assign _0228_ = _0217_ & ~_0206_;
	assign _0238_ = io_in[13] | ~_0022_;
	assign _0249_ = io_in[13] | ~_0021_;
	assign _0260_ = _0249_ | _0238_;
	assign _0271_ = _0228_ & ~_0260_;
	assign _0282_ = _0271_ & ~_0195_;
	assign _0293_ = _0282_ & ~_0184_;
	assign _0304_ = _0044_ & ~io_in[13];
	assign _0315_ = _0043_ & ~io_in[13];
	assign _0325_ = _0315_ | _0304_;
	assign _0336_ = _0046_ & ~io_in[13];
	assign _0347_ = _0045_ & ~io_in[13];
	assign _0358_ = _0347_ | _0336_;
	assign _0369_ = _0358_ | _0325_;
	assign _0380_ = _0050_ & ~io_in[13];
	assign _0390_ = _0049_ & ~io_in[13];
	assign _0401_ = _0390_ | _0380_;
	assign _0412_ = _0048_ & ~io_in[13];
	assign _0423_ = _0047_ & ~io_in[13];
	assign _0434_ = _0423_ | _0412_;
	assign _0445_ = _0434_ | _0401_;
	assign _0456_ = _0445_ | _0369_;
	assign _0467_ = _0026_ & ~io_in[13];
	assign _0478_ = _0025_ & ~io_in[13];
	assign _0489_ = _0478_ | _0467_;
	assign _0500_ = _0489_ | _0456_;
	assign _0511_ = _0028_ & ~io_in[13];
	assign _0522_ = _0027_ & ~io_in[13];
	assign _0533_ = _0522_ & _0511_;
	assign _0544_ = _0030_ & ~io_in[13];
	assign _0555_ = _0029_ & ~io_in[13];
	assign _0566_ = ~(_0555_ & _0544_);
	assign _0577_ = _0566_ | ~_0533_;
	assign _0588_ = _0031_ & ~io_in[13];
	assign _0599_ = _0577_ | ~_0588_;
	assign _0610_ = _0500_ & ~_0599_;
	assign _0621_ = ~(_0610_ | _0293_);
	assign _0632_ = ~_0282_;
	assign _0641_ = _0184_ & ~_0632_;
	assign _0652_ = ~(_0599_ | _0500_);
	assign _0663_ = _0652_ | _0641_;
	assign _0674_ = _0062_ & ~io_in[13];
	assign _0684_ = _0061_ & ~io_in[13];
	assign _0695_ = ~(_0684_ | _0674_);
	assign _0705_ = _0663_ & ~_0695_;
	assign _0714_ = _0060_ & ~io_in[13];
	assign _0724_ = _0059_ & ~io_in[13];
	assign _0735_ = _0724_ | ~_0714_;
	assign _0746_ = _0695_ & ~_0735_;
	assign _0757_ = _0024_ & ~io_in[13];
	assign _0768_ = _0757_ ^ _0746_;
	assign _0779_ = _0032_ & ~io_in[13];
	assign _0790_ = _0779_ ^ _0768_;
	assign _0801_ = _0790_ | ~_0705_;
	assign _0812_ = ~_0141_;
	assign _0823_ = ~_0315_;
	assign _0834_ = _0315_ & _2533_;
	assign _0845_ = _0304_ & _2566_;
	assign _0856_ = _0347_ & _2577_;
	assign _0867_ = _0856_ ^ _0845_;
	assign _0878_ = _0315_ & _2544_;
	assign _0889_ = ~(_0878_ ^ _0867_);
	assign _0900_ = ~(_0336_ & _0064_);
	assign _0911_ = _0423_ & _0097_;
	assign _0922_ = _0900_ | ~_0911_;
	assign _0933_ = _0347_ & _2599_;
	assign _0944_ = ~(_0911_ ^ _0900_);
	assign _0955_ = _0944_ & _0933_;
	assign _0966_ = _0922_ & ~_0955_;
	assign _0977_ = _0966_ | _0889_;
	assign _0988_ = _0315_ & _2566_;
	assign _0999_ = _0304_ & _2577_;
	assign _1010_ = _0999_ & _0988_;
	assign _1021_ = _0966_ ^ _0889_;
	assign _1032_ = _1021_ & _1010_;
	assign _1043_ = _0977_ & ~_1032_;
	assign _1054_ = _0834_ & ~_1043_;
	assign _1065_ = _0390_ & _0141_;
	assign _1076_ = _0412_ & _0130_;
	assign _1087_ = _1076_ & _1065_;
	assign _1098_ = _0423_ & _0108_;
	assign _1109_ = _1076_ ^ _1065_;
	assign _1120_ = _1109_ & _1098_;
	assign _1131_ = ~(_1120_ | _1087_);
	assign _1142_ = _0390_ & _0130_;
	assign _1153_ = _0380_ & _0141_;
	assign _1164_ = _1153_ ^ _1142_;
	assign _1175_ = _0412_ & _0108_;
	assign _1186_ = _1175_ ^ _1164_;
	assign _1197_ = _1186_ & ~_1131_;
	assign _1208_ = _0944_ ^ _0933_;
	assign _1219_ = ~(_1186_ ^ _1131_);
	assign _1230_ = _1219_ & _1208_;
	assign _1241_ = ~(_1230_ | _1197_);
	assign _1252_ = _1153_ & _1142_;
	assign _1263_ = _1175_ & _1164_;
	assign _1274_ = ~(_1263_ | _1252_);
	assign _1285_ = _0380_ & _0130_;
	assign _1296_ = _0478_ & _0141_;
	assign _1307_ = _1296_ ^ _1285_;
	assign _1318_ = _0390_ & _0108_;
	assign _1329_ = _1318_ ^ _1307_;
	assign _1340_ = ~(_1329_ ^ _1274_);
	assign _1351_ = _0336_ & _2599_;
	assign _1362_ = _0412_ & _0097_;
	assign _1373_ = _0423_ & _0064_;
	assign _1383_ = _1373_ ^ _1362_;
	assign _1393_ = _1383_ ^ _1351_;
	assign _1404_ = _1393_ ^ _1340_;
	assign _1415_ = _1404_ & ~_1241_;
	assign _1426_ = _1021_ ^ _1010_;
	assign _1437_ = ~(_1404_ ^ _1241_);
	assign _1448_ = _1437_ & _1426_;
	assign _1459_ = ~(_1448_ | _1415_);
	assign _1469_ = _1329_ & ~_1274_;
	assign _1480_ = _1393_ & _1340_;
	assign _1491_ = ~(_1480_ | _1469_);
	assign _1501_ = _1296_ & _1285_;
	assign _1512_ = _1318_ & _1307_;
	assign _1523_ = ~(_1512_ | _1501_);
	assign _1533_ = _0478_ & _0130_;
	assign _1544_ = _0467_ & _0141_;
	assign _1555_ = _1544_ ^ _1533_;
	assign _1566_ = _0380_ & _0108_;
	assign _1577_ = _1566_ ^ _1555_;
	assign _1587_ = ~(_1577_ ^ _1523_);
	assign _1598_ = _0423_ & _2599_;
	assign _1609_ = ~(_0412_ & _0064_);
	assign _1620_ = _0390_ & _0097_;
	assign _1631_ = ~(_1620_ ^ _1609_);
	assign _1641_ = _1631_ ^ _1598_;
	assign _1652_ = _1641_ ^ _1587_;
	assign _1663_ = ~(_1652_ ^ _1491_);
	assign _1674_ = _0856_ & _0845_;
	assign _1685_ = _0878_ & _0867_;
	assign _1695_ = _1685_ | _1674_;
	assign _1706_ = _0347_ & _2566_;
	assign _1717_ = _0336_ & _2577_;
	assign _1728_ = _1717_ ^ _1706_;
	assign _1739_ = _0304_ & _2544_;
	assign _1750_ = ~(_1739_ ^ _1728_);
	assign _1760_ = _1373_ & _1362_;
	assign _1771_ = ~(_1383_ & _1351_);
	assign _1782_ = _1771_ & ~_1760_;
	assign _1793_ = _1782_ ^ _1750_;
	assign _1804_ = _1793_ ^ _1695_;
	assign _1814_ = _1804_ ^ _1663_;
	assign _1825_ = _1814_ & ~_1459_;
	assign _1836_ = ~(_1043_ ^ _0834_);
	assign _1847_ = ~(_1814_ ^ _1459_);
	assign _1858_ = _1847_ & _1836_;
	assign _1864_ = ~(_1858_ | _1825_);
	assign _1865_ = _0304_ & _2533_;
	assign _1866_ = _1782_ | _1750_;
	assign _1867_ = _1793_ & _1695_;
	assign _1868_ = _1866_ & ~_1867_;
	assign _1869_ = ~(_1868_ ^ _1865_);
	assign _1870_ = ~(_1869_ ^ _0823_);
	assign _1871_ = _1652_ & ~_1491_;
	assign _1872_ = _1804_ & _1663_;
	assign _1873_ = ~(_1872_ | _1871_);
	assign _1874_ = ~(_1717_ & _1706_);
	assign _1875_ = _1739_ & _1728_;
	assign _1876_ = _1874_ & ~_1875_;
	assign _1877_ = _0347_ & _2544_;
	assign _1878_ = _0336_ & _2566_;
	assign _1879_ = _0423_ & _2577_;
	assign _1880_ = _1879_ ^ _1878_;
	assign _1881_ = _1880_ ^ _1877_;
	assign _1882_ = _1609_ | ~_1620_;
	assign _1883_ = _1631_ & _1598_;
	assign _1884_ = _1882_ & ~_1883_;
	assign _1885_ = _1884_ ^ _1881_;
	assign _1886_ = _1885_ ^ _1876_;
	assign _1887_ = _1577_ & ~_1523_;
	assign _1888_ = _1641_ & _1587_;
	assign _1889_ = ~(_1888_ | _1887_);
	assign _1890_ = ~(_0390_ & _0064_);
	assign _1891_ = _0380_ & _0097_;
	assign _1892_ = ~(_1891_ ^ _1890_);
	assign _1893_ = _0412_ & _2599_;
	assign _1894_ = _1893_ ^ _1892_;
	assign _1895_ = _1544_ & _1533_;
	assign _1896_ = _1566_ & _1555_;
	assign _1897_ = ~(_1896_ | _1895_);
	assign _1898_ = _0478_ & _0108_;
	assign _1899_ = _0467_ & _0130_;
	assign _1900_ = _1899_ ^ _0141_;
	assign _1901_ = _1900_ ^ _1898_;
	assign _1902_ = ~(_1901_ ^ _1897_);
	assign _1903_ = _1902_ ^ _1894_;
	assign _1904_ = ~(_1903_ ^ _1889_);
	assign _1905_ = _1904_ ^ _1886_;
	assign _1906_ = ~(_1905_ ^ _1873_);
	assign _1907_ = _1906_ ^ _1870_;
	assign _1908_ = ~(_1907_ ^ _1864_);
	assign _1909_ = _1908_ ^ _1054_;
	assign _1910_ = _1847_ ^ _1836_;
	assign _1911_ = _0412_ & _0141_;
	assign _1912_ = _0423_ & _0130_;
	assign _1913_ = _1912_ & _1911_;
	assign _1914_ = _0336_ & _0108_;
	assign _1915_ = _1912_ ^ _1911_;
	assign _1916_ = _1915_ & _1914_;
	assign _1917_ = ~(_1916_ | _1913_);
	assign _1918_ = _1109_ ^ _1098_;
	assign _1919_ = _1918_ & ~_1917_;
	assign _1920_ = _0304_ & _2599_;
	assign _1921_ = _0347_ & _0064_;
	assign _1922_ = _0336_ & _0097_;
	assign _1923_ = _1922_ ^ _1921_;
	assign _1924_ = _1923_ ^ _1920_;
	assign _1925_ = ~(_1918_ ^ _1917_);
	assign _1926_ = _1925_ & _1924_;
	assign _1927_ = ~(_1926_ | _1919_);
	assign _1928_ = _1219_ ^ _1208_;
	assign _1929_ = _1927_ | ~_1928_;
	assign _1930_ = _0999_ ^ _0988_;
	assign _1931_ = ~(_1922_ & _1921_);
	assign _1932_ = _1923_ & _1920_;
	assign _1933_ = _1931_ & ~_1932_;
	assign _1934_ = ~(_1933_ ^ _1930_);
	assign _1935_ = ~(_1928_ ^ _1927_);
	assign _1936_ = _1935_ & _1934_;
	assign _1937_ = _1929_ & ~_1936_;
	assign _1938_ = _1437_ ^ _1426_;
	assign _1939_ = _1937_ | ~_1938_;
	assign _1940_ = _1930_ & ~_1933_;
	assign _1941_ = ~(_1938_ ^ _1937_);
	assign _1942_ = _1941_ & _1940_;
	assign _1943_ = _1939_ & ~_1942_;
	assign _1944_ = _1910_ & ~_1943_;
	assign _1945_ = _1944_ & _1909_;
	assign _1946_ = _1944_ ^ _1909_;
	assign _1947_ = _0423_ & _0141_;
	assign _1948_ = _0336_ & _0130_;
	assign _1949_ = _1948_ & _1947_;
	assign _1950_ = _0347_ & _0108_;
	assign _1951_ = _1948_ ^ _1947_;
	assign _1952_ = _1951_ & _1950_;
	assign _1953_ = ~(_1952_ | _1949_);
	assign _1954_ = _1915_ ^ _1914_;
	assign _1955_ = _1954_ & ~_1953_;
	assign _1956_ = _0315_ & _2599_;
	assign _1957_ = ~(_0304_ & _0064_);
	assign _1958_ = _0347_ & _0097_;
	assign _1959_ = ~(_1958_ ^ _1957_);
	assign _1960_ = _1959_ ^ _1956_;
	assign _1961_ = ~(_1954_ ^ _1953_);
	assign _1962_ = _1961_ & _1960_;
	assign _1963_ = ~(_1962_ | _1955_);
	assign _1964_ = _1925_ ^ _1924_;
	assign _1965_ = _1964_ & ~_1963_;
	assign _1966_ = _0315_ & _2577_;
	assign _1967_ = _1957_ | ~_1958_;
	assign _1968_ = _1959_ & _1956_;
	assign _1969_ = _1967_ & ~_1968_;
	assign _1970_ = ~(_1969_ ^ _1966_);
	assign _1971_ = ~(_1964_ ^ _1963_);
	assign _1972_ = _1971_ & _1970_;
	assign _1973_ = ~(_1972_ | _1965_);
	assign _1974_ = _1935_ ^ _1934_;
	assign _1975_ = _1974_ & ~_1973_;
	assign _1976_ = _1966_ & ~_1969_;
	assign _1977_ = ~(_1974_ ^ _1973_);
	assign _1978_ = _1977_ & _1976_;
	assign _1979_ = ~(_1978_ | _1975_);
	assign _1980_ = _1941_ ^ _1940_;
	assign _1981_ = _1980_ & ~_1979_;
	assign _1982_ = ~(_1943_ ^ _1910_);
	assign _1983_ = _1982_ & _1981_;
	assign _1984_ = ~(_1980_ ^ _1979_);
	assign _1985_ = _1971_ ^ _1970_;
	assign _1986_ = _0336_ & _0141_;
	assign _1987_ = _0347_ & _0130_;
	assign _1988_ = _1987_ & _1986_;
	assign _1989_ = _0304_ & _0108_;
	assign _1990_ = _1987_ ^ _1986_;
	assign _1991_ = _1990_ & _1989_;
	assign _1992_ = ~(_1991_ | _1988_);
	assign _1993_ = _1951_ ^ _1950_;
	assign _1994_ = _1993_ & ~_1992_;
	assign _1995_ = _0315_ & _0064_;
	assign _1996_ = _0304_ & _0097_;
	assign _1997_ = _1996_ ^ _1995_;
	assign _1998_ = ~(_1993_ ^ _1992_);
	assign _1999_ = _1998_ & _1997_;
	assign _2000_ = ~(_1999_ | _1994_);
	assign _2001_ = _1961_ ^ _1960_;
	assign _2002_ = _2000_ | ~_2001_;
	assign _2003_ = _1996_ & _1995_;
	assign _2004_ = ~(_2001_ ^ _2000_);
	assign _2005_ = _2004_ & _2003_;
	assign _2006_ = _2002_ & ~_2005_;
	assign _2007_ = _1985_ & ~_2006_;
	assign _2008_ = _1977_ ^ _1976_;
	assign _2009_ = _2008_ & _2007_;
	assign _2010_ = _2009_ & _1984_;
	assign _2011_ = _1982_ ^ _1981_;
	assign _2012_ = _2011_ & _2010_;
	assign _2013_ = ~(_2012_ | _1983_);
	assign _2014_ = _2009_ ^ _1984_;
	assign _2015_ = _2014_ & _2011_;
	assign _2016_ = _0315_ & _0130_;
	assign _2017_ = _0304_ & _0141_;
	assign _2018_ = _2017_ & _2016_;
	assign _2019_ = _0347_ & _0141_;
	assign _2020_ = _0304_ & _0130_;
	assign _2021_ = _2020_ ^ _2019_;
	assign _2022_ = _0315_ & _0108_;
	assign _2023_ = _2022_ ^ _2021_;
	assign _2024_ = _2023_ & _2018_;
	assign _2025_ = _2020_ & _2019_;
	assign _2026_ = _2022_ & _2021_;
	assign _2027_ = ~(_2026_ | _2025_);
	assign _2028_ = _1990_ ^ _1989_;
	assign _2029_ = ~(_2028_ ^ _2027_);
	assign _2030_ = _0315_ & _0097_;
	assign _2031_ = _2030_ ^ _2029_;
	assign _2032_ = _2031_ & _2024_;
	assign _2033_ = _2028_ & ~_2027_;
	assign _2034_ = _2030_ & _2029_;
	assign _2035_ = ~(_2034_ | _2033_);
	assign _2036_ = _1998_ ^ _1997_;
	assign _2037_ = ~(_2036_ ^ _2035_);
	assign _2038_ = _2037_ & _2032_;
	assign _2039_ = _2036_ & ~_2035_;
	assign _2040_ = _2004_ ^ _2003_;
	assign _2041_ = _2040_ ^ _2039_;
	assign _2042_ = _2041_ & _2038_;
	assign _2043_ = ~_2039_;
	assign _2044_ = _2040_ & ~_2043_;
	assign _2045_ = ~(_2006_ ^ _1985_);
	assign _2046_ = _2045_ ^ _2044_;
	assign _2047_ = _2046_ & _2042_;
	assign _2048_ = _2045_ & _2044_;
	assign _2049_ = _2008_ ^ _2007_;
	assign _2050_ = ~(_2049_ ^ _2048_);
	assign _2051_ = _2047_ & ~_2050_;
	assign _2052_ = _2049_ & _2048_;
	assign _2053_ = ~(_2052_ | _2051_);
	assign _2054_ = _2015_ & ~_2053_;
	assign _2055_ = _2013_ & ~_2054_;
	assign _2056_ = _1946_ & ~_2055_;
	assign _2057_ = ~(_2056_ | _1945_);
	assign _2058_ = _1864_ | ~_1907_;
	assign _2059_ = _1908_ & _1054_;
	assign _2060_ = _2058_ & ~_2059_;
	assign _2061_ = _1865_ & ~_1868_;
	assign _2062_ = _1869_ & ~_0823_;
	assign _2063_ = _2062_ | _2061_;
	assign _2064_ = _1905_ & ~_1873_;
	assign _2065_ = _1906_ & _1870_;
	assign _2066_ = ~(_2065_ | _2064_);
	assign _2067_ = ~_0304_;
	assign _2068_ = _0347_ & _2533_;
	assign _2069_ = _1885_ | _1876_;
	assign _2070_ = _1881_ & ~_1884_;
	assign _2071_ = _2069_ & ~_2070_;
	assign _2072_ = ~(_2071_ ^ _2068_);
	assign _2073_ = ~(_2072_ ^ _2067_);
	assign _2074_ = _1903_ & ~_1889_;
	assign _2075_ = _1904_ & _1886_;
	assign _2076_ = ~(_2075_ | _2074_);
	assign _2077_ = ~(_1879_ & _1878_);
	assign _2078_ = _1880_ & _1877_;
	assign _2079_ = _2077_ & ~_2078_;
	assign _2080_ = _0336_ & _2544_;
	assign _2081_ = _0423_ & _2566_;
	assign _2082_ = _0412_ & _2577_;
	assign _2083_ = _2082_ ^ _2081_;
	assign _2084_ = _2083_ ^ _2080_;
	assign _2085_ = _1890_ | ~_1891_;
	assign _2086_ = _1893_ & _1892_;
	assign _2087_ = _2085_ & ~_2086_;
	assign _2088_ = _2087_ ^ _2084_;
	assign _2089_ = _2088_ ^ _2079_;
	assign _2090_ = _1901_ & ~_1897_;
	assign _2091_ = _1902_ & _1894_;
	assign _2092_ = ~(_2091_ | _2090_);
	assign _2093_ = _0390_ & _2599_;
	assign _2094_ = ~(_0380_ & _0064_);
	assign _2095_ = _0478_ & _0097_;
	assign _2096_ = ~(_2095_ ^ _2094_);
	assign _2097_ = _2096_ ^ _2093_;
	assign _2098_ = _1899_ & ~_0812_;
	assign _2099_ = _1900_ & _1898_;
	assign _2100_ = ~(_2099_ | _2098_);
	assign _2101_ = _0467_ & _0108_;
	assign _2102_ = _2101_ ^ _0130_;
	assign _2103_ = ~(_2102_ ^ _2100_);
	assign _2104_ = _2103_ ^ _2097_;
	assign _2105_ = ~(_2104_ ^ _2092_);
	assign _2106_ = _2105_ ^ _2089_;
	assign _2107_ = ~(_2106_ ^ _2076_);
	assign _2108_ = _2107_ ^ _2073_;
	assign _2109_ = ~(_2108_ ^ _2066_);
	assign _2110_ = _2109_ ^ _2063_;
	assign _2111_ = ~(_2110_ ^ _2060_);
	assign _2112_ = ~(_2111_ ^ _2057_);
	assign _2113_ = ~_2533_;
	assign _2114_ = ~_2544_;
	assign _2115_ = ~_2566_;
	assign _2116_ = _0467_ & _2544_;
	assign _2117_ = _2116_ & ~_2115_;
	assign _2118_ = _2117_ & ~_2114_;
	assign _2119_ = _2118_ & ~_2113_;
	assign _2120_ = ~_0467_;
	assign _2121_ = _2118_ ^ _2533_;
	assign _2122_ = _2121_ & ~_2120_;
	assign _2123_ = ~(_2122_ | _2119_);
	assign _2124_ = ~_2123_;
	assign _2125_ = ~(_2121_ ^ _2120_);
	assign _2126_ = _2117_ ^ _2544_;
	assign _2127_ = ~_0478_;
	assign _2128_ = ~_2577_;
	assign _2129_ = _0467_ & _2566_;
	assign _2130_ = _2129_ & ~_2128_;
	assign _2131_ = _0478_ & _2544_;
	assign _2132_ = ~_2131_;
	assign _2133_ = _2129_ ^ _2577_;
	assign _2134_ = _2133_ & ~_2132_;
	assign _2135_ = ~(_2134_ | _2130_);
	assign _2136_ = _2116_ ^ _2566_;
	assign _2137_ = _2136_ & ~_2135_;
	assign _2138_ = _0467_ & _2533_;
	assign _2139_ = _2138_ ^ _2137_;
	assign _2140_ = ~(_2139_ ^ _2127_);
	assign _2141_ = _2140_ & _2126_;
	assign _2142_ = ~(_2141_ & _2125_);
	assign _2143_ = _2138_ & _2137_;
	assign _2144_ = _2139_ & ~_2127_;
	assign _2145_ = ~(_2144_ | _2143_);
	assign _2146_ = _2141_ ^ _2125_;
	assign _2147_ = _2146_ & ~_2145_;
	assign _2148_ = _2142_ & ~_2147_;
	assign _2149_ = _2148_ | _2124_;
	assign _2150_ = _2148_ ^ _2124_;
	assign _2151_ = _2140_ ^ _2126_;
	assign _2152_ = ~(_2136_ ^ _2135_);
	assign _2153_ = ~_0380_;
	assign _2154_ = _0478_ & _2533_;
	assign _2155_ = _0478_ & _2566_;
	assign _2156_ = _0467_ & _2577_;
	assign _2157_ = _2156_ & _2155_;
	assign _2158_ = _0380_ & _2544_;
	assign _2159_ = _2156_ ^ _2155_;
	assign _2160_ = _2159_ & _2158_;
	assign _2161_ = ~(_2160_ | _2157_);
	assign _2162_ = _2133_ ^ _2131_;
	assign _2163_ = _2162_ & ~_2161_;
	assign _2164_ = _2163_ ^ _2154_;
	assign _2165_ = ~(_2164_ ^ _2153_);
	assign _2166_ = _2165_ & _2152_;
	assign _2167_ = _2166_ & _2151_;
	assign _2168_ = _2163_ & _2154_;
	assign _2169_ = _2164_ & ~_2153_;
	assign _2170_ = ~(_2169_ | _2168_);
	assign _2171_ = _2166_ ^ _2151_;
	assign _2172_ = _2171_ & ~_2170_;
	assign _2173_ = ~(_2172_ | _2167_);
	assign _2174_ = ~(_2146_ ^ _2145_);
	assign _2175_ = _2173_ | ~_2174_;
	assign _2176_ = ~(_2174_ ^ _2173_);
	assign _2177_ = ~(_2162_ ^ _2161_);
	assign _2178_ = ~_2599_;
	assign _2179_ = _0380_ & _2566_;
	assign _2180_ = _0478_ & _2577_;
	assign _2181_ = ~(_2180_ & _2179_);
	assign _2182_ = _0390_ & _2544_;
	assign _2183_ = _2180_ ^ _2179_;
	assign _2184_ = _2183_ & _2182_;
	assign _2185_ = _2181_ & ~_2184_;
	assign _2186_ = _2159_ ^ _2158_;
	assign _2187_ = ~_0064_;
	assign _2188_ = _0467_ & _2599_;
	assign _2189_ = _2188_ & ~_2187_;
	assign _2190_ = ~_2189_;
	assign _2191_ = _2190_ ^ _2186_;
	assign _2192_ = _2191_ ^ _2185_;
	assign _2193_ = _2192_ & ~_2178_;
	assign _2194_ = _2193_ & _2177_;
	assign _2195_ = _2193_ ^ _2177_;
	assign _2196_ = ~_0390_;
	assign _2197_ = _0380_ & _2533_;
	assign _2198_ = _2191_ | _2185_;
	assign _2199_ = _2186_ & ~_2190_;
	assign _2200_ = _2198_ & ~_2199_;
	assign _2201_ = ~(_2200_ ^ _2197_);
	assign _2202_ = ~(_2201_ ^ _2196_);
	assign _2203_ = _2202_ & _2195_;
	assign _2204_ = ~(_2203_ | _2194_);
	assign _2205_ = _2165_ ^ _2152_;
	assign _2206_ = _2205_ & ~_2204_;
	assign _2207_ = _2197_ & ~_2200_;
	assign _2208_ = _2201_ & ~_2196_;
	assign _2209_ = _2208_ | _2207_;
	assign _2210_ = ~(_2205_ ^ _2204_);
	assign _2211_ = _2210_ & _2209_;
	assign _2212_ = ~(_2211_ | _2206_);
	assign _2213_ = ~(_2171_ ^ _2170_);
	assign _2214_ = _2212_ | ~_2213_;
	assign _2215_ = _2176_ & ~_2214_;
	assign _2216_ = _2175_ & ~_2215_;
	assign _2217_ = ~(_2213_ ^ _2212_);
	assign _2218_ = _2217_ & _2176_;
	assign _2219_ = _2192_ ^ _2599_;
	assign _2220_ = _2188_ ^ _0064_;
	assign _2221_ = _0380_ & _2577_;
	assign _2222_ = _0390_ & _2566_;
	assign _2223_ = _2222_ & _2221_;
	assign _2224_ = _0412_ & _2544_;
	assign _2225_ = _2222_ ^ _2221_;
	assign _2226_ = _2225_ & _2224_;
	assign _2227_ = _2226_ | _2223_;
	assign _2228_ = ~(_2183_ ^ _2182_);
	assign _2229_ = _0467_ & _0064_;
	assign _2230_ = ~(_2229_ & _0097_);
	assign _2231_ = _0478_ & _2599_;
	assign _2232_ = _2229_ ^ _0097_;
	assign _2233_ = _2232_ & _2231_;
	assign _2234_ = _2230_ & ~_2233_;
	assign _2235_ = _2234_ ^ _2228_;
	assign _2236_ = _2235_ ^ _2227_;
	assign _2237_ = _2236_ & _2220_;
	assign _2238_ = _2237_ & _2219_;
	assign _2239_ = _2237_ ^ _2219_;
	assign _2240_ = ~_0412_;
	assign _2241_ = _0390_ & _2533_;
	assign _2242_ = _2234_ | _2228_;
	assign _2243_ = _2235_ & _2227_;
	assign _2244_ = _2242_ & ~_2243_;
	assign _2245_ = ~(_2244_ ^ _2241_);
	assign _2246_ = ~(_2245_ ^ _2240_);
	assign _2247_ = _2246_ & _2239_;
	assign _2248_ = ~(_2247_ | _2238_);
	assign _2249_ = _2202_ ^ _2195_;
	assign _2250_ = _2248_ | ~_2249_;
	assign _2251_ = _2241_ & ~_2244_;
	assign _2252_ = _2245_ & ~_2240_;
	assign _2253_ = _2252_ | _2251_;
	assign _2254_ = ~(_2249_ ^ _2248_);
	assign _2255_ = _2254_ & _2253_;
	assign _2256_ = _2250_ & ~_2255_;
	assign _2257_ = _2210_ ^ _2209_;
	assign _2258_ = _2256_ | ~_2257_;
	assign _2259_ = ~_0108_;
	assign _2260_ = ~_0130_;
	assign _2261_ = _2101_ & ~_2260_;
	assign _2262_ = _2261_ & ~_2259_;
	assign _2263_ = _2261_ ^ _0108_;
	assign _2264_ = _0380_ & _2599_;
	assign _2265_ = ~(_0478_ & _0064_);
	assign _2266_ = _0467_ & _0097_;
	assign _2267_ = ~(_2266_ ^ _2265_);
	assign _2268_ = _2267_ ^ _2264_;
	assign _2269_ = _2268_ & _2263_;
	assign _2270_ = ~(_2269_ | _2262_);
	assign _2271_ = _2232_ ^ _2231_;
	assign _2272_ = _2271_ & ~_2270_;
	assign _2273_ = ~(_2271_ ^ _2270_);
	assign _2274_ = _0390_ & _2577_;
	assign _2275_ = _0412_ & _2566_;
	assign _2276_ = _2275_ & _2274_;
	assign _2277_ = _0423_ & _2544_;
	assign _2278_ = ~_2277_;
	assign _2279_ = _2275_ ^ _2274_;
	assign _2280_ = _2279_ & ~_2278_;
	assign _2281_ = _2280_ | _2276_;
	assign _2282_ = ~(_2225_ ^ _2224_);
	assign _2283_ = _2265_ | ~_2266_;
	assign _2284_ = _2267_ & _2264_;
	assign _2285_ = _2283_ & ~_2284_;
	assign _2286_ = _2285_ ^ _2282_;
	assign _2287_ = _2286_ ^ _2281_;
	assign _2288_ = _2287_ & _2273_;
	assign _2289_ = ~(_2288_ | _2272_);
	assign _2290_ = _2236_ ^ _2220_;
	assign _2291_ = _2290_ & ~_2289_;
	assign _2292_ = ~(_2290_ ^ _2289_);
	assign _2293_ = ~_0423_;
	assign _2294_ = _0412_ & _2533_;
	assign _2295_ = _2285_ | _2282_;
	assign _2296_ = _2286_ & _2281_;
	assign _2297_ = _2295_ & ~_2296_;
	assign _2298_ = ~(_2297_ ^ _2294_);
	assign _2299_ = ~(_2298_ ^ _2293_);
	assign _2300_ = _2299_ & _2292_;
	assign _2301_ = ~(_2300_ | _2291_);
	assign _2302_ = _2246_ ^ _2239_;
	assign _2303_ = _2302_ & ~_2301_;
	assign _2304_ = _2294_ & ~_2297_;
	assign _2305_ = _2298_ & ~_2293_;
	assign _2306_ = _2305_ | _2304_;
	assign _2307_ = ~(_2302_ ^ _2301_);
	assign _2308_ = _2307_ & _2306_;
	assign _2309_ = ~(_2308_ | _2303_);
	assign _2310_ = _2254_ ^ _2253_;
	assign _2311_ = _2310_ & ~_2309_;
	assign _2312_ = ~(_2257_ ^ _2256_);
	assign _2313_ = _2312_ & _2311_;
	assign _2314_ = _2258_ & ~_2313_;
	assign _2315_ = _2218_ & ~_2314_;
	assign _2316_ = _2216_ & ~_2315_;
	assign _2317_ = _2310_ ^ _2309_;
	assign _2318_ = _2312_ & ~_2317_;
	assign _2319_ = _2318_ & _2218_;
	assign _2320_ = _2102_ & ~_2100_;
	assign _2321_ = _2103_ & _2097_;
	assign _2322_ = ~(_2321_ | _2320_);
	assign _2323_ = _2268_ ^ _2263_;
	assign _2324_ = _2323_ & ~_2322_;
	assign _2325_ = _2082_ & _2081_;
	assign _2326_ = _2083_ & _2080_;
	assign _2327_ = _2326_ | _2325_;
	assign _2328_ = _2279_ ^ _2278_;
	assign _2329_ = _2094_ | ~_2095_;
	assign _2330_ = _2096_ & _2093_;
	assign _2331_ = _2329_ & ~_2330_;
	assign _2332_ = _2331_ ^ _2328_;
	assign _2333_ = _2332_ ^ _2327_;
	assign _2334_ = ~(_2323_ ^ _2322_);
	assign _2335_ = _2334_ & _2333_;
	assign _2336_ = ~(_2335_ | _2324_);
	assign _2337_ = _2287_ ^ _2273_;
	assign _2338_ = _2337_ & ~_2336_;
	assign _2339_ = ~_0336_;
	assign _2340_ = _0423_ & _2533_;
	assign _2341_ = _2331_ | _2328_;
	assign _2342_ = _2332_ & _2327_;
	assign _2343_ = _2341_ & ~_2342_;
	assign _2344_ = ~(_2343_ ^ _2340_);
	assign _2345_ = ~(_2344_ ^ _2339_);
	assign _2346_ = ~(_2337_ ^ _2336_);
	assign _2347_ = _2346_ & _2345_;
	assign _2348_ = ~(_2347_ | _2338_);
	assign _2349_ = _2299_ ^ _2292_;
	assign _2350_ = _2348_ | ~_2349_;
	assign _2351_ = _2340_ & ~_2343_;
	assign _2352_ = _2344_ & ~_2339_;
	assign _2353_ = _2352_ | _2351_;
	assign _2354_ = ~(_2349_ ^ _2348_);
	assign _2355_ = _2354_ & _2353_;
	assign _2356_ = _2350_ & ~_2355_;
	assign _2357_ = _2307_ ^ _2306_;
	assign _2358_ = _2356_ | ~_2357_;
	assign _2359_ = _2104_ & ~_2092_;
	assign _2360_ = _2105_ & _2089_;
	assign _2361_ = ~(_2360_ | _2359_);
	assign _2362_ = _2334_ ^ _2333_;
	assign _2363_ = _2362_ & ~_2361_;
	assign _2364_ = ~_0347_;
	assign _2365_ = _0336_ & _2533_;
	assign _2366_ = _2088_ | _2079_;
	assign _2367_ = _2084_ & ~_2087_;
	assign _2368_ = _2366_ & ~_2367_;
	assign _2369_ = ~(_2368_ ^ _2365_);
	assign _2370_ = ~(_2369_ ^ _2364_);
	assign _2371_ = ~(_2362_ ^ _2361_);
	assign _2372_ = _2371_ & _2370_;
	assign _2373_ = ~(_2372_ | _2363_);
	assign _2374_ = _2346_ ^ _2345_;
	assign _2375_ = _2374_ & ~_2373_;
	assign _2376_ = _2365_ & ~_2368_;
	assign _2377_ = _2369_ & ~_2364_;
	assign _2379_ = _2377_ | _2376_;
	assign _2380_ = ~(_2374_ ^ _2373_);
	assign _2381_ = _2380_ & _2379_;
	assign _2382_ = ~(_2381_ | _2375_);
	assign _2383_ = _2354_ ^ _2353_;
	assign _2384_ = _2383_ & ~_2382_;
	assign _2385_ = ~(_2357_ ^ _2356_);
	assign _2386_ = _2385_ & _2384_;
	assign _2387_ = _2358_ & ~_2386_;
	assign _2388_ = _2383_ ^ _2382_;
	assign _2390_ = _2385_ & ~_2388_;
	assign _2391_ = _2106_ & ~_2076_;
	assign _2392_ = _2107_ & _2073_;
	assign _2393_ = ~(_2392_ | _2391_);
	assign _2394_ = _2371_ ^ _2370_;
	assign _2395_ = _2393_ | ~_2394_;
	assign _2396_ = _2068_ & ~_2071_;
	assign _2397_ = _2072_ & ~_2067_;
	assign _2398_ = _2397_ | _2396_;
	assign _2399_ = ~(_2394_ ^ _2393_);
	assign _2400_ = _2399_ & _2398_;
	assign _2401_ = _2395_ & ~_2400_;
	assign _2402_ = _2380_ ^ _2379_;
	assign _2403_ = _2401_ | ~_2402_;
	assign _2404_ = _2108_ & ~_2066_;
	assign _2405_ = _2109_ & _2063_;
	assign _2406_ = ~(_2405_ | _2404_);
	assign _2407_ = _2399_ ^ _2398_;
	assign _2408_ = _2407_ & ~_2406_;
	assign _2409_ = ~(_2402_ ^ _2401_);
	assign _2411_ = _2409_ & _2408_;
	assign _2412_ = _2403_ & ~_2411_;
	assign _2413_ = _2390_ & ~_2412_;
	assign _2414_ = _2387_ & ~_2413_;
	assign _2415_ = _2407_ ^ _2406_;
	assign _2416_ = _2415_ | ~_2409_;
	assign _2417_ = _2390_ & ~_2416_;
	assign _2418_ = _2060_ | ~_2110_;
	assign _2419_ = _2111_ & _1945_;
	assign _2420_ = _2418_ & ~_2419_;
	assign _2421_ = ~(_2111_ & _1946_);
	assign _2422_ = ~(_2421_ | _2013_);
	assign _2423_ = _2420_ & ~_2422_;
	assign _2424_ = _2417_ & ~_2423_;
	assign _2425_ = _2414_ & ~_2424_;
	assign _2426_ = ~_2053_;
	assign _2427_ = _2421_ | ~_2015_;
	assign _2428_ = _2427_ | ~_2417_;
	assign _2429_ = _2426_ & ~_2428_;
	assign _2430_ = _2425_ & ~_2429_;
	assign _2432_ = _2319_ & ~_2430_;
	assign _2433_ = _2316_ & ~_2432_;
	assign _2434_ = _2150_ & ~_2433_;
	assign _2435_ = _2149_ & ~_2434_;
	assign _2436_ = _2435_ ^ _2123_;
	assign _2437_ = ~(_2055_ ^ _1946_);
	assign _2438_ = (_2436_ ? _2112_ : _2437_);
	assign _2439_ = ~_2438_;
	assign _2440_ = _2426_ & ~_2427_;
	assign _2441_ = _2423_ & ~_2440_;
	assign _2442_ = _2441_ ^ _2415_;
	assign _2443_ = (_2436_ ? _2442_ : _2112_);
	assign _2444_ = _2443_ & _2438_;
	assign _2445_ = ~(_2441_ | _2416_);
	assign _2446_ = _2412_ & ~_2445_;
	assign _2447_ = ~(_2446_ ^ _2388_);
	assign _2448_ = _2441_ | _2415_;
	assign _2449_ = _2448_ & ~_2408_;
	assign _2450_ = ~(_2449_ ^ _2409_);
	assign _2451_ = ~_2450_;
	assign _2452_ = (_2436_ ? _2447_ : _2451_);
	assign _2453_ = (_2436_ ? _2450_ : _2442_);
	assign _2454_ = _2452_ | ~_2453_;
	assign _2455_ = _2444_ & ~_2454_;
	assign _2456_ = _2430_ | _2317_;
	assign _2457_ = _2456_ & ~_2311_;
	assign _2458_ = ~(_2457_ ^ _2312_);
	assign _2459_ = _2430_ ^ _2317_;
	assign _2460_ = (_2436_ ? _2458_ : _2459_);
	assign _2461_ = ~_2458_;
	assign _2463_ = _2318_ & ~_2430_;
	assign _2464_ = _2314_ & ~_2463_;
	assign _2465_ = _2464_ ^ _2217_;
	assign _2466_ = (_2436_ ? _2465_ : _2461_);
	assign _2467_ = _2466_ | ~_2460_;
	assign _2468_ = _2446_ | _2388_;
	assign _2469_ = _2468_ & ~_2384_;
	assign _2470_ = _2469_ ^ _2385_;
	assign _2471_ = (_2436_ ? _2470_ : _2447_);
	assign _2472_ = ~_2459_;
	assign _2473_ = (_2436_ ? _2472_ : _2470_);
	assign _2474_ = _2473_ | _2471_;
	assign _2475_ = ~(_2474_ | _2467_);
	assign _2476_ = ~(_2475_ & _2455_);
	assign _2477_ = _2217_ & ~_2464_;
	assign _2478_ = _2214_ & ~_2477_;
	assign _2479_ = _2478_ ^ _2176_;
	assign _2480_ = (_2436_ ? _2479_ : _2465_);
	assign _2481_ = ~(_2433_ ^ _2150_);
	assign _2482_ = ~_2481_;
	assign _2483_ = (_2436_ ? _2482_ : _2479_);
	assign _2484_ = _2483_ | _2480_;
	assign _2485_ = _2484_ | _2476_;
	assign _2486_ = _2482_ & ~_2436_;
	assign _2487_ = ~(_2486_ | _2485_);
	assign _2488_ = ~(_2443_ ^ _2438_);
	assign _2489_ = (_2487_ ? _2488_ : _2438_);
	assign _2490_ = ~_2453_;
	assign _2491_ = ~_2014_;
	assign _2492_ = _2053_ | _2491_;
	assign _2493_ = _2492_ & ~_2010_;
	assign _2494_ = ~(_2493_ ^ _2011_);
	assign _2495_ = (_2436_ ? _2437_ : _2494_);
	assign _2496_ = ~_2495_;
	assign _2497_ = _2053_ ^ _2491_;
	assign _2498_ = (_2436_ ? _2494_ : _2497_);
	assign _2499_ = _0315_ & _0141_;
	assign _2500_ = _2017_ ^ _2016_;
	assign _2501_ = _2499_ & ~_2500_;
	assign _2502_ = _2023_ ^ _2018_;
	assign _2503_ = _2031_ ^ _2024_;
	assign _2504_ = _2503_ | _2502_;
	assign _2505_ = _2501_ & ~_2504_;
	assign _2506_ = _2046_ ^ _2042_;
	assign _2507_ = ~(_2050_ ^ _2047_);
	assign _2508_ = _2507_ | _2506_;
	assign _2509_ = _2037_ ^ _2032_;
	assign _2510_ = _2041_ ^ _2038_;
	assign _2511_ = _2510_ | _2509_;
	assign _2512_ = _2511_ | _2508_;
	assign _2513_ = _2505_ & ~_2512_;
	assign _2514_ = _2502_ | _2500_;
	assign _2515_ = _2509_ | _2503_;
	assign _2516_ = _2515_ | _2514_;
	assign _2517_ = _2510_ | _2506_;
	assign _2518_ = _2517_ | _2516_;
	assign _2519_ = _2518_ | _2507_;
	assign _2520_ = _2519_ | _2513_;
	assign _2521_ = _2520_ | _2498_;
	assign _2522_ = _2495_ & ~_2521_;
	assign _2524_ = (_2522_ ? _2490_ : _2496_);
	assign _2525_ = (_2524_ ? _2439_ : _2489_);
	assign _2526_ = _0195_ & ~_0271_;
	assign _2527_ = ~(_0555_ & _0511_);
	assign _2528_ = _0588_ | ~_0522_;
	assign _2529_ = _2528_ | _2527_;
	assign _2530_ = _0544_ & ~_2529_;
	assign _2531_ = ~(_2530_ | _0588_);
	assign _2532_ = ~(_2531_ | _2526_);
	assign _2534_ = _0022_ & ~io_in[13];
	assign _2535_ = _2531_ & _2526_;
	assign _2536_ = _2531_ & ~_2526_;
	assign _2537_ = _0228_ & ~_0249_;
	assign _2538_ = _2537_ ^ _0238_;
	assign _2539_ = _2526_ & ~_2531_;
	assign _2540_ = (_2539_ ? _2534_ : _2538_);
	assign _2541_ = (_2536_ ? _2538_ : _2540_);
	assign _2542_ = (_2535_ ? _2534_ : _2541_);
	assign _2543_ = ~_0544_;
	assign _2545_ = ~_0555_;
	assign _2546_ = _0533_ & ~_2545_;
	assign _2547_ = _2546_ ^ _2543_;
	assign _2548_ = (_2536_ ? _0544_ : _2547_);
	assign _2549_ = (_2535_ ? _0544_ : _2548_);
	assign _2550_ = ~(_2549_ | _2542_);
	assign _2551_ = _0021_ & ~io_in[13];
	assign _2552_ = _2551_ ^ _0228_;
	assign _2553_ = (_2539_ ? _0249_ : _2552_);
	assign _2554_ = (_2536_ ? _2552_ : _2553_);
	assign _2556_ = (_2535_ ? _0249_ : _2554_);
	assign _2557_ = _0555_ ^ _0533_;
	assign _2558_ = (_2536_ ? _2545_ : _2557_);
	assign _2559_ = (_2535_ ? _2545_ : _2558_);
	assign _2560_ = _2559_ & _2556_;
	assign _2561_ = _2542_ | ~_2549_;
	assign _2562_ = _2549_ | ~_2542_;
	assign _2563_ = _2562_ & _2561_;
	assign _2564_ = _2560_ & ~_2563_;
	assign _2565_ = ~(_2564_ | _2550_);
	assign _2567_ = _0020_ & ~io_in[13];
	assign _2568_ = _0217_ | _2567_;
	assign _2569_ = _0228_ | ~_2568_;
	assign _2570_ = (_2539_ ? _2567_ : _2569_);
	assign _2571_ = (_2536_ ? _2569_ : _2570_);
	assign _2572_ = (_2535_ ? _2567_ : _2571_);
	assign _2573_ = ~(_0522_ ^ _0511_);
	assign _2574_ = (_2536_ ? _0511_ : _2573_);
	assign _2575_ = (_2535_ ? _0511_ : _2574_);
	assign _2576_ = ~(_2575_ | _2572_);
	assign _2578_ = ~(_0522_ | _0217_);
	assign _2579_ = _2572_ | ~_2575_;
	assign _2580_ = _2575_ | ~_2572_;
	assign _2581_ = _2580_ & _2579_;
	assign _2582_ = _2578_ & ~_2581_;
	assign _2583_ = _2582_ | _2576_;
	assign _2584_ = _2556_ & ~_2559_;
	assign _2585_ = _2559_ & ~_2556_;
	assign _2586_ = ~(_2585_ | _2584_);
	assign _2587_ = _2563_ | _2586_;
	assign _2589_ = _2583_ & ~_2587_;
	assign _2590_ = _2565_ & ~_2589_;
	assign _2591_ = _0588_ ^ _0577_;
	assign _2592_ = (_2536_ ? _0588_ : _2591_);
	assign _2593_ = (_2535_ ? _0588_ : _2592_);
	assign _2594_ = _2593_ ^ _0282_;
	assign _2595_ = ~(_2594_ ^ _2590_);
	assign _2596_ = _2593_ & ~_0282_;
	assign _2597_ = _2593_ ^ _0632_;
	assign _2598_ = ~_2585_;
	assign _2600_ = _2563_ & ~_2598_;
	assign _2601_ = _2562_ & ~_2600_;
	assign _2602_ = _2563_ & _2586_;
	assign _2603_ = _0217_ | ~_0522_;
	assign _2604_ = ~_2603_;
	assign _2605_ = _2581_ & ~_2604_;
	assign _2606_ = _2580_ & ~_2605_;
	assign _2607_ = _2602_ & ~_2606_;
	assign _2608_ = _2601_ & ~_2607_;
	assign _2609_ = _2597_ & ~_2608_;
	assign _0065_ = _2609_ | _2596_;
	assign _0066_ = _0217_ & ~_0522_;
	assign _0067_ = _2603_ & ~_0066_;
	assign _0068_ = ~_0067_;
	assign _0069_ = _2581_ & ~_0068_;
	assign _0070_ = ~(_0069_ & _2602_);
	assign _0071_ = _2597_ & ~_0070_;
	assign _0072_ = _0065_ & ~_0071_;
	assign _0073_ = _2536_ & ~_0072_;
	assign _0074_ = _2563_ & _2584_;
	assign _0076_ = _2561_ & ~_0074_;
	assign _0077_ = _2581_ & ~_0066_;
	assign _0078_ = _2579_ & ~_0077_;
	assign _0079_ = _2602_ & ~_0078_;
	assign _0080_ = _0076_ & ~_0079_;
	assign _0081_ = ~(_0080_ ^ _2597_);
	assign _0082_ = _0072_ & _2536_;
	assign _0083_ = ~(_2608_ ^ _2597_);
	assign _0084_ = ~(_0071_ | _0065_);
	assign _0085_ = _0084_ | ~_2539_;
	assign _0087_ = _2539_ & ~_0065_;
	assign _0088_ = _0081_ & _0087_;
	assign _0089_ = (_0085_ ? _0088_ : _0083_);
	assign _0090_ = (_0082_ ? _0083_ : _0089_);
	assign _0091_ = (_0073_ ? _0081_ : _0090_);
	assign _0092_ = (_2535_ ? _2595_ : _0091_);
	assign _0093_ = (_2532_ ? _2595_ : _0092_);
	assign _0094_ = _2583_ & ~_2586_;
	assign _0095_ = ~(_2560_ | _0094_);
	assign _0096_ = _2563_ ^ _0095_;
	assign _0098_ = ~_2563_;
	assign _0099_ = _0078_ | ~_2586_;
	assign _0100_ = _0099_ & ~_2584_;
	assign _0101_ = _0100_ ^ _0098_;
	assign _0102_ = _2586_ & ~_2606_;
	assign _0103_ = _2598_ & ~_0102_;
	assign _0104_ = _0103_ ^ _0098_;
	assign _0105_ = _0101_ & _0087_;
	assign _0106_ = (_0085_ ? _0105_ : _0104_);
	assign _0107_ = (_0082_ ? _0104_ : _0106_);
	assign _0109_ = (_0073_ ? _0101_ : _0107_);
	assign _0110_ = (_2535_ ? _0096_ : _0109_);
	assign _0111_ = (_2532_ ? _0096_ : _0110_);
	assign _0112_ = _0085_ & _0087_;
	assign _0113_ = (_2536_ ? _0072_ : _0112_);
	assign _0114_ = ~(_0113_ | _2535_);
	assign _0115_ = ~(_0114_ | _2532_);
	assign _0116_ = ~_0115_;
	assign _0117_ = _0111_ & ~_0116_;
	assign _0118_ = ~(_2586_ ^ _2583_);
	assign _0120_ = ~(_0078_ ^ _2586_);
	assign _0121_ = ~(_2606_ ^ _2586_);
	assign _0122_ = _0120_ & _0087_;
	assign _0123_ = (_0085_ ? _0122_ : _0121_);
	assign _0124_ = (_0082_ ? _0121_ : _0123_);
	assign _0125_ = (_0073_ ? _0120_ : _0124_);
	assign _0126_ = (_2535_ ? _0118_ : _0125_);
	assign _0127_ = (_2532_ ? _0118_ : _0126_);
	assign _0128_ = _0127_ & ~_0116_;
	assign _0129_ = _0115_ ^ _0111_;
	assign _0131_ = _0129_ & _0128_;
	assign _0132_ = ~(_0131_ | _0117_);
	assign _0133_ = _0127_ ^ _0115_;
	assign _0134_ = _0133_ & _0129_;
	assign _0135_ = ~(_2581_ ^ _2578_);
	assign _0136_ = ~(_0066_ ^ _2581_);
	assign _0137_ = ~(_2604_ ^ _2581_);
	assign _0138_ = _0136_ & _0087_;
	assign _0139_ = (_0085_ ? _0138_ : _0137_);
	assign _0140_ = (_0082_ ? _0137_ : _0139_);
	assign _0142_ = (_0073_ ? _0136_ : _0140_);
	assign _0143_ = (_2535_ ? _0135_ : _0142_);
	assign _0144_ = (_2532_ ? _0135_ : _0143_);
	assign _0145_ = ~(_0144_ & _0115_);
	assign _0146_ = _0144_ ^ _0115_;
	assign _0147_ = _0522_ ^ _0217_;
	assign _0148_ = _0147_ & _0146_;
	assign _0149_ = _0145_ & ~_0148_;
	assign _0150_ = _0134_ & ~_0149_;
	assign _0151_ = _0132_ & ~_0150_;
	assign _0153_ = _0093_ ^ _0115_;
	assign _0154_ = ~(_0153_ ^ _0151_);
	assign _0155_ = (_2436_ ? _0154_ : _0093_);
	assign _0156_ = ~_0155_;
	assign _0157_ = ~_0133_;
	assign _0158_ = _0149_ | _0157_;
	assign _0159_ = _0158_ & ~_0128_;
	assign _0160_ = ~(_0159_ ^ _0129_);
	assign _0161_ = _0149_ ^ _0157_;
	assign _0163_ = ~(_0161_ | _0160_);
	assign _0164_ = _0163_ & _0148_;
	assign _0165_ = _0164_ & ~_0154_;
	assign _0166_ = _0115_ & ~_0165_;
	assign _0167_ = (_2436_ ? _0166_ : _0115_);
	assign _0168_ = (_2436_ ? _0160_ : _0111_);
	assign _0169_ = (_2436_ ? _0161_ : _0127_);
	assign _0170_ = _0169_ | _0168_;
	assign _0171_ = _0147_ ^ _0146_;
	assign _0172_ = (_2436_ ? _0171_ : _0144_);
	assign _0174_ = _0147_ ^ _2436_;
	assign _0175_ = ~(_0174_ | _0172_);
	assign _0176_ = _0175_ & ~_0170_;
	assign _0177_ = _0176_ ^ _0156_;
	assign _0178_ = _0167_ & ~_0177_;
	assign _0179_ = ~_0178_;
	assign _0180_ = (_2487_ ? _0179_ : _0156_);
	assign _0181_ = (_2524_ ? _0156_ : _0180_);
	assign _0182_ = _0174_ ^ _0172_;
	assign _0183_ = _0167_ & ~_0182_;
	assign _0185_ = _0167_ & ~_0174_;
	assign _0186_ = _0185_ | _0183_;
	assign _0187_ = ~_0169_;
	assign _0188_ = ~(_0175_ & _0187_);
	assign _0189_ = _0188_ ^ _0168_;
	assign _0190_ = _0167_ & ~_0189_;
	assign _0191_ = _0175_ ^ _0187_;
	assign _0192_ = _0167_ & ~_0191_;
	assign _0193_ = _0192_ | _0190_;
	assign _0194_ = _0193_ | _0186_;
	assign _0196_ = _0179_ & ~_0194_;
	assign _0197_ = _0167_ & ~_0196_;
	assign _0198_ = (_2487_ ? _0197_ : _0167_);
	assign _0199_ = (_2524_ ? _0167_ : _0198_);
	assign _0200_ = ~(_0199_ | _0181_);
	assign _0201_ = _0200_ | _2525_;
	assign _0202_ = (_2487_ ? _0192_ : _0169_);
	assign _0203_ = (_2524_ ? _0169_ : _0202_);
	assign _0204_ = (_2487_ ? _0190_ : _0168_);
	assign _0205_ = (_2524_ ? _0168_ : _0204_);
	assign _0207_ = _0205_ & _0203_;
	assign _0208_ = (_2487_ ? _0183_ : _0172_);
	assign _0209_ = (_2524_ ? _0172_ : _0208_);
	assign _0210_ = (_2487_ ? _0185_ : _0174_);
	assign _0211_ = (_2524_ ? _0174_ : _0210_);
	assign _0212_ = _0209_ & ~_0211_;
	assign _0213_ = _0212_ & _0207_;
	assign _0214_ = ~(_0213_ & _0181_);
	assign _0215_ = ~(_0211_ & _0209_);
	assign _0216_ = _0207_ & ~_0215_;
	assign _0218_ = _0181_ & ~_0216_;
	assign _0219_ = _0214_ & ~_0218_;
	assign _0220_ = _0199_ & ~_0219_;
	assign _0221_ = (_0220_ ? _2525_ : _0201_);
	assign _0222_ = _0199_ & ~_0218_;
	assign _0223_ = _0222_ | _0221_;
	assign _0224_ = ~(_0724_ | _0714_);
	assign _0225_ = _0588_ ^ _0195_;
	assign _0226_ = _0544_ ^ _0238_;
	assign _0227_ = _0555_ ^ _2551_;
	assign _0229_ = _0226_ & ~_0227_;
	assign _0230_ = _0511_ ^ _2567_;
	assign _0231_ = ~(_0230_ | _0147_);
	assign _0232_ = ~(_0231_ & _0229_);
	assign _0233_ = _0225_ & ~_0232_;
	assign _0234_ = _0467_ ^ _2533_;
	assign _0235_ = ~_0234_;
	assign _0236_ = _2533_ & ~_0467_;
	assign _0237_ = _2544_ & ~_0478_;
	assign _0239_ = _0237_ & ~_0234_;
	assign _0240_ = _0239_ | _0236_;
	assign _0241_ = _0478_ ^ _2544_;
	assign _0242_ = ~(_0241_ | _0234_);
	assign _0243_ = _0380_ | ~_2566_;
	assign _0244_ = _0380_ ^ _2566_;
	assign _0245_ = _2577_ & ~_0390_;
	assign _0246_ = _0245_ & ~_0244_;
	assign _0247_ = _0243_ & ~_0246_;
	assign _0248_ = _0390_ ^ _2577_;
	assign _0250_ = ~(_0248_ | _0244_);
	assign _0251_ = _0412_ | ~_2599_;
	assign _0252_ = _0423_ | ~_0064_;
	assign _0253_ = ~(_0412_ ^ _2599_);
	assign _0254_ = _0253_ & ~_0252_;
	assign _0255_ = _0251_ & ~_0254_;
	assign _0256_ = _0250_ & ~_0255_;
	assign _0257_ = _0247_ & ~_0256_;
	assign _0258_ = _0423_ ^ _0064_;
	assign _0259_ = _0258_ | ~_0253_;
	assign _0261_ = _0250_ & ~_0259_;
	assign _0262_ = _0336_ | ~_0097_;
	assign _0263_ = ~(_0336_ ^ _0097_);
	assign _0264_ = _0347_ | ~_0108_;
	assign _0265_ = _0263_ & ~_0264_;
	assign _0266_ = _0262_ & ~_0265_;
	assign _0267_ = _0347_ ^ _0108_;
	assign _0268_ = _0263_ & ~_0267_;
	assign _0269_ = _0304_ | ~_0130_;
	assign _0270_ = ~(_0304_ ^ _0130_);
	assign _0272_ = _0315_ & ~_0141_;
	assign _0273_ = _0270_ & ~_0272_;
	assign _0274_ = _0269_ & ~_0273_;
	assign _0275_ = _0268_ & ~_0274_;
	assign _0276_ = _0266_ & ~_0275_;
	assign _0277_ = _0261_ & ~_0276_;
	assign _0278_ = _0257_ & ~_0277_;
	assign _0279_ = _0242_ & ~_0278_;
	assign _0280_ = _0279_ | _0240_;
	assign _0281_ = (_0280_ ? _2127_ : _2114_);
	assign _0283_ = (_0280_ ? _2114_ : _2127_);
	assign _0284_ = _0281_ & ~_0283_;
	assign _0285_ = ~(_0467_ ^ _2533_);
	assign _0286_ = ~_0285_;
	assign _0287_ = _0284_ & ~_0286_;
	assign _0288_ = _0235_ & ~_0287_;
	assign _0289_ = (_0280_ ? _2153_ : _2115_);
	assign _0290_ = (_0280_ ? _2115_ : _2153_);
	assign _0291_ = _0290_ | ~_0289_;
	assign _0292_ = (_0280_ ? _2196_ : _2128_);
	assign _0294_ = (_0280_ ? _2128_ : _2196_);
	assign _0295_ = _0292_ & ~_0294_;
	assign _0296_ = ~(_0380_ ^ _2566_);
	assign _0297_ = ~_0296_;
	assign _0298_ = _0295_ & ~_0297_;
	assign _0299_ = _0291_ & ~_0298_;
	assign _0300_ = (_0280_ ? _0423_ : _0064_);
	assign _0301_ = (_0280_ ? _2187_ : _2293_);
	assign _0302_ = _0301_ | _0300_;
	assign _0303_ = _0253_ & ~_0302_;
	assign _0305_ = (_0280_ ? _2240_ : _2178_);
	assign _0306_ = (_0280_ ? _2178_ : _2240_);
	assign _0307_ = _0305_ & ~_0306_;
	assign _0308_ = ~(_0307_ | _0303_);
	assign _0309_ = _0248_ | ~_0296_;
	assign _0310_ = ~(_0309_ | _0308_);
	assign _0311_ = _0299_ & ~_0310_;
	assign _0312_ = ~_0097_;
	assign _0313_ = (_0280_ ? _2339_ : _0312_);
	assign _0314_ = (_0280_ ? _0312_ : _2339_);
	assign _0316_ = _0314_ | ~_0313_;
	assign _0317_ = (_0280_ ? _2364_ : _2259_);
	assign _0318_ = (_0280_ ? _2259_ : _2364_);
	assign _0319_ = _0317_ & ~_0318_;
	assign _0320_ = ~_0263_;
	assign _0321_ = _0319_ & ~_0320_;
	assign _0322_ = _0316_ & ~_0321_;
	assign _0323_ = (_0280_ ? _0812_ : _0823_);
	assign _0324_ = (_0280_ ? _0823_ : _0812_);
	assign _0326_ = _0323_ & ~_0324_;
	assign _0327_ = _0326_ | ~_0270_;
	assign _0328_ = (_0280_ ? _2067_ : _2260_);
	assign _0329_ = (_0280_ ? _2260_ : _2067_);
	assign _0330_ = _0328_ & ~_0329_;
	assign _0331_ = _0327_ & ~_0330_;
	assign _0332_ = _0267_ | ~_0263_;
	assign _0333_ = ~(_0332_ | _0331_);
	assign _0334_ = _0322_ & ~_0333_;
	assign _0335_ = _0309_ | _0259_;
	assign _0337_ = ~(_0335_ | _0334_);
	assign _0338_ = _0311_ & ~_0337_;
	assign _0339_ = _0241_ | ~_0285_;
	assign _0340_ = ~(_0339_ | _0338_);
	assign _0341_ = _0288_ & ~_0340_;
	assign _0342_ = _0341_ | ~_0790_;
	assign _0343_ = ~(_0588_ | _0195_);
	assign _0344_ = _0544_ ^ _2534_;
	assign _0345_ = _0555_ | _0249_;
	assign _0346_ = _0345_ | _0344_;
	assign _0348_ = _2534_ & ~_0544_;
	assign _0349_ = _0346_ & ~_0348_;
	assign _0350_ = _0511_ | _0206_;
	assign _0351_ = _2603_ & ~_0230_;
	assign _0352_ = _0350_ & ~_0351_;
	assign _0353_ = _0229_ & ~_0352_;
	assign _0354_ = _0349_ & ~_0353_;
	assign _0355_ = _0225_ & ~_0354_;
	assign _0356_ = _0355_ | _0343_;
	assign _0357_ = (_0356_ ? _2534_ : _0544_);
	assign _0359_ = (_0356_ ? _0544_ : _2534_);
	assign _0360_ = _0357_ & ~_0359_;
	assign _0361_ = (_0356_ ? _0249_ : _2545_);
	assign _0362_ = (_0356_ ? _0555_ : _2551_);
	assign _0363_ = _0362_ | _0361_;
	assign _0364_ = _0226_ & ~_0363_;
	assign _0365_ = _0364_ | _0360_;
	assign _0366_ = (_0356_ ? _0217_ : _0522_);
	assign _0367_ = ~_0217_;
	assign _0368_ = ~_0522_;
	assign _0370_ = (_0356_ ? _0368_ : _0367_);
	assign _0371_ = ~(_0370_ | _0366_);
	assign _0372_ = _0511_ ^ _0206_;
	assign _0373_ = _0371_ | ~_0372_;
	assign _0374_ = (_0356_ ? _2567_ : _0511_);
	assign _0375_ = (_0356_ ? _0511_ : _2567_);
	assign _0376_ = _0374_ & ~_0375_;
	assign _0377_ = _0373_ & ~_0376_;
	assign _0378_ = _0229_ & ~_0377_;
	assign _0379_ = _0378_ | _0365_;
	assign _0381_ = _0225_ ^ _0379_;
	assign _0382_ = ~(_0377_ | _0227_);
	assign _0383_ = _0363_ & ~_0382_;
	assign _0384_ = _0383_ ^ _0344_;
	assign _0385_ = _0377_ ^ _0227_;
	assign _0386_ = _0372_ ^ _0371_;
	assign _0387_ = (_0356_ ? _2127_ : _2114_);
	assign _0388_ = (_0356_ ? _0467_ : _2533_);
	assign _0389_ = ~_0388_;
	assign _0391_ = (_0067_ ? _0387_ : _0389_);
	assign _0392_ = (_0386_ ? _0391_ : _0068_);
	assign _0393_ = _0392_ | _0385_;
	assign _0394_ = _0393_ | _0384_;
	assign _0395_ = ~(_0394_ | _0381_);
	assign _0396_ = (_0356_ ? _2114_ : _2127_);
	assign _0397_ = ~(_0396_ | _0395_);
	assign _0398_ = _0067_ & ~_0388_;
	assign _0399_ = (_0356_ ? _2153_ : _2115_);
	assign _0400_ = (_0067_ ? _0399_ : _0387_);
	assign _0402_ = (_0386_ ? _0400_ : _0398_);
	assign _0403_ = _0402_ | _0385_;
	assign _0404_ = _0403_ | _0384_;
	assign _0405_ = ~(_0404_ | _0381_);
	assign _0406_ = (_0356_ ? _2115_ : _2153_);
	assign _0407_ = ~(_0406_ | _0405_);
	assign _0408_ = _0396_ ^ _0395_;
	assign _0409_ = _0408_ & _0407_;
	assign _0410_ = _0409_ | _0397_;
	assign _0411_ = (_0356_ ? _0390_ : _2577_);
	assign _0413_ = ~_0411_;
	assign _0414_ = (_0067_ ? _0413_ : _0399_);
	assign _0415_ = (_0386_ ? _0414_ : _0391_);
	assign _0416_ = ~(_0386_ & _0067_);
	assign _0417_ = (_0385_ ? _0416_ : _0415_);
	assign _0418_ = _0417_ | _0384_;
	assign _0419_ = ~(_0418_ | _0381_);
	assign _0420_ = (_0356_ ? _2128_ : _2196_);
	assign _0421_ = ~(_0420_ | _0419_);
	assign _0422_ = (_0356_ ? _0412_ : _2599_);
	assign _0424_ = ~_0422_;
	assign _0425_ = (_0067_ ? _0424_ : _0413_);
	assign _0426_ = (_0386_ ? _0425_ : _0400_);
	assign _0427_ = _0398_ | ~_0386_;
	assign _0428_ = (_0385_ ? _0427_ : _0426_);
	assign _0429_ = _0428_ | _0384_;
	assign _0430_ = ~(_0429_ | _0381_);
	assign _0431_ = (_0356_ ? _2178_ : _2240_);
	assign _0432_ = ~(_0431_ | _0430_);
	assign _0433_ = _0420_ ^ _0419_;
	assign _0435_ = _0433_ & _0432_;
	assign _0436_ = ~(_0435_ | _0421_);
	assign _0437_ = _0406_ ^ _0405_;
	assign _0438_ = ~(_0437_ & _0408_);
	assign _0439_ = ~(_0438_ | _0436_);
	assign _0440_ = _0439_ | _0410_;
	assign _0441_ = (_0356_ ? _0423_ : _0064_);
	assign _0442_ = ~_0441_;
	assign _0443_ = (_0067_ ? _0442_ : _0424_);
	assign _0444_ = (_0386_ ? _0443_ : _0414_);
	assign _0446_ = (_0385_ ? _0392_ : _0444_);
	assign _0447_ = _0446_ | _0384_;
	assign _0448_ = _0447_ | _0381_;
	assign _0449_ = (_0356_ ? _0064_ : _0423_);
	assign _0450_ = _0449_ & _0448_;
	assign _0451_ = (_0356_ ? _0336_ : _0097_);
	assign _0452_ = ~_0451_;
	assign _0453_ = (_0067_ ? _0452_ : _0442_);
	assign _0454_ = (_0386_ ? _0453_ : _0425_);
	assign _0455_ = (_0385_ ? _0402_ : _0454_);
	assign _0457_ = _0455_ | _0384_;
	assign _0458_ = ~(_0457_ | _0381_);
	assign _0459_ = (_0356_ ? _0312_ : _2339_);
	assign _0460_ = ~(_0459_ | _0458_);
	assign _0461_ = ~(_0449_ ^ _0448_);
	assign _0462_ = _0460_ & ~_0461_;
	assign _0463_ = _0462_ | _0450_;
	assign _0464_ = _0416_ | _0385_;
	assign _0465_ = (_0356_ ? _0347_ : _0108_);
	assign _0466_ = ~_0465_;
	assign _0468_ = (_0067_ ? _0466_ : _0452_);
	assign _0469_ = (_0386_ ? _0468_ : _0443_);
	assign _0470_ = (_0385_ ? _0415_ : _0469_);
	assign _0471_ = (_0384_ ? _0464_ : _0470_);
	assign _0472_ = _0471_ | _0381_;
	assign _0473_ = (_0356_ ? _0108_ : _0347_);
	assign _0474_ = _0473_ & _0472_;
	assign _0475_ = _0427_ | _0385_;
	assign _0476_ = (_0356_ ? _0304_ : _0130_);
	assign _0477_ = ~_0476_;
	assign _0479_ = (_0067_ ? _0477_ : _0466_);
	assign _0480_ = (_0386_ ? _0479_ : _0453_);
	assign _0481_ = (_0385_ ? _0426_ : _0480_);
	assign _0482_ = (_0384_ ? _0475_ : _0481_);
	assign _0483_ = ~(_0482_ | _0381_);
	assign _0484_ = (_0356_ ? _2260_ : _2067_);
	assign _0485_ = ~(_0484_ | _0483_);
	assign _0486_ = ~(_0473_ ^ _0472_);
	assign _0487_ = _0485_ & ~_0486_;
	assign _0488_ = ~(_0487_ | _0474_);
	assign _0490_ = _0459_ ^ _0458_;
	assign _0491_ = _0461_ | ~_0490_;
	assign _0492_ = ~(_0491_ | _0488_);
	assign _0493_ = _0492_ | _0463_;
	assign _0494_ = (_0356_ ? _0315_ : _0141_);
	assign _0495_ = ~_0494_;
	assign _0496_ = (_0067_ ? _0495_ : _0477_);
	assign _0497_ = (_0386_ ? _0496_ : _0468_);
	assign _0498_ = (_0385_ ? _0444_ : _0497_);
	assign _0499_ = (_0384_ ? _0393_ : _0498_);
	assign _0501_ = _0499_ | _0381_;
	assign _0502_ = (_0356_ ? _0812_ : _0823_);
	assign _0503_ = _0501_ & ~_0502_;
	assign _0504_ = _0496_ | _0386_;
	assign _0505_ = (_0385_ ? _0469_ : _0504_);
	assign _0506_ = (_0384_ ? _0417_ : _0505_);
	assign _0507_ = _0506_ | _0381_;
	assign _0508_ = _0385_ | _0384_;
	assign _0509_ = ~(_0386_ & _0068_);
	assign _0510_ = _0509_ | _0508_;
	assign _0512_ = ~(_0510_ | _0381_);
	assign _0513_ = _0379_ | ~_0225_;
	assign _0514_ = _0381_ | ~_0513_;
	assign _0515_ = _0386_ | _0068_;
	assign _0516_ = _0515_ | _0508_;
	assign _0517_ = ~(_0516_ | _0514_);
	assign _0518_ = _0386_ | _0067_;
	assign _0519_ = ~_0385_;
	assign _0520_ = ~(_0519_ & _0384_);
	assign _0521_ = _0518_ & ~_0520_;
	assign _0523_ = _0384_ & ~_0521_;
	assign _0524_ = _0523_ | _0514_;
	assign _0525_ = _0513_ & ~_0524_;
	assign _0526_ = _0520_ | _0515_;
	assign _0527_ = _0526_ | _0514_;
	assign _0528_ = _0513_ & ~_0527_;
	assign _0529_ = _0399_ & ~_0411_;
	assign _0530_ = _0441_ | _0422_;
	assign _0531_ = _0529_ & ~_0530_;
	assign _0532_ = _0494_ | _0476_;
	assign _0534_ = _0465_ | _0451_;
	assign _0535_ = _0534_ | _0532_;
	assign _0536_ = _0531_ & ~_0535_;
	assign _0537_ = _0528_ & ~_0536_;
	assign _0538_ = _0525_ & ~_0537_;
	assign _0539_ = _0520_ | _0509_;
	assign _0540_ = ~(_0539_ | _0514_);
	assign _0541_ = _0535_ | _0530_;
	assign _0542_ = _0413_ & ~_0541_;
	assign _0543_ = _0540_ & ~_0542_;
	assign _0545_ = _0538_ & ~_0543_;
	assign _0546_ = _0520_ | _0416_;
	assign _0547_ = _0546_ | _0514_;
	assign _0548_ = _0541_ & ~_0547_;
	assign _0549_ = _0545_ & ~_0548_;
	assign _0550_ = _0519_ | _0384_;
	assign _0551_ = _0550_ | _0518_;
	assign _0552_ = ~(_0551_ | _0514_);
	assign _0553_ = _0442_ & ~_0535_;
	assign _0554_ = _0552_ & ~_0553_;
	assign _0556_ = _0549_ & ~_0554_;
	assign _0557_ = _0550_ | _0515_;
	assign _0558_ = _0557_ | _0514_;
	assign _0559_ = _0535_ & ~_0558_;
	assign _0560_ = _0556_ & ~_0559_;
	assign _0561_ = _0550_ | _0509_;
	assign _0562_ = ~(_0561_ | _0514_);
	assign _0563_ = _0466_ & ~_0532_;
	assign _0564_ = _0562_ & ~_0563_;
	assign _0565_ = _0560_ & ~_0564_;
	assign _0567_ = _0550_ | _0416_;
	assign _0568_ = _0567_ | _0514_;
	assign _0569_ = _0532_ & ~_0568_;
	assign _0570_ = _0565_ & ~_0569_;
	assign _0571_ = _0508_ | _0518_;
	assign _0572_ = _0571_ | _0514_;
	assign _0573_ = ~(_0572_ | _0495_);
	assign _0574_ = _0570_ & ~_0573_;
	assign _0575_ = _0574_ | _0517_;
	assign _0576_ = ~(_0575_ | _0512_);
	assign _0578_ = _0507_ & ~_0576_;
	assign _0579_ = ~(_0494_ & _0068_);
	assign _0580_ = (_0386_ ? _0579_ : _0479_);
	assign _0581_ = (_0385_ ? _0454_ : _0580_);
	assign _0582_ = (_0384_ ? _0403_ : _0581_);
	assign _0583_ = ~(_0582_ | _0381_);
	assign _0584_ = _0502_ ^ _0501_;
	assign _0585_ = _0584_ | _0583_;
	assign _0586_ = _0578_ & ~_0585_;
	assign _0587_ = _0586_ | _0503_;
	assign _0589_ = _0484_ ^ _0483_;
	assign _0590_ = _0486_ | ~_0589_;
	assign _0591_ = _0590_ | _0491_;
	assign _0592_ = _0587_ & ~_0591_;
	assign _0593_ = _0592_ | _0493_;
	assign _0594_ = _0431_ ^ _0430_;
	assign _0595_ = ~(_0594_ & _0433_);
	assign _0596_ = _0595_ | _0438_;
	assign _0597_ = _0593_ & ~_0596_;
	assign _0598_ = _0597_ | _0440_;
	assign _0600_ = _0475_ | _0384_;
	assign _0601_ = ~(_0600_ | _0381_);
	assign _0602_ = (_0356_ ? _2533_ : _0467_);
	assign _0603_ = ~(_0602_ ^ _0601_);
	assign _0604_ = _0464_ | _0384_;
	assign _0605_ = _0604_ | _0381_;
	assign _0606_ = _0605_ | ~_0603_;
	assign _0607_ = _0606_ | ~_0598_;
	assign _0608_ = _0602_ & ~_0601_;
	assign _0609_ = _0605_ | _0608_;
	assign _0611_ = _0607_ & ~_0609_;
	assign _0612_ = _0405_ & ~_0406_;
	assign _0613_ = _0419_ & ~_0420_;
	assign _0614_ = ~(_0406_ ^ _0405_);
	assign _0615_ = _0614_ & _0613_;
	assign _0616_ = _0615_ | _0612_;
	assign _0617_ = _0448_ | ~_0449_;
	assign _0618_ = ~(_0617_ | _0594_);
	assign _0619_ = _0430_ & ~_0431_;
	assign _0620_ = ~(_0619_ | _0618_);
	assign _0622_ = ~(_0420_ ^ _0419_);
	assign _0623_ = ~(_0622_ & _0614_);
	assign _0624_ = ~(_0623_ | _0620_);
	assign _0625_ = _0624_ | _0616_;
	assign _0626_ = _0458_ & ~_0459_;
	assign _0627_ = _0472_ | ~_0473_;
	assign _0628_ = ~(_0627_ | _0490_);
	assign _0629_ = _0628_ | _0626_;
	assign _0630_ = _0483_ & ~_0484_;
	assign _0631_ = ~(_0502_ | _0501_);
	assign _0633_ = _0631_ & ~_0589_;
	assign _0634_ = _0633_ | _0630_;
	assign _0635_ = _0490_ | ~_0486_;
	assign _0636_ = _0634_ & ~_0635_;
	assign _0637_ = _0636_ | _0629_;
	assign _0638_ = _0594_ | ~_0461_;
	assign _0639_ = _0638_ | _0623_;
	assign _0640_ = _0637_ & ~_0639_;
	assign _0642_ = _0640_ | _0625_;
	assign _0643_ = ~(_0396_ ^ _0395_);
	assign _0644_ = _0602_ ^ _0601_;
	assign _0645_ = ~(_0644_ & _0643_);
	assign _0646_ = _0642_ & ~_0645_;
	assign _0647_ = _0602_ & _0601_;
	assign _0648_ = _0395_ & ~_0396_;
	assign _0649_ = _0644_ & _0648_;
	assign _0650_ = _0649_ | _0647_;
	assign _0651_ = ~(_0650_ | _0646_);
	assign _0653_ = ~(_0651_ & _0605_);
	assign _0654_ = (_0790_ ? _0611_ : _0653_);
	assign _0655_ = (_0233_ ? _0342_ : _0654_);
	assign _0656_ = _0195_ & ~_0588_;
	assign _0657_ = (_0280_ ? _2551_ : _0555_);
	assign _0658_ = ~_0361_;
	assign _0659_ = (_0233_ ? _0657_ : _0658_);
	assign _0660_ = (_0280_ ? _2534_ : _0544_);
	assign _0661_ = (_0233_ ? _0660_ : _0357_);
	assign _0662_ = _0661_ & _0659_;
	assign _0664_ = (_0280_ ? _0217_ : _0522_);
	assign _0665_ = (_0233_ ? _0664_ : _0366_);
	assign _0666_ = (_0280_ ? _2567_ : _0511_);
	assign _0667_ = (_0233_ ? _0666_ : _0374_);
	assign _0668_ = _0667_ & ~_0665_;
	assign _0669_ = ~(_0668_ & _0662_);
	assign _0670_ = ~(_0669_ | _0656_);
	assign _0671_ = ~_0656_;
	assign _0672_ = _0667_ & _0665_;
	assign _0673_ = ~(_0672_ & _0662_);
	assign _0675_ = _0671_ & ~_0673_;
	assign _0676_ = _0675_ | _0670_;
	assign _0677_ = ~(_0326_ ^ _0270_);
	assign _0678_ = ~(_0270_ ^ _2499_);
	assign _0679_ = (_0790_ ? _0677_ : _0678_);
	assign _0680_ = ~_0589_;
	assign _0681_ = ~_0631_;
	assign _0682_ = (_0790_ ? _0587_ : _0681_);
	assign _0683_ = ~(_0682_ ^ _0680_);
	assign _0685_ = (_0233_ ? _0679_ : _0683_);
	assign _0686_ = _0685_ & ~_0676_;
	assign _0687_ = ~_0686_;
	assign _0688_ = _0315_ ^ _0141_;
	assign _0689_ = ~_0688_;
	assign _0690_ = ~_0584_;
	assign _0691_ = _0578_ & ~_0583_;
	assign _0692_ = _0691_ ^ _0584_;
	assign _0693_ = (_0790_ ? _0692_ : _0690_);
	assign _0694_ = (_0233_ ? _0689_ : _0693_);
	assign _0696_ = _0244_ & _2274_;
	assign _0697_ = _0696_ | _2179_;
	assign _0698_ = _1373_ & ~_0253_;
	assign _0699_ = ~(_0698_ | _1893_);
	assign _0700_ = ~(_0248_ & _0244_);
	assign _0701_ = ~(_0700_ | _0699_);
	assign _0702_ = _0701_ | _0697_;
	assign _0703_ = _1950_ & ~_0263_;
	assign _0704_ = _0703_ | _1922_;
	assign _0706_ = _2499_ & ~_0270_;
	assign _0707_ = ~(_0706_ | _2020_);
	assign _0708_ = _0267_ & ~_0263_;
	assign _0709_ = _0708_ & ~_0707_;
	assign _0710_ = _0709_ | _0704_;
	assign _0711_ = _0253_ | ~_0258_;
	assign _0712_ = _0711_ | _0700_;
	assign _0713_ = _0710_ & ~_0712_;
	assign _0715_ = _0713_ | _0702_;
	assign _0716_ = ~(_0241_ & _0234_);
	assign _0717_ = _0715_ & ~_0716_;
	assign _0718_ = _0234_ & _2131_;
	assign _0719_ = _0718_ | _2138_;
	assign _0720_ = _0719_ | _0717_;
	assign _0721_ = (_0790_ ? _0341_ : _0720_);
	assign _0722_ = ~(_0603_ & _0598_);
	assign _0723_ = _0608_ | ~_0722_;
	assign _0725_ = (_0790_ ? _0723_ : _0651_);
	assign _0726_ = ~(_0725_ ^ _0605_);
	assign _0727_ = (_0233_ ? _0721_ : _0726_);
	assign _0728_ = _0338_ | _0241_;
	assign _0729_ = _0728_ & ~_0284_;
	assign _0730_ = _0729_ ^ _0286_;
	assign _0731_ = _0241_ & _0715_;
	assign _0732_ = _2132_ & ~_0731_;
	assign _0733_ = _0732_ ^ _0235_;
	assign _0734_ = (_0790_ ? _0730_ : _0733_);
	assign _0736_ = _0603_ ^ _0598_;
	assign _0737_ = ~(_0643_ & _0642_);
	assign _0738_ = _0737_ & ~_0648_;
	assign _0739_ = ~(_0738_ ^ _0644_);
	assign _0740_ = (_0790_ ? _0736_ : _0739_);
	assign _0741_ = (_0233_ ? _0734_ : _0740_);
	assign _0742_ = _0656_ & ~_0661_;
	assign _0743_ = ~(_0667_ | _0659_);
	assign _0744_ = _0743_ & _0742_;
	assign _0745_ = ~_0790_;
	assign _0747_ = ~(_0583_ ^ _0578_);
	assign _0748_ = (_0790_ ? _0747_ : _0583_);
	assign _0749_ = _0233_ | ~_0748_;
	assign _0750_ = ~(_0749_ | _0744_);
	assign _0751_ = ~_0750_;
	assign _0752_ = _0338_ ^ _0241_;
	assign _0753_ = _0241_ ^ _0715_;
	assign _0754_ = (_0790_ ? _0752_ : _0753_);
	assign _0755_ = ~_0437_;
	assign _0756_ = _0593_ & ~_0595_;
	assign _0758_ = _0436_ & ~_0756_;
	assign _0759_ = _0758_ | _0755_;
	assign _0760_ = _0759_ & ~_0407_;
	assign _0761_ = ~(_0760_ ^ _0408_);
	assign _0762_ = _0643_ ^ _0642_;
	assign _0763_ = (_0790_ ? _0761_ : _0762_);
	assign _0764_ = (_0233_ ? _0754_ : _0763_);
	assign _0765_ = ~(_0661_ | _0659_);
	assign _0766_ = _0672_ | ~_0765_;
	assign _0767_ = _0656_ & ~_0766_;
	assign _0769_ = _0576_ ^ _0507_;
	assign _0770_ = (_0790_ ? _0769_ : _0507_);
	assign _0771_ = _0770_ | _0233_;
	assign _0772_ = ~(_0771_ | _0767_);
	assign _0773_ = ~_0772_;
	assign _0774_ = ~(_0334_ | _0259_);
	assign _0775_ = _0308_ & ~_0774_;
	assign _0776_ = _0775_ | _0248_;
	assign _0777_ = _0776_ & ~_0295_;
	assign _0778_ = _0777_ ^ _0297_;
	assign _0780_ = ~_0248_;
	assign _0781_ = _0710_ & ~_0711_;
	assign _0782_ = _0699_ & ~_0781_;
	assign _0783_ = _0782_ | _0780_;
	assign _0784_ = _0783_ & ~_2274_;
	assign _0785_ = ~(_0784_ ^ _0244_);
	assign _0786_ = (_0790_ ? _0778_ : _0785_);
	assign _0787_ = _0758_ ^ _0755_;
	assign _0788_ = ~_0622_;
	assign _0789_ = _0637_ & ~_0638_;
	assign _0791_ = _0620_ & ~_0789_;
	assign _0792_ = _0791_ | _0788_;
	assign _0793_ = _0792_ & ~_0613_;
	assign _0794_ = ~(_0793_ ^ _0614_);
	assign _0795_ = (_0790_ ? _0787_ : _0794_);
	assign _0796_ = (_0233_ ? _0786_ : _0795_);
	assign _0797_ = _0765_ & ~_0671_;
	assign _0798_ = _0233_ | ~_0576_;
	assign _0799_ = _0798_ | _0797_;
	assign _0800_ = _0799_ | ~_0796_;
	assign _0802_ = (_0764_ ? _0773_ : _0800_);
	assign _0803_ = (_0741_ ? _0751_ : _0802_);
	assign _0804_ = (_0727_ ? _0694_ : _0803_);
	assign _0805_ = (_0655_ ? _0687_ : _0804_);
	assign _0806_ = ~_0805_;
	assign _0807_ = ~(_0676_ | _0665_);
	assign _0808_ = ~(_0744_ | _0665_);
	assign _0809_ = _0665_ & ~_0767_;
	assign _0810_ = ~(_0797_ | _0665_);
	assign _0811_ = ~_0765_;
	assign _0813_ = _0659_ & ~_0661_;
	assign _0814_ = ~(_0667_ | _0665_);
	assign _0815_ = _0814_ & _0813_;
	assign _0816_ = _0811_ & ~_0815_;
	assign _0817_ = _0656_ & ~_0816_;
	assign _0818_ = _0665_ & ~_0817_;
	assign _0819_ = _0775_ ^ _0248_;
	assign _0820_ = _0782_ ^ _0780_;
	assign _0821_ = (_0790_ ? _0819_ : _0820_);
	assign _0822_ = ~(_0594_ & _0593_);
	assign _0824_ = _0822_ & ~_0432_;
	assign _0825_ = ~(_0824_ ^ _0433_);
	assign _0826_ = _0791_ ^ _0788_;
	assign _0827_ = (_0790_ ? _0825_ : _0826_);
	assign _0828_ = (_0233_ ? _0821_ : _0827_);
	assign _0829_ = _0667_ & _0659_;
	assign _0830_ = _0742_ & ~_0829_;
	assign _0831_ = ~(_0830_ | _0665_);
	assign _0832_ = ~(_0334_ | _0258_);
	assign _0833_ = _0302_ & ~_0832_;
	assign _0835_ = ~(_0833_ ^ _0253_);
	assign _0836_ = ~(_0258_ & _0710_);
	assign _0837_ = _0836_ & ~_1373_;
	assign _0838_ = _0837_ ^ _0253_;
	assign _0839_ = (_0790_ ? _0835_ : _0838_);
	assign _0840_ = _0594_ ^ _0593_;
	assign _0841_ = _0461_ & _0637_;
	assign _0842_ = _0617_ & ~_0841_;
	assign _0843_ = _0842_ ^ _0594_;
	assign _0844_ = (_0790_ ? _0840_ : _0843_);
	assign _0846_ = (_0233_ ? _0839_ : _0844_);
	assign _0847_ = _0813_ & ~_0672_;
	assign _0848_ = _0811_ & ~_0847_;
	assign _0849_ = _0656_ & ~_0848_;
	assign _0850_ = _0665_ & ~_0849_;
	assign _0851_ = _0334_ ^ _0258_;
	assign _0852_ = _0258_ ^ _0710_;
	assign _0853_ = (_0790_ ? _0851_ : _0852_);
	assign _0854_ = ~_0490_;
	assign _0855_ = _0587_ & ~_0590_;
	assign _0857_ = _0488_ & ~_0855_;
	assign _0858_ = _0857_ | _0854_;
	assign _0859_ = _0858_ & ~_0460_;
	assign _0860_ = _0859_ ^ _0461_;
	assign _0861_ = _0461_ ^ _0637_;
	assign _0862_ = (_0790_ ? _0860_ : _0861_);
	assign _0863_ = (_0233_ ? _0853_ : _0862_);
	assign _0864_ = ~(_0742_ | _0665_);
	assign _0865_ = _0331_ | _0267_;
	assign _0866_ = _0865_ & ~_0319_;
	assign _0868_ = _0267_ & ~_0707_;
	assign _0869_ = _0868_ | _1950_;
	assign _0870_ = (_0790_ ? _0866_ : _0869_);
	assign _0871_ = _0870_ ^ _0320_;
	assign _0872_ = _0857_ ^ _0854_;
	assign _0873_ = _0486_ & _0634_;
	assign _0874_ = _0627_ & ~_0873_;
	assign _0875_ = _0874_ ^ _0490_;
	assign _0876_ = (_0790_ ? _0872_ : _0875_);
	assign _0877_ = (_0233_ ? _0871_ : _0876_);
	assign _0879_ = _0659_ | ~_0661_;
	assign _0880_ = _0814_ & ~_0879_;
	assign _0881_ = _0661_ & ~_0880_;
	assign _0882_ = _0656_ & ~_0881_;
	assign _0883_ = _0665_ & ~_0882_;
	assign _0884_ = _0331_ ^ _0267_;
	assign _0885_ = ~(_0267_ ^ _0707_);
	assign _0886_ = (_0790_ ? _0884_ : _0885_);
	assign _0887_ = _0680_ | ~_0587_;
	assign _0888_ = _0887_ & ~_0485_;
	assign _0890_ = _0888_ ^ _0486_;
	assign _0891_ = _0486_ ^ _0634_;
	assign _0892_ = (_0790_ ? _0890_ : _0891_);
	assign _0893_ = (_0233_ ? _0886_ : _0892_);
	assign _0894_ = ~(_0661_ & _0656_);
	assign _0895_ = _0743_ & ~_0894_;
	assign _0896_ = ~(_0895_ | _0742_);
	assign _0897_ = _0896_ & ~_0665_;
	assign _0898_ = ~(_0879_ | _0672_);
	assign _0899_ = _0661_ & ~_0898_;
	assign _0901_ = _0656_ & ~_0899_;
	assign _0902_ = _0665_ & ~_0901_;
	assign _0903_ = _0656_ & ~_0662_;
	assign _0904_ = ~(_0903_ | _0665_);
	assign _0905_ = (_0694_ ? _0904_ : _0902_);
	assign _0906_ = (_0685_ ? _0897_ : _0905_);
	assign _0907_ = (_0893_ ? _0883_ : _0906_);
	assign _0908_ = (_0877_ ? _0864_ : _0907_);
	assign _0909_ = (_0863_ ? _0850_ : _0908_);
	assign _0910_ = (_0846_ ? _0831_ : _0909_);
	assign _0912_ = (_0828_ ? _0818_ : _0910_);
	assign _0913_ = (_0796_ ? _0810_ : _0912_);
	assign _0914_ = (_0764_ ? _0809_ : _0913_);
	assign _0915_ = (_0741_ ? _0808_ : _0914_);
	assign _0916_ = (_0727_ ? _0665_ : _0915_);
	assign _0917_ = (_0655_ ? _0807_ : _0916_);
	assign _0918_ = _0814_ | _0672_;
	assign _0919_ = _0918_ | _0676_;
	assign _0920_ = ~_0667_;
	assign _0921_ = _0744_ | ~_0918_;
	assign _0923_ = _0767_ | _0667_;
	assign _0924_ = _0918_ | _0797_;
	assign _0925_ = _0817_ | ~_0667_;
	assign _0926_ = _0830_ | ~_0918_;
	assign _0927_ = _0849_ | _0667_;
	assign _0928_ = _0918_ | _0742_;
	assign _0929_ = _0882_ | ~_0667_;
	assign _0930_ = ~(_0918_ & _0896_);
	assign _0931_ = _0901_ | _0667_;
	assign _0932_ = _0918_ | _0903_;
	assign _0934_ = (_0694_ ? _0932_ : _0931_);
	assign _0935_ = (_0685_ ? _0930_ : _0934_);
	assign _0936_ = (_0893_ ? _0929_ : _0935_);
	assign _0937_ = (_0877_ ? _0928_ : _0936_);
	assign _0938_ = (_0863_ ? _0927_ : _0937_);
	assign _0939_ = (_0846_ ? _0926_ : _0938_);
	assign _0940_ = (_0828_ ? _0925_ : _0939_);
	assign _0941_ = (_0796_ ? _0924_ : _0940_);
	assign _0942_ = (_0764_ ? _0923_ : _0941_);
	assign _0943_ = (_0741_ ? _0921_ : _0942_);
	assign _0945_ = (_0727_ ? _0920_ : _0943_);
	assign _0946_ = (_0655_ ? _0919_ : _0945_);
	assign _0947_ = ~(_0946_ | _0917_);
	assign _0948_ = ~_0659_;
	assign _0949_ = _0672_ & ~_0948_;
	assign _0950_ = _0948_ & ~_0672_;
	assign _0951_ = _0950_ | _0949_;
	assign _0952_ = ~(_0951_ | _0676_);
	assign _0953_ = _0814_ ^ _0948_;
	assign _0954_ = ~(_0953_ | _0744_);
	assign _0956_ = ~(_0829_ | _0743_);
	assign _0957_ = ~(_0956_ | _0767_);
	assign _0958_ = _0672_ ^ _0659_;
	assign _0959_ = ~(_0958_ | _0797_);
	assign _0960_ = ~(_0817_ | _0659_);
	assign _0961_ = _0659_ & ~_0814_;
	assign _0962_ = _0814_ & ~_0659_;
	assign _0963_ = _0962_ | _0961_;
	assign _0964_ = ~(_0963_ | _0830_);
	assign _0965_ = _0956_ & ~_0849_;
	assign _0967_ = ~(_0951_ | _0742_);
	assign _0968_ = _0659_ & ~_0882_;
	assign _0969_ = _0896_ & ~_0953_;
	assign _0970_ = ~(_0956_ | _0901_);
	assign _0971_ = ~(_0958_ | _0903_);
	assign _0972_ = (_0694_ ? _0971_ : _0970_);
	assign _0973_ = (_0685_ ? _0969_ : _0972_);
	assign _0974_ = (_0893_ ? _0968_ : _0973_);
	assign _0975_ = (_0877_ ? _0967_ : _0974_);
	assign _0976_ = (_0863_ ? _0965_ : _0975_);
	assign _0978_ = (_0846_ ? _0964_ : _0976_);
	assign _0979_ = (_0828_ ? _0960_ : _0978_);
	assign _0980_ = (_0796_ ? _0959_ : _0979_);
	assign _0981_ = (_0764_ ? _0957_ : _0980_);
	assign _0982_ = (_0741_ ? _0954_ : _0981_);
	assign _0983_ = (_0727_ ? _0659_ : _0982_);
	assign _0984_ = (_0655_ ? _0952_ : _0983_);
	assign _0985_ = ~_0661_;
	assign _0986_ = _0949_ ^ _0985_;
	assign _0987_ = ~(_0986_ | _0676_);
	assign _0989_ = ~_0987_;
	assign _0990_ = _0962_ ^ _0985_;
	assign _0991_ = ~(_0990_ | _0744_);
	assign _0992_ = ~_0991_;
	assign _0993_ = _0743_ ^ _0985_;
	assign _0994_ = ~(_0993_ | _0767_);
	assign _0995_ = ~_0994_;
	assign _0996_ = _0950_ ^ _0985_;
	assign _0997_ = ~(_0996_ | _0797_);
	assign _0998_ = ~_0997_;
	assign _1000_ = ~(_0765_ | _0662_);
	assign _1001_ = ~(_1000_ | _0817_);
	assign _1002_ = ~_1001_;
	assign _1003_ = _0961_ ^ _0661_;
	assign _1004_ = ~(_1003_ | _0830_);
	assign _1005_ = ~_1004_;
	assign _1006_ = _0829_ ^ _0661_;
	assign _1007_ = ~(_1006_ | _0849_);
	assign _1008_ = ~_1007_;
	assign _1009_ = _0949_ ^ _0661_;
	assign _1011_ = ~(_1009_ | _0742_);
	assign _1012_ = ~_1011_;
	assign _1013_ = _0671_ & ~_0661_;
	assign _1014_ = ~_1013_;
	assign _1015_ = _0962_ ^ _0661_;
	assign _1016_ = _0896_ & ~_1015_;
	assign _1017_ = ~_1016_;
	assign _1018_ = _0743_ & ~_0661_;
	assign _1019_ = _0661_ & ~_0743_;
	assign _1020_ = _1019_ | _1018_;
	assign _1022_ = ~(_1020_ | _0901_);
	assign _1023_ = ~_1022_;
	assign _1024_ = _0950_ ^ _0661_;
	assign _1025_ = ~(_1024_ | _0903_);
	assign _1026_ = ~_1025_;
	assign _1027_ = (_0694_ ? _1026_ : _1023_);
	assign _1028_ = (_0685_ ? _1017_ : _1027_);
	assign _1029_ = (_0893_ ? _1014_ : _1028_);
	assign _1030_ = (_0877_ ? _1012_ : _1029_);
	assign _1031_ = (_0863_ ? _1008_ : _1030_);
	assign _1033_ = (_0846_ ? _1005_ : _1031_);
	assign _1034_ = (_0828_ ? _1002_ : _1033_);
	assign _1035_ = (_0796_ ? _0998_ : _1034_);
	assign _1036_ = (_0764_ ? _0995_ : _1035_);
	assign _1037_ = (_0741_ ? _0992_ : _1036_);
	assign _1038_ = (_0727_ ? _0985_ : _1037_);
	assign _1039_ = (_0655_ ? _0989_ : _1038_);
	assign _1040_ = _1039_ | ~_0984_;
	assign _1041_ = _0947_ & ~_1040_;
	assign _1042_ = _0672_ & _0662_;
	assign _1044_ = _1042_ ^ _0656_;
	assign _1045_ = ~(_1044_ | _0676_);
	assign _1046_ = _0814_ & _0765_;
	assign _1047_ = _1046_ ^ _0656_;
	assign _1048_ = ~(_1047_ | _0744_);
	assign _1049_ = _1018_ ^ _0656_;
	assign _1050_ = ~(_1049_ | _0767_);
	assign _1051_ = _0765_ & ~_0672_;
	assign _1052_ = _1051_ ^ _0656_;
	assign _1053_ = ~(_1052_ | _0797_);
	assign _1055_ = _0671_ & ~_0765_;
	assign _1056_ = _0813_ & ~_0814_;
	assign _1057_ = _0985_ & ~_1056_;
	assign _1058_ = _1057_ ^ _0656_;
	assign _1059_ = ~(_1058_ | _0830_);
	assign _1060_ = _0985_ & ~_0829_;
	assign _1061_ = _1060_ ^ _0656_;
	assign _1062_ = ~(_1061_ | _0849_);
	assign _1063_ = _0813_ & _0672_;
	assign _1064_ = _0985_ & ~_1063_;
	assign _1066_ = _1064_ ^ _0656_;
	assign _1067_ = ~(_1066_ | _0742_);
	assign _1068_ = _0661_ & ~_0656_;
	assign _1069_ = ~_0896_;
	assign _1070_ = ~_0662_;
	assign _1071_ = ~(_0879_ | _0814_);
	assign _1072_ = _1070_ & ~_1071_;
	assign _1073_ = _1072_ ^ _0656_;
	assign _1074_ = ~(_1073_ | _1069_);
	assign _1075_ = _1019_ ^ _0671_;
	assign _1077_ = ~(_1075_ | _0901_);
	assign _1078_ = _0672_ & ~_0879_;
	assign _1079_ = _1070_ & ~_1078_;
	assign _1080_ = _1079_ ^ _0656_;
	assign _1081_ = ~(_1080_ | _0903_);
	assign _1082_ = (_0694_ ? _1081_ : _1077_);
	assign _1083_ = (_0685_ ? _1074_ : _1082_);
	assign _1084_ = (_0893_ ? _1068_ : _1083_);
	assign _1085_ = (_0877_ ? _1067_ : _1084_);
	assign _1086_ = (_0863_ ? _1062_ : _1085_);
	assign _1088_ = (_0846_ ? _1059_ : _1086_);
	assign _1089_ = (_0828_ ? _1055_ : _1088_);
	assign _1090_ = (_0796_ ? _1053_ : _1089_);
	assign _1091_ = (_0764_ ? _1050_ : _1090_);
	assign _1092_ = (_0741_ ? _1048_ : _1091_);
	assign _1093_ = (_0727_ ? _0671_ : _1092_);
	assign _1094_ = (_0655_ ? _1045_ : _1093_);
	assign _1095_ = ~_1094_;
	assign _1096_ = _1041_ & ~_1095_;
	assign _1097_ = _0946_ | ~_0917_;
	assign _1099_ = _1097_ | _1040_;
	assign _1100_ = _1094_ & ~_1099_;
	assign _1101_ = _1100_ | _1096_;
	assign _1102_ = _0676_ | ~_0893_;
	assign _1103_ = ~_0685_;
	assign _1104_ = _0694_ | _0744_;
	assign _1105_ = _0749_ | _0767_;
	assign _1106_ = _0771_ | _0797_;
	assign _1107_ = _0798_ | _0817_;
	assign _1108_ = _1107_ | ~_0828_;
	assign _1110_ = (_0796_ ? _1106_ : _1108_);
	assign _1111_ = (_0764_ ? _1105_ : _1110_);
	assign _1112_ = (_0741_ ? _1104_ : _1111_);
	assign _1113_ = (_0727_ ? _1103_ : _1112_);
	assign _1114_ = (_0655_ ? _1102_ : _1113_);
	assign _1115_ = ~(_0805_ ^ _1114_);
	assign _1116_ = _1115_ | _1101_;
	assign _1117_ = ~_0744_;
	assign _1118_ = ~_0767_;
	assign _1119_ = ~_0797_;
	assign _1121_ = ~_0817_;
	assign _1122_ = ~_0830_;
	assign _1123_ = ~_0849_;
	assign _1124_ = ~_0742_;
	assign _1125_ = ~_0882_;
	assign _1126_ = ~_0901_;
	assign _1127_ = ~(_0749_ | _0903_);
	assign _1128_ = (_0694_ ? _1127_ : _1126_);
	assign _1129_ = (_0685_ ? _0896_ : _1128_);
	assign _1130_ = (_0893_ ? _1125_ : _1129_);
	assign _1132_ = (_0877_ ? _1124_ : _1130_);
	assign _1133_ = (_0863_ ? _1123_ : _1132_);
	assign _1134_ = (_0846_ ? _1122_ : _1133_);
	assign _1135_ = (_0828_ ? _1121_ : _1134_);
	assign _1136_ = (_0796_ ? _1119_ : _1135_);
	assign _1137_ = (_0764_ ? _1118_ : _1136_);
	assign _1138_ = (_0741_ ? _1117_ : _1137_);
	assign _1139_ = ~(_1138_ | _0727_);
	assign _1140_ = (_0655_ ? _0676_ : _1139_);
	assign _1141_ = _0676_ | ~_0741_;
	assign _1143_ = ~_0764_;
	assign _1144_ = ~(_0796_ & _1117_);
	assign _1145_ = _0767_ | ~_0828_;
	assign _1146_ = ~(_0846_ & _1119_);
	assign _1147_ = _0817_ | ~_0863_;
	assign _1148_ = ~(_0877_ & _1122_);
	assign _1149_ = _0849_ | ~_0893_;
	assign _1150_ = ~(_0685_ & _1124_);
	assign _1151_ = _0694_ | _0882_;
	assign _1152_ = _0749_ | _1069_;
	assign _1154_ = _0771_ | _0901_;
	assign _1155_ = _0798_ | _0903_;
	assign _1156_ = (_0694_ ? _1155_ : _1154_);
	assign _1157_ = (_0685_ ? _1152_ : _1156_);
	assign _1158_ = (_0893_ ? _1151_ : _1157_);
	assign _1159_ = (_0877_ ? _1150_ : _1158_);
	assign _1160_ = (_0863_ ? _1149_ : _1159_);
	assign _1161_ = (_0846_ ? _1148_ : _1160_);
	assign _1162_ = (_0828_ ? _1147_ : _1161_);
	assign _1163_ = (_0796_ ? _1146_ : _1162_);
	assign _1165_ = (_0764_ ? _1145_ : _1163_);
	assign _1166_ = (_0741_ ? _1144_ : _1165_);
	assign _1167_ = (_0727_ ? _1143_ : _1166_);
	assign _1168_ = (_0655_ ? _1141_ : _1167_);
	assign _1169_ = _0676_ | ~_0727_;
	assign _1170_ = ~_0741_;
	assign _1171_ = _0744_ | ~_0764_;
	assign _1172_ = _0767_ | ~_0796_;
	assign _1173_ = _0797_ | ~_0828_;
	assign _1174_ = _0817_ | ~_0846_;
	assign _1176_ = ~(_0863_ & _1122_);
	assign _1177_ = _0849_ | ~_0877_;
	assign _1178_ = ~(_0893_ & _1124_);
	assign _1179_ = _0882_ | ~_0685_;
	assign _1180_ = _0694_ | _1069_;
	assign _1181_ = _0749_ | _0901_;
	assign _1182_ = _0771_ | _0903_;
	assign _1183_ = (_0694_ ? _1182_ : _1181_);
	assign _1184_ = (_0685_ ? _1180_ : _1183_);
	assign _1185_ = (_0893_ ? _1179_ : _1184_);
	assign _1187_ = (_0877_ ? _1178_ : _1185_);
	assign _1188_ = (_0863_ ? _1177_ : _1187_);
	assign _1189_ = (_0846_ ? _1176_ : _1188_);
	assign _1190_ = (_0828_ ? _1174_ : _1189_);
	assign _1191_ = (_0796_ ? _1173_ : _1190_);
	assign _1192_ = (_0764_ ? _1172_ : _1191_);
	assign _1193_ = (_0741_ ? _1171_ : _1192_);
	assign _1194_ = (_0727_ ? _1170_ : _1193_);
	assign _1195_ = (_0655_ ? _1169_ : _1194_);
	assign _1196_ = _1195_ | _1168_;
	assign _1198_ = ~(_0805_ | _1114_);
	assign _1199_ = _0877_ & ~_0676_;
	assign _1200_ = ~_1199_;
	assign _1201_ = ~_0893_;
	assign _1202_ = _0685_ & ~_0744_;
	assign _1203_ = ~_1202_;
	assign _1204_ = _1118_ & ~_0694_;
	assign _1205_ = ~_1204_;
	assign _1206_ = ~(_0749_ | _0797_);
	assign _1207_ = ~_1206_;
	assign _1209_ = ~(_0771_ | _0817_);
	assign _1210_ = ~_1209_;
	assign _1211_ = _0798_ | _0830_;
	assign _1212_ = _1211_ | ~_0846_;
	assign _1213_ = (_0828_ ? _1210_ : _1212_);
	assign _1214_ = (_0796_ ? _1207_ : _1213_);
	assign _1215_ = (_0764_ ? _1205_ : _1214_);
	assign _1216_ = (_0741_ ? _1203_ : _1215_);
	assign _1217_ = (_0727_ ? _1201_ : _1216_);
	assign _1218_ = (_0655_ ? _1200_ : _1217_);
	assign _1220_ = _0676_ | ~_0863_;
	assign _1221_ = ~_0877_;
	assign _1222_ = ~(_0893_ & _1117_);
	assign _1223_ = ~(_0685_ & _1118_);
	assign _1224_ = _0694_ | _0797_;
	assign _1225_ = _0749_ | _0817_;
	assign _1226_ = _0771_ | _0830_;
	assign _1227_ = _0798_ | _0849_;
	assign _1228_ = _1227_ | ~_0863_;
	assign _1229_ = (_0846_ ? _1226_ : _1228_);
	assign _1231_ = (_0828_ ? _1225_ : _1229_);
	assign _1232_ = (_0796_ ? _1224_ : _1231_);
	assign _1233_ = (_0764_ ? _1223_ : _1232_);
	assign _1234_ = (_0741_ ? _1222_ : _1233_);
	assign _1235_ = (_0727_ ? _1221_ : _1234_);
	assign _1236_ = (_0655_ ? _1220_ : _1235_);
	assign _1237_ = _1236_ | _1218_;
	assign _1238_ = _1198_ & ~_1237_;
	assign _1239_ = _0676_ | ~_0846_;
	assign _1240_ = ~_0863_;
	assign _1242_ = ~(_0877_ & _1117_);
	assign _1243_ = ~(_0893_ & _1118_);
	assign _1244_ = ~(_0685_ & _1119_);
	assign _1245_ = _0694_ | _0817_;
	assign _1246_ = _0749_ | _0830_;
	assign _1247_ = _0771_ | _0849_;
	assign _1248_ = _0798_ | _0742_;
	assign _1249_ = _1248_ | ~_0877_;
	assign _1250_ = (_0863_ ? _1247_ : _1249_);
	assign _1251_ = (_0846_ ? _1246_ : _1250_);
	assign _1253_ = (_0828_ ? _1245_ : _1251_);
	assign _1254_ = (_0796_ ? _1244_ : _1253_);
	assign _1255_ = (_0764_ ? _1243_ : _1254_);
	assign _1256_ = (_0741_ ? _1242_ : _1255_);
	assign _1257_ = (_0727_ ? _1240_ : _1256_);
	assign _1258_ = (_0655_ ? _1239_ : _1257_);
	assign _1259_ = _0676_ | ~_0828_;
	assign _1260_ = ~_0846_;
	assign _1261_ = ~(_0863_ & _1117_);
	assign _1262_ = ~(_0877_ & _1118_);
	assign _1264_ = ~(_0893_ & _1119_);
	assign _1265_ = _0817_ | ~_0685_;
	assign _1266_ = _0694_ | _0830_;
	assign _1267_ = _0749_ | _0849_;
	assign _1268_ = _0771_ | _0742_;
	assign _1269_ = _0798_ | _0882_;
	assign _1270_ = _1269_ | ~_0893_;
	assign _1271_ = (_0877_ ? _1268_ : _1270_);
	assign _1272_ = (_0863_ ? _1267_ : _1271_);
	assign _1273_ = (_0846_ ? _1266_ : _1272_);
	assign _1275_ = (_0828_ ? _1265_ : _1273_);
	assign _1276_ = (_0796_ ? _1264_ : _1275_);
	assign _1277_ = (_0764_ ? _1262_ : _1276_);
	assign _1278_ = (_0741_ ? _1261_ : _1277_);
	assign _1279_ = (_0727_ ? _1260_ : _1278_);
	assign _1280_ = (_0655_ ? _1259_ : _1279_);
	assign _1281_ = _1280_ | _1258_;
	assign _1282_ = _0796_ & ~_0676_;
	assign _1283_ = _0846_ & ~_0744_;
	assign _1284_ = ~(_0863_ & _1118_);
	assign _1286_ = ~_1284_;
	assign _1287_ = _0877_ & ~_0797_;
	assign _1288_ = ~(_0893_ & _1121_);
	assign _1289_ = ~_1288_;
	assign _1290_ = _0685_ & ~_0830_;
	assign _1291_ = ~(_0694_ | _0849_);
	assign _1292_ = ~(_0749_ | _0742_);
	assign _1293_ = ~(_0771_ | _0882_);
	assign _1294_ = _0798_ | _1069_;
	assign _1295_ = _0685_ & ~_1294_;
	assign _1297_ = (_0893_ ? _1293_ : _1295_);
	assign _1298_ = (_0877_ ? _1292_ : _1297_);
	assign _1299_ = (_0863_ ? _1291_ : _1298_);
	assign _1300_ = (_0846_ ? _1290_ : _1299_);
	assign _1301_ = (_0828_ ? _1289_ : _1300_);
	assign _1302_ = (_0796_ ? _1287_ : _1301_);
	assign _1303_ = (_0764_ ? _1286_ : _1302_);
	assign _1304_ = (_0741_ ? _1283_ : _1303_);
	assign _1305_ = (_0727_ ? _0828_ : _1304_);
	assign _1306_ = (_0655_ ? _1282_ : _1305_);
	assign _1308_ = _0676_ | ~_0764_;
	assign _1309_ = ~_0796_;
	assign _1310_ = _0744_ | ~_0828_;
	assign _1311_ = ~(_0846_ & _1118_);
	assign _1312_ = ~(_0863_ & _1119_);
	assign _1313_ = _0817_ | ~_0877_;
	assign _1314_ = ~(_0893_ & _1122_);
	assign _1315_ = _0849_ | ~_0685_;
	assign _1316_ = _0694_ | _0742_;
	assign _1317_ = _0749_ | _0882_;
	assign _1319_ = _0771_ | _1069_;
	assign _1320_ = _0798_ | _0901_;
	assign _1321_ = _1320_ | _0694_;
	assign _1322_ = (_0685_ ? _1319_ : _1321_);
	assign _1323_ = (_0893_ ? _1317_ : _1322_);
	assign _1324_ = (_0877_ ? _1316_ : _1323_);
	assign _1325_ = (_0863_ ? _1315_ : _1324_);
	assign _1326_ = (_0846_ ? _1314_ : _1325_);
	assign _1327_ = (_0828_ ? _1313_ : _1326_);
	assign _1328_ = (_0796_ ? _1312_ : _1327_);
	assign _1330_ = (_0764_ ? _1311_ : _1328_);
	assign _1331_ = (_0741_ ? _1310_ : _1330_);
	assign _1332_ = (_0727_ ? _1309_ : _1331_);
	assign _1333_ = (_0655_ ? _1308_ : _1332_);
	assign _1334_ = _1333_ | ~_1306_;
	assign _1335_ = ~(_1334_ | _1281_);
	assign _1336_ = ~(_1335_ & _1238_);
	assign _1337_ = _1336_ | _1196_;
	assign _1338_ = _1337_ | _1140_;
	assign _1339_ = (_1338_ ? _0806_ : _1116_);
	assign _1341_ = _0694_ | _0676_;
	assign _1342_ = _0771_ | _0744_;
	assign _1343_ = _0798_ | _0767_;
	assign _1344_ = _1343_ | ~_0764_;
	assign _1345_ = (_0741_ ? _1342_ : _1344_);
	assign _1346_ = (_0727_ ? _0749_ : _1345_);
	assign _1347_ = (_0655_ ? _1341_ : _1346_);
	assign _1348_ = ~(_0749_ | _0676_);
	assign _1349_ = ~_0771_;
	assign _1350_ = _0798_ | _0744_;
	assign _1352_ = _0741_ & ~_1350_;
	assign _1353_ = (_0727_ ? _1349_ : _1352_);
	assign _1354_ = (_0655_ ? _1348_ : _1353_);
	assign _1355_ = _0798_ & _0771_;
	assign _1356_ = ~(_1355_ | _0676_);
	assign _1357_ = _0727_ & ~_0798_;
	assign _1358_ = (_0655_ ? _1356_ : _1357_);
	assign _1359_ = _1358_ | _1354_;
	assign _1360_ = ~(_1359_ | _1347_);
	assign _1361_ = (_1360_ ? _0805_ : _1347_);
	assign _1363_ = (_1361_ ? _0805_ : _1339_);
	assign _1364_ = ~_0903_;
	assign _1365_ = (_0694_ ? _1364_ : _1126_);
	assign _1366_ = (_0685_ ? _0896_ : _1365_);
	assign _1367_ = (_0893_ ? _1125_ : _1366_);
	assign _1368_ = (_0877_ ? _1124_ : _1367_);
	assign _1369_ = (_0863_ ? _1123_ : _1368_);
	assign _1370_ = (_0846_ ? _1122_ : _1369_);
	assign _1371_ = (_0828_ ? _1121_ : _1370_);
	assign _1372_ = (_0796_ ? _1119_ : _1371_);
	assign _1374_ = (_0764_ ? _1118_ : _1372_);
	assign _1375_ = (_0741_ ? _1117_ : _1374_);
	assign _1376_ = ~(_1375_ | _0727_);
	assign _1377_ = (_0655_ ? _0676_ : _1376_);
	assign _1378_ = _1377_ | _1363_;
	assign _1379_ = (_0224_ ? _0223_ : _1378_);
	assign _1380_ = ~_0224_;
	assign _1381_ = ~(_0344_ | _0227_);
	assign _1382_ = ~(_1381_ & _0225_);
	assign _1384_ = ~(_0372_ & _0067_);
	assign _1385_ = _1384_ | _0339_;
	assign _1386_ = _1385_ | _1382_;
	assign _1387_ = _0688_ | ~_0270_;
	assign _1388_ = _1387_ | _0332_;
	assign _1389_ = _1388_ | _0335_;
	assign _1390_ = _1389_ | _1386_;
	assign _1391_ = _1390_ | _0745_;
	assign _1392_ = _1380_ & ~_1391_;
	assign _1394_ = _1392_ | _1379_;
	assign _1395_ = ~_0695_;
	assign _1396_ = ~_0195_;
	assign _1397_ = _2551_ | _2534_;
	assign _1398_ = _1397_ | _2568_;
	assign _1399_ = _1398_ | _1396_;
	assign _1400_ = _1395_ & ~_1399_;
	assign _1401_ = _1400_ | _1394_;
	assign _1402_ = ~(_1399_ | _0735_);
	assign _1403_ = (_1402_ ? _0823_ : _1401_);
	assign _1405_ = _0714_ | ~_0724_;
	assign _1406_ = ~(_1405_ | _1399_);
	assign _1407_ = (_1406_ ? _0823_ : _1403_);
	assign _1408_ = _0555_ | _0544_;
	assign _1409_ = _0522_ | _0511_;
	assign _1410_ = _1409_ | _1408_;
	assign _1411_ = _1410_ | _0588_;
	assign _1412_ = _1395_ & ~_1411_;
	assign _1413_ = _1412_ | _1407_;
	assign _1414_ = _1380_ & ~_1411_;
	assign _1416_ = (_1414_ ? _0812_ : _1413_);
	assign _1417_ = _1411_ | _1399_;
	assign _1418_ = ~(_1417_ | _0224_);
	assign _1419_ = _1418_ | _1416_;
	assign _1420_ = _0790_ & _0705_;
	assign _1421_ = _1420_ | _1419_;
	assign _1422_ = _0801_ & ~_1421_;
	assign _1423_ = _0641_ & ~_0224_;
	assign _1424_ = (_1423_ ? _0141_ : _1422_);
	assign _1425_ = _0652_ & ~_0224_;
	assign _1427_ = (_1425_ ? _0315_ : _1424_);
	assign _1428_ = ~(_0652_ & _0641_);
	assign _1429_ = _1428_ | ~_0790_;
	assign _1430_ = ~(_1429_ | _0224_);
	assign _1431_ = _1430_ | _1427_;
	assign _1432_ = _0621_ & ~_1431_;
	assign _1433_ = _2523_ & ~_1432_;
	assign _1434_ = ~_0621_;
	assign _1435_ = ~(_2480_ ^ _2476_);
	assign _1436_ = ~(_2480_ | _2476_);
	assign _1438_ = _1436_ ^ _2483_;
	assign _1439_ = (_2487_ ? _1438_ : _1435_);
	assign _1440_ = (_2524_ ? _2480_ : _1439_);
	assign _1441_ = _1440_ | _0200_;
	assign _1442_ = (_0220_ ? _1440_ : _1441_);
	assign _1443_ = _1442_ | _0222_;
	assign _1444_ = ~(_1336_ | _1168_);
	assign _1445_ = _1444_ ^ _1195_;
	assign _1446_ = _1445_ | _1101_;
	assign _1447_ = ~(_1336_ ^ _1168_);
	assign _1449_ = (_1338_ ? _1447_ : _1446_);
	assign _1450_ = (_1361_ ? _1168_ : _1449_);
	assign _1451_ = _1450_ | _1377_;
	assign _1452_ = (_0224_ ? _1443_ : _1451_);
	assign _1453_ = _1452_ | _1392_;
	assign _1454_ = _1453_ | _1400_;
	assign _1455_ = (_1402_ ? _2127_ : _1454_);
	assign _1456_ = (_1406_ ? _2127_ : _1455_);
	assign _1457_ = _1456_ | _1412_;
	assign _1458_ = (_1414_ ? _2114_ : _1457_);
	assign _1460_ = _1458_ | _1418_;
	assign _1461_ = _1460_ | _1420_;
	assign _1462_ = _0801_ & ~_1461_;
	assign _1463_ = (_1423_ ? _2544_ : _1462_);
	assign _1464_ = (_1425_ ? _0478_ : _1463_);
	assign _1465_ = _1464_ | _1430_;
	assign _1466_ = _1465_ | _1434_;
	assign _0008_ = (\mchip.in1.start  ? _1466_ : _1433_);
	assign _1467_ = ~_2443_;
	assign _1468_ = _2490_ ^ _2444_;
	assign _1470_ = (_2487_ ? _1468_ : _2488_);
	assign _1471_ = (_2524_ ? _1467_ : _1470_);
	assign _1472_ = _1471_ | _0200_;
	assign _1473_ = (_0220_ ? _1471_ : _1472_);
	assign _1474_ = _1473_ | _0222_;
	assign _1475_ = _1218_ ^ _1198_;
	assign _1476_ = _1475_ | _1101_;
	assign _1477_ = (_1338_ ? _1115_ : _1476_);
	assign _1478_ = (_1361_ ? _1114_ : _1477_);
	assign _1479_ = _1478_ | _1377_;
	assign _1481_ = (_0224_ ? _1474_ : _1479_);
	assign _1482_ = _1481_ | _1392_;
	assign _1483_ = _1482_ | _1400_;
	assign _1484_ = (_1402_ ? _2067_ : _1483_);
	assign _1485_ = (_1406_ ? _2067_ : _1484_);
	assign _1486_ = _1485_ | _1412_;
	assign _1487_ = (_1414_ ? _2260_ : _1486_);
	assign _1488_ = _1487_ | _1418_;
	assign _1489_ = _1488_ | _1420_;
	assign _1490_ = _0801_ & ~_1489_;
	assign _1492_ = (_1423_ ? _0130_ : _1490_);
	assign _1493_ = (_1425_ ? _0304_ : _1492_);
	assign _1494_ = _1493_ | _1430_;
	assign _1495_ = _0621_ & ~_1494_;
	assign _1496_ = _2523_ & ~_1495_;
	assign _1497_ = _1438_ | _2487_;
	assign _1498_ = (_2524_ ? _2483_ : _1497_);
	assign _1499_ = _1498_ | _0200_;
	assign _1500_ = (_0220_ ? _1498_ : _1499_);
	assign _1502_ = _1500_ | _0222_;
	assign _1503_ = ~(_1337_ ^ _1140_);
	assign _1504_ = _1503_ | _1101_;
	assign _1505_ = (_1338_ ? _1445_ : _1504_);
	assign _1506_ = (_1361_ ? _1195_ : _1505_);
	assign _1507_ = _1506_ | _1377_;
	assign _1508_ = (_0224_ ? _1502_ : _1507_);
	assign _1509_ = _1508_ | _1392_;
	assign _1510_ = _1509_ | _1400_;
	assign _1511_ = (_1402_ ? _2120_ : _1510_);
	assign _1513_ = (_1406_ ? _2120_ : _1511_);
	assign _1514_ = _1513_ | _1412_;
	assign _1515_ = (_1414_ ? _2113_ : _1514_);
	assign _1516_ = _1515_ | _1418_;
	assign _1517_ = _1516_ | _1420_;
	assign _1518_ = _0801_ & ~_1517_;
	assign _1519_ = (_1423_ ? _2533_ : _1518_);
	assign _1520_ = (_1425_ ? _0467_ : _1519_);
	assign _1521_ = _1520_ | _1430_;
	assign _1522_ = _1521_ | _1434_;
	assign _0009_ = (\mchip.in1.start  ? _1522_ : _1496_);
	assign _1524_ = _2444_ & ~_2490_;
	assign _1525_ = _1524_ ^ _2452_;
	assign _1526_ = (_2487_ ? _1525_ : _1468_);
	assign _1527_ = (_2524_ ? _2490_ : _1526_);
	assign _1528_ = _1527_ | _0200_;
	assign _1529_ = (_0220_ ? _1527_ : _1528_);
	assign _1530_ = _1529_ | _0222_;
	assign _1531_ = _1198_ & ~_1218_;
	assign _1532_ = _1531_ ^ _1236_;
	assign _1534_ = _1532_ | _1101_;
	assign _1535_ = (_1338_ ? _1475_ : _1534_);
	assign _1536_ = (_1361_ ? _1218_ : _1535_);
	assign _1537_ = _1536_ | _1377_;
	assign _1538_ = (_0224_ ? _1530_ : _1537_);
	assign _1539_ = _1538_ | _1392_;
	assign _1540_ = _1539_ | _1400_;
	assign _1541_ = (_1402_ ? _2364_ : _1540_);
	assign _1542_ = (_1406_ ? _2364_ : _1541_);
	assign _1543_ = _1542_ | _1412_;
	assign _1545_ = (_1414_ ? _2259_ : _1543_);
	assign _1546_ = _1545_ | _1418_;
	assign _1547_ = _1546_ | _1420_;
	assign _1548_ = _0801_ & ~_1547_;
	assign _1549_ = (_1423_ ? _0108_ : _1548_);
	assign _1550_ = (_1425_ ? _0347_ : _1549_);
	assign _1551_ = _1550_ | _1430_;
	assign _1552_ = _0621_ & ~_1551_;
	assign _1553_ = _2523_ & ~_1552_;
	assign _1554_ = _0211_ & ~_0200_;
	assign _1556_ = (_0220_ ? _0211_ : _1554_);
	assign _1557_ = _1556_ | _0222_;
	assign _1558_ = ~(_0655_ & _0676_);
	assign _1559_ = ~_0917_;
	assign _1560_ = _0917_ & ~_1101_;
	assign _1561_ = (_1338_ ? _1559_ : _1560_);
	assign _1562_ = (_1361_ ? _1559_ : _1561_);
	assign _1563_ = (_1377_ ? _1558_ : _1562_);
	assign _1564_ = (_0224_ ? _1557_ : _1563_);
	assign _1565_ = _1564_ | _1392_;
	assign _1567_ = _1565_ | _1400_;
	assign _1568_ = (_1402_ ? _0368_ : _1567_);
	assign _1569_ = (_1406_ ? _0368_ : _1568_);
	assign _1570_ = _1569_ | _1412_;
	assign _1571_ = (_1414_ ? _0367_ : _1570_);
	assign _1572_ = ~(_1571_ | _1418_);
	assign _1573_ = _1572_ | _1420_;
	assign _1574_ = _1573_ | ~_0801_;
	assign _1575_ = (_1423_ ? _0217_ : _1574_);
	assign _1576_ = (_1425_ ? _0522_ : _1575_);
	assign _1578_ = _1576_ | _1430_;
	assign _1579_ = _1578_ | _1434_;
	assign _0010_ = (\mchip.in1.start  ? _1579_ : _1553_);
	assign _1580_ = _2471_ ^ _2455_;
	assign _1581_ = (_2487_ ? _1580_ : _1525_);
	assign _1582_ = (_2524_ ? _2452_ : _1581_);
	assign _1583_ = _1582_ | _0200_;
	assign _1584_ = (_0220_ ? _1582_ : _1583_);
	assign _1585_ = _1584_ | _0222_;
	assign _1586_ = _1258_ ^ _1238_;
	assign _1588_ = _1586_ | _1101_;
	assign _1589_ = (_1338_ ? _1532_ : _1588_);
	assign _1590_ = (_1361_ ? _1236_ : _1589_);
	assign _1591_ = _1590_ | _1377_;
	assign _1592_ = (_0224_ ? _1585_ : _1591_);
	assign _1593_ = _1592_ | _1392_;
	assign _1594_ = _1593_ | _1400_;
	assign _1595_ = (_1402_ ? _2339_ : _1594_);
	assign _1596_ = (_1406_ ? _2339_ : _1595_);
	assign _1597_ = _1596_ | _1412_;
	assign _1599_ = (_1414_ ? _0312_ : _1597_);
	assign _1600_ = _1599_ | _1418_;
	assign _1601_ = _1600_ | _1420_;
	assign _1602_ = _0801_ & ~_1601_;
	assign _1603_ = (_1423_ ? _0097_ : _1602_);
	assign _1604_ = (_1425_ ? _0336_ : _1603_);
	assign _1605_ = _1604_ | _1430_;
	assign _1606_ = _0621_ & ~_1605_;
	assign _1607_ = _2523_ & ~_1606_;
	assign _1608_ = ~(_0211_ | _0209_);
	assign _1610_ = _1608_ | ~_0215_;
	assign _1611_ = ~(_1610_ | _0200_);
	assign _1612_ = (_0220_ ? _0209_ : _1611_);
	assign _1613_ = _1612_ | _0222_;
	assign _1614_ = ~(_0946_ ^ _0917_);
	assign _1615_ = ~(_1614_ | _1101_);
	assign _1616_ = (_1338_ ? _0946_ : _1615_);
	assign _1617_ = (_1361_ ? _0946_ : _1616_);
	assign _1618_ = (_1377_ ? _1558_ : _1617_);
	assign _1619_ = (_0224_ ? _1613_ : _1618_);
	assign _1621_ = _1619_ | _1392_;
	assign _1622_ = ~(_1621_ | _1400_);
	assign _1623_ = (_1402_ ? _0511_ : _1622_);
	assign _1624_ = (_1406_ ? _0511_ : _1623_);
	assign _1625_ = _1412_ | ~_1624_;
	assign _1626_ = (_1414_ ? _0206_ : _1625_);
	assign _1627_ = ~(_1626_ | _1418_);
	assign _1628_ = _1627_ | _1420_;
	assign _1629_ = _1628_ | ~_0801_;
	assign _1630_ = (_1423_ ? _2567_ : _1629_);
	assign _1632_ = (_1425_ ? _0511_ : _1630_);
	assign _1633_ = _1632_ | _1430_;
	assign _1634_ = _1633_ | _1434_;
	assign _0011_ = (\mchip.in1.start  ? _1634_ : _1607_);
	assign _1635_ = _2455_ & ~_2471_;
	assign _1636_ = _1635_ ^ _2473_;
	assign _1637_ = (_2487_ ? _1636_ : _1580_);
	assign _1638_ = (_2524_ ? _2471_ : _1637_);
	assign _1639_ = _1638_ | _0200_;
	assign _1640_ = (_0220_ ? _1638_ : _1639_);
	assign _1642_ = _1640_ | _0222_;
	assign _1643_ = _1238_ & ~_1258_;
	assign _1644_ = _1643_ ^ _1280_;
	assign _1645_ = _1644_ | _1101_;
	assign _1646_ = (_1338_ ? _1586_ : _1645_);
	assign _1647_ = (_1361_ ? _1258_ : _1646_);
	assign _1648_ = _1647_ | _1377_;
	assign _1649_ = (_0224_ ? _1642_ : _1648_);
	assign _1650_ = _1649_ | _1392_;
	assign _1651_ = _1650_ | _1400_;
	assign _1653_ = (_1402_ ? _2293_ : _1651_);
	assign _1654_ = (_1406_ ? _2293_ : _1653_);
	assign _1655_ = _1654_ | _1412_;
	assign _1656_ = (_1414_ ? _2187_ : _1655_);
	assign _1657_ = _1656_ | _1418_;
	assign _1658_ = _1657_ | _1420_;
	assign _1659_ = _0801_ & ~_1658_;
	assign _1660_ = (_1423_ ? _0064_ : _1659_);
	assign _1661_ = (_1425_ ? _0423_ : _1660_);
	assign _1662_ = _1661_ | _1430_;
	assign _1664_ = _0621_ & ~_1662_;
	assign _1665_ = _2523_ & ~_1664_;
	assign _1666_ = _1608_ ^ _0203_;
	assign _1667_ = ~(_1666_ | _0200_);
	assign _1668_ = (_0220_ ? _0203_ : _1667_);
	assign _1669_ = _1668_ | _0222_;
	assign _1670_ = ~_0984_;
	assign _1671_ = _1097_ ^ _1670_;
	assign _1672_ = ~(_1671_ | _1101_);
	assign _1673_ = (_1338_ ? _1670_ : _1672_);
	assign _1675_ = (_1361_ ? _1670_ : _1673_);
	assign _1676_ = (_1377_ ? _1558_ : _1675_);
	assign _1677_ = (_0224_ ? _1669_ : _1676_);
	assign _1678_ = _1677_ | _1392_;
	assign _1679_ = _1678_ | _1400_;
	assign _1680_ = (_1402_ ? _2545_ : _1679_);
	assign _1681_ = (_1406_ ? _2545_ : _1680_);
	assign _1682_ = _1681_ | _1412_;
	assign _1683_ = (_1414_ ? _0249_ : _1682_);
	assign _1684_ = ~(_1683_ | _1418_);
	assign _1686_ = _1684_ | _1420_;
	assign _1687_ = _1686_ | ~_0801_;
	assign _1688_ = (_1423_ ? _2551_ : _1687_);
	assign _1689_ = (_1425_ ? _0555_ : _1688_);
	assign _1690_ = _1689_ | _1430_;
	assign _1691_ = _1690_ | _1434_;
	assign _0012_ = (\mchip.in1.start  ? _1691_ : _1665_);
	assign _1692_ = ~_2460_;
	assign _1693_ = _2455_ & ~_2474_;
	assign _1694_ = _1693_ ^ _1692_;
	assign _1696_ = (_2487_ ? _1694_ : _1636_);
	assign _1697_ = (_2524_ ? _2473_ : _1696_);
	assign _1698_ = _1697_ | _0200_;
	assign _1699_ = (_0220_ ? _1697_ : _1698_);
	assign _1700_ = _1699_ | _0222_;
	assign _1701_ = ~_1306_;
	assign _1702_ = _1238_ & ~_1281_;
	assign _1703_ = _1702_ ^ _1701_;
	assign _1704_ = _1703_ | _1101_;
	assign _1705_ = (_1338_ ? _1644_ : _1704_);
	assign _1707_ = (_1361_ ? _1280_ : _1705_);
	assign _1708_ = _1707_ | _1377_;
	assign _1709_ = (_0224_ ? _1700_ : _1708_);
	assign _1710_ = _1709_ | _1392_;
	assign _1711_ = _1710_ | _1400_;
	assign _1712_ = (_1402_ ? _2240_ : _1711_);
	assign _1713_ = (_1406_ ? _2240_ : _1712_);
	assign _1714_ = _1713_ | _1412_;
	assign _1715_ = (_1414_ ? _2178_ : _1714_);
	assign _1716_ = _1715_ | _1418_;
	assign _1718_ = _1716_ | _1420_;
	assign _1719_ = _0801_ & ~_1718_;
	assign _1720_ = (_1423_ ? _2599_ : _1719_);
	assign _1721_ = (_1425_ ? _0412_ : _1720_);
	assign _1722_ = _1721_ | _1430_;
	assign _1723_ = _0621_ & ~_1722_;
	assign _1724_ = _2523_ & ~_1723_;
	assign _1725_ = _1608_ & ~_0203_;
	assign _1726_ = _1725_ ^ _0205_;
	assign _1727_ = ~(_1726_ | _0200_);
	assign _1729_ = (_0220_ ? _0205_ : _1727_);
	assign _1730_ = _1729_ | _0222_;
	assign _1731_ = _1097_ | _1670_;
	assign _1732_ = _1731_ ^ _1039_;
	assign _1733_ = ~(_1732_ | _1101_);
	assign _1734_ = (_1338_ ? _1039_ : _1733_);
	assign _1735_ = (_1361_ ? _1039_ : _1734_);
	assign _1736_ = (_1377_ ? _1558_ : _1735_);
	assign _1737_ = (_0224_ ? _1730_ : _1736_);
	assign _1738_ = _1737_ | _1392_;
	assign _1740_ = _1738_ | _1400_;
	assign _1741_ = (_1402_ ? _2543_ : _1740_);
	assign _1742_ = (_1406_ ? _2543_ : _1741_);
	assign _1743_ = _1742_ | _1412_;
	assign _1744_ = (_1414_ ? _0238_ : _1743_);
	assign _1745_ = ~(_1744_ | _1418_);
	assign _1746_ = _1745_ | _1420_;
	assign _1747_ = _1746_ | ~_0801_;
	assign _1748_ = (_1423_ ? _2534_ : _1747_);
	assign _1749_ = (_1425_ ? _0544_ : _1748_);
	assign _1751_ = _1749_ | _1430_;
	assign _1752_ = _1751_ | _1434_;
	assign _0013_ = (\mchip.in1.start  ? _1752_ : _1724_);
	assign _1753_ = _1693_ & ~_1692_;
	assign _1754_ = _1753_ ^ _2466_;
	assign _1755_ = (_2487_ ? _1754_ : _1694_);
	assign _1756_ = (_2524_ ? _1692_ : _1755_);
	assign _1757_ = _1756_ | _0200_;
	assign _1758_ = (_0220_ ? _1756_ : _1757_);
	assign _1759_ = _1758_ | _0222_;
	assign _1761_ = _1702_ & ~_1701_;
	assign _1762_ = _1761_ ^ _1333_;
	assign _1763_ = _1762_ | _1101_;
	assign _1764_ = (_1338_ ? _1703_ : _1763_);
	assign _1765_ = (_1361_ ? _1701_ : _1764_);
	assign _1766_ = _1765_ | _1377_;
	assign _1767_ = (_0224_ ? _1759_ : _1766_);
	assign _1768_ = _1767_ | _1392_;
	assign _1769_ = _1768_ | _1400_;
	assign _1770_ = (_1402_ ? _2196_ : _1769_);
	assign _1772_ = (_1406_ ? _2196_ : _1770_);
	assign _1773_ = _1772_ | _1412_;
	assign _1774_ = (_1414_ ? _2128_ : _1773_);
	assign _1775_ = _1774_ | _1418_;
	assign _1776_ = _1775_ | _1420_;
	assign _1777_ = _0801_ & ~_1776_;
	assign _1778_ = (_1423_ ? _2577_ : _1777_);
	assign _1779_ = (_1425_ ? _0390_ : _1778_);
	assign _1780_ = _1779_ | _1430_;
	assign _1781_ = _0621_ & ~_1780_;
	assign _1783_ = _2523_ & ~_1781_;
	assign _1784_ = _0205_ | _0203_;
	assign _1785_ = _1608_ & ~_1784_;
	assign _1786_ = _1785_ ^ _0181_;
	assign _1787_ = ~(_1786_ | _0200_);
	assign _1788_ = (_0220_ ? _0181_ : _1787_);
	assign _1789_ = _1788_ | _0222_;
	assign _1790_ = ~(_1097_ | _1040_);
	assign _1791_ = _1790_ ^ _1094_;
	assign _1792_ = ~(_1791_ | _1101_);
	assign _1794_ = (_1338_ ? _1095_ : _1792_);
	assign _1795_ = (_1361_ ? _1095_ : _1794_);
	assign _1796_ = (_1377_ ? _1558_ : _1795_);
	assign _1797_ = (_0224_ ? _1789_ : _1796_);
	assign _1798_ = _1797_ | _1392_;
	assign _1799_ = ~(_1798_ | _1400_);
	assign _1800_ = (_1402_ ? _0588_ : _1799_);
	assign _1801_ = (_1406_ ? _0588_ : _1800_);
	assign _1802_ = _1412_ | ~_1801_;
	assign _1803_ = (_1414_ ? _0195_ : _1802_);
	assign _1805_ = ~(_1803_ | _1418_);
	assign _1806_ = _1805_ | _1420_;
	assign _1807_ = _1806_ | ~_0801_;
	assign _1808_ = (_1423_ ? _1396_ : _1807_);
	assign _1809_ = (_1425_ ? _0588_ : _1808_);
	assign _1810_ = _1809_ | _1430_;
	assign _1811_ = _1810_ | _1434_;
	assign _0014_ = (\mchip.in1.start  ? _1811_ : _1783_);
	assign _1812_ = (_2487_ ? _1435_ : _1754_);
	assign _1813_ = (_2524_ ? _2466_ : _1812_);
	assign _1815_ = _1813_ | _0200_;
	assign _1816_ = (_0220_ ? _1813_ : _1815_);
	assign _1817_ = _1816_ | _0222_;
	assign _1818_ = _1447_ | _1101_;
	assign _1819_ = (_1338_ ? _1762_ : _1818_);
	assign _1820_ = (_1361_ ? _1333_ : _1819_);
	assign _1821_ = _1820_ | _1377_;
	assign _1822_ = (_0224_ ? _1817_ : _1821_);
	assign _1823_ = _1822_ | _1392_;
	assign _1824_ = _1823_ | _1400_;
	assign _1826_ = (_1402_ ? _2153_ : _1824_);
	assign _1827_ = (_1406_ ? _2153_ : _1826_);
	assign _1828_ = _1827_ | _1412_;
	assign _1829_ = (_1414_ ? _2115_ : _1828_);
	assign _1830_ = _1829_ | _1418_;
	assign _1831_ = _1830_ | _1420_;
	assign _1832_ = _0801_ & ~_1831_;
	assign _1833_ = (_1423_ ? _2566_ : _1832_);
	assign _1834_ = (_1425_ ? _0380_ : _1833_);
	assign _1835_ = _1834_ | _1430_;
	assign _1837_ = _0621_ & ~_1835_;
	assign _1838_ = _2523_ & ~_1837_;
	assign _1839_ = ~_0768_;
	assign _1840_ = ~_0779_;
	assign _1841_ = (_0280_ ? _1839_ : _1840_);
	assign _1842_ = (_0356_ ? _1839_ : _1840_);
	assign _1843_ = (_0233_ ? _1841_ : _1842_);
	assign _1844_ = _1843_ | ~_0676_;
	assign _1845_ = _1843_ | _1375_;
	assign _1846_ = _1845_ | _0727_;
	assign _1848_ = (_0655_ ? _1844_ : _1846_);
	assign _1849_ = (_1377_ ? _1848_ : _1843_);
	assign _1850_ = (_0224_ ? _0745_ : _1849_);
	assign _1851_ = _1850_ | _1392_;
	assign _1852_ = _1851_ | _1400_;
	assign _1853_ = (_1402_ ? _0779_ : _1852_);
	assign _1854_ = (_1406_ ? _1840_ : _1853_);
	assign _1855_ = _1854_ | _1412_;
	assign _1856_ = (_1414_ ? _1839_ : _1855_);
	assign _1857_ = ~(_1856_ | _1418_);
	assign _1859_ = (_0705_ ? _0790_ : _1857_);
	assign _1860_ = (_1423_ ? _0768_ : _1859_);
	assign _1861_ = (_1425_ ? _0779_ : _1860_);
	assign _1862_ = _1861_ | _1430_;
	assign _1863_ = _1862_ | _1434_;
	assign _0015_ = (\mchip.in1.start  ? _1863_ : _1838_);
	assign _0007_ = _2523_ | \mchip.in1.start ;
	assign io_out[1] = _0033_ & ~io_in[13];
	assign io_out[2] = _0034_ & ~io_in[13];
	assign io_out[3] = _0035_ & ~io_in[13];
	assign io_out[4] = _0036_ & ~io_in[13];
	assign io_out[5] = _0037_ & ~io_in[13];
	assign io_out[6] = _0038_ & ~io_in[13];
	assign io_out[7] = _0039_ & ~io_in[13];
	assign io_out[8] = _0040_ & ~io_in[13];
	assign io_out[9] = _0041_ & ~io_in[13];
	always @(posedge io_in[12])
		if (io_in[13])
			_0016_ <= 1'h0;
		else if (!_0000_)
			_0016_ <= _0006_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0017_ <= 1'h0;
		else if (_0003_)
			_0017_ <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0018_ <= 1'h0;
		else if (_0003_)
			_0018_ <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0019_ <= 1'h0;
		else if (_0003_)
			_0019_ <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0020_ <= 1'h0;
		else if (_0003_)
			_0020_ <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0021_ <= 1'h0;
		else if (_0003_)
			_0021_ <= io_in[6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0022_ <= 1'h0;
		else if (_0003_)
			_0022_ <= io_in[7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0023_ <= 1'h0;
		else if (_0003_)
			_0023_ <= io_in[8];
	always @(posedge io_in[12])
		if (io_in[13])
			_0024_ <= 1'h0;
		else if (_0003_)
			_0024_ <= io_in[9];
	always @(posedge io_in[12])
		if (io_in[13])
			_0025_ <= 1'h0;
		else if (_0005_)
			_0025_ <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0026_ <= 1'h0;
		else if (_0005_)
			_0026_ <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0027_ <= 1'h0;
		else if (_0005_)
			_0027_ <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0028_ <= 1'h0;
		else if (_0005_)
			_0028_ <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0029_ <= 1'h0;
		else if (_0005_)
			_0029_ <= io_in[6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0030_ <= 1'h0;
		else if (_0005_)
			_0030_ <= io_in[7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0031_ <= 1'h0;
		else if (_0005_)
			_0031_ <= io_in[8];
	always @(posedge io_in[12])
		if (io_in[13])
			_0032_ <= 1'h0;
		else if (_0005_)
			_0032_ <= io_in[9];
	always @(posedge io_in[12])
		if (io_in[13])
			_0033_ <= 1'h0;
		else
			_0033_ <= _0007_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0034_ <= 1'h0;
		else
			_0034_ <= _0008_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0035_ <= 1'h0;
		else
			_0035_ <= _0009_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0036_ <= 1'h0;
		else
			_0036_ <= _0010_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0037_ <= 1'h0;
		else
			_0037_ <= _0011_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0038_ <= 1'h0;
		else
			_0038_ <= _0012_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0039_ <= 1'h0;
		else
			_0039_ <= _0013_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0040_ <= 1'h0;
		else
			_0040_ <= _0014_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0041_ <= 1'h0;
		else
			_0041_ <= _0015_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0042_ <= 1'h0;
		else
			_0042_ <= \mchip.in1.start ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0043_ <= 1'h0;
		else if (_0004_)
			_0043_ <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0044_ <= 1'h0;
		else if (_0004_)
			_0044_ <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0045_ <= 1'h0;
		else if (_0004_)
			_0045_ <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0046_ <= 1'h0;
		else if (_0004_)
			_0046_ <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0047_ <= 1'h0;
		else if (_0004_)
			_0047_ <= io_in[6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0048_ <= 1'h0;
		else if (_0004_)
			_0048_ <= io_in[7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0049_ <= 1'h0;
		else if (_0004_)
			_0049_ <= io_in[8];
	always @(posedge io_in[12])
		if (io_in[13])
			_0050_ <= 1'h0;
		else if (_0004_)
			_0050_ <= io_in[9];
	always @(posedge io_in[12])
		if (io_in[13])
			_0051_ <= 1'h0;
		else if (_0002_)
			_0051_ <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0052_ <= 1'h0;
		else if (_0002_)
			_0052_ <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0053_ <= 1'h0;
		else if (_0002_)
			_0053_ <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0054_ <= 1'h0;
		else if (_0002_)
			_0054_ <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0055_ <= 1'h0;
		else if (_0002_)
			_0055_ <= io_in[6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0056_ <= 1'h0;
		else if (_0002_)
			_0056_ <= io_in[7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0057_ <= 1'h0;
		else if (_0002_)
			_0057_ <= io_in[8];
	always @(posedge io_in[12])
		if (io_in[13])
			_0058_ <= 1'h0;
		else if (_0002_)
			_0058_ <= io_in[9];
	always @(posedge io_in[12])
		if (io_in[13])
			_0059_ <= 1'h0;
		else if (_0001_)
			_0059_ <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0060_ <= 1'h0;
		else if (_0001_)
			_0060_ <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0061_ <= 1'h0;
		else if (_0001_)
			_0061_ <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0062_ <= 1'h0;
		else if (_0001_)
			_0062_ <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0063_ <= 1'h0;
		else if (_0000_)
			_0063_ <= _0001_;
	assign {io_out[13:10], io_out[0]} = {4'h0, io_out[1]};
	assign \mchip.calc.b [15] = 1'h0;
	assign \mchip.calc.max_exp  = 5'h1e;
	assign \mchip.calc.min_exp  = 5'h01;
	assign \mchip.clock  = io_in[12];
	assign \mchip.in1.clock  = io_in[12];
	assign \mchip.in1.data_in  = io_in[9:0];
	assign \mchip.in1.reset  = io_in[13];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {2'h0, io_out[9:1], io_out[1]};
	assign \mchip.out1.clock  = io_in[12];
	assign \mchip.out1.data_out  = {io_out[9:1], io_out[1]};
	assign \mchip.out1.done_calc  = \mchip.in1.start ;
	assign \mchip.out1.reset  = io_in[13];
	assign \mchip.reset  = io_in[13];
	assign \mchip.signal  = \mchip.in1.start ;
endmodule
`default_nettype none
module multiplexer (
	io_in,
	io_out,
	des_sel,
	hold_if_not_sel,
	sync_inputs,
	des_io_in,
	des_reset,
	des_io_out,
	clock,
	reset
);
	input wire [11:0] io_in;
	output reg [11:0] io_out;
	input wire [5:0] des_sel;
	input wire hold_if_not_sel;
	input wire sync_inputs;
	output reg [767:0] des_io_in;
	output reg [0:63] des_reset;
	input wire [767:0] des_io_out;
	input wire clock;
	input wire reset;
	reg [12:0] io_in_sync1;
	reg [12:0] io_in_sync2;
	reg [12:0] io_in_sync3;
	reg [63:0] des_sel_dec;
	always @(posedge clock) begin
		des_sel_dec <= 1'sb0;
		des_sel_dec[des_sel] <= 1;
		io_in_sync3 <= io_in_sync2;
		io_in_sync2 <= io_in_sync1;
		io_in_sync1 <= {reset, io_in};
	end
	integer i;
	always @(*) begin
		io_out = 1'sb0;
		for (i = 0; i < 64; i = i + 1)
			begin
				if (des_sel_dec[i])
					io_out = des_io_out[(63 - i) * 12+:12];
				if (hold_if_not_sel && !des_sel_dec[i]) begin
					des_io_in[(63 - i) * 12+:12] = 1'sb0;
					des_reset[i] = 1'sb1;
				end
				else begin
					des_io_in[(63 - i) * 12+:12] = (sync_inputs ? io_in_sync3[11:0] : io_in);
					des_reset[i] = (sync_inputs ? io_in_sync3[12] : reset);
				end
			end
	end
endmodule
`default_nettype none
module design_instantiations (
	io_in,
	io_out,
	des_sel,
	hold_if_not_sel,
	sync_inputs,
	clock,
	reset
);
	input wire [11:0] io_in;
	output wire [11:0] io_out;
	input wire [5:0] des_sel;
	input wire hold_if_not_sel;
	input wire sync_inputs;
	input wire clock;
	input wire reset;
	wire [767:0] des_io_in;
	wire [767:0] des_io_out;
	wire [0:63] des_reset;
	multiplexer mux(
		.io_in(io_in),
		.io_out(io_out),
		.des_sel(des_sel),
		.hold_if_not_sel(hold_if_not_sel),
		.sync_inputs(sync_inputs),
		.des_io_in(des_io_in),
		.des_reset(des_reset),
		.des_io_out(des_io_out),
		.clock(clock),
		.reset(reset)
	);
	assign des_io_out[756+:12] = 12'h000;
	d01_example_adder inst1(
		.io_in({des_reset[1], clock, des_io_in[744+:12]}),
		.io_out(des_io_out[744+:12])
	);
	d02_example_counter inst2(
		.io_in({des_reset[2], clock, des_io_in[732+:12]}),
		.io_out(des_io_out[732+:12])
	);
	d03_example_iotest inst3(
		.io_in({des_reset[3], clock, des_io_in[720+:12]}),
		.io_out(des_io_out[720+:12])
	);
	assign des_io_out[708+:12] = 12'h000;
	d05_meta_info inst5(
		.io_in({des_reset[5], clock, des_io_in[696+:12]}),
		.io_out(des_io_out[696+:12])
	);
	d06_demo_vgapong inst6(
		.io_in({des_reset[6], clock, des_io_in[684+:12]}),
		.io_out(des_io_out[684+:12])
	);
	d07_demo_vgarunner inst7(
		.io_in({des_reset[7], clock, des_io_in[672+:12]}),
		.io_out(des_io_out[672+:12])
	);
	assign des_io_out[660+:12] = 12'h000;
	assign des_io_out[648+:12] = 12'h000;
	d10_jjalacce_connect4 inst10(
		.io_in({des_reset[10], clock, des_io_in[636+:12]}),
		.io_out(des_io_out[636+:12])
	);
	d11_zhexic_i2cdriver inst11(
		.io_in({des_reset[11], clock, des_io_in[624+:12]}),
		.io_out(des_io_out[624+:12])
	);
	d12_sjg2_tiny_game_of_life inst12(
		.io_in({des_reset[12], clock, des_io_in[612+:12]}),
		.io_out(des_io_out[612+:12])
	);
	d13_thomaska_cordic inst13(
		.io_in({des_reset[13], clock, des_io_in[600+:12]}),
		.io_out(des_io_out[600+:12])
	);
	d14_siyuanl4_matrixcalc inst14(
		.io_in({des_reset[14], clock, des_io_in[588+:12]}),
		.io_out(des_io_out[588+:12])
	);
	d15_spencer2_pianotiles inst15(
		.io_in({des_reset[15], clock, des_io_in[576+:12]}),
		.io_out(des_io_out[576+:12])
	);
	d16_jaehyun3_bobatc inst16(
		.io_in({des_reset[16], clock, des_io_in[564+:12]}),
		.io_out(des_io_out[564+:12])
	);
	d17_cporco_clockbox inst17(
		.io_in({des_reset[17], clock, des_io_in[552+:12]}),
		.io_out(des_io_out[552+:12])
	);
	d18_vrajesh_motorcontroller inst18(
		.io_in({des_reset[18], clock, des_io_in[540+:12]}),
		.io_out(des_io_out[540+:12])
	);
	d19_gsavant_16bit_serial_cpu inst19(
		.io_in({des_reset[19], clock, des_io_in[528+:12]}),
		.io_out(des_io_out[528+:12])
	);
	d20_zhehuax_16bit_fpu inst20(
		.io_in({des_reset[20], clock, des_io_in[516+:12]}),
		.io_out(des_io_out[516+:12])
	);
	assign des_io_out[504+:12] = 12'h000;
	assign des_io_out[492+:12] = 12'h000;
	assign des_io_out[480+:12] = 12'h000;
	assign des_io_out[468+:12] = 12'h000;
	assign des_io_out[456+:12] = 12'h000;
	assign des_io_out[444+:12] = 12'h000;
	assign des_io_out[432+:12] = 12'h000;
	assign des_io_out[420+:12] = 12'h000;
	assign des_io_out[408+:12] = 12'h000;
	assign des_io_out[396+:12] = 12'h000;
	assign des_io_out[384+:12] = 12'h000;
	assign des_io_out[372+:12] = 12'h000;
	assign des_io_out[360+:12] = 12'h000;
	assign des_io_out[348+:12] = 12'h000;
	assign des_io_out[336+:12] = 12'h000;
	assign des_io_out[324+:12] = 12'h000;
	assign des_io_out[312+:12] = 12'h000;
	assign des_io_out[300+:12] = 12'h000;
	assign des_io_out[288+:12] = 12'h000;
	assign des_io_out[276+:12] = 12'h000;
	assign des_io_out[264+:12] = 12'h000;
	assign des_io_out[252+:12] = 12'h000;
	assign des_io_out[240+:12] = 12'h000;
	assign des_io_out[228+:12] = 12'h000;
	assign des_io_out[216+:12] = 12'h000;
	assign des_io_out[204+:12] = 12'h000;
	assign des_io_out[192+:12] = 12'h000;
	assign des_io_out[180+:12] = 12'h000;
	assign des_io_out[168+:12] = 12'h000;
	assign des_io_out[156+:12] = 12'h000;
	assign des_io_out[144+:12] = 12'h000;
	assign des_io_out[132+:12] = 12'h000;
	assign des_io_out[120+:12] = 12'h000;
	assign des_io_out[108+:12] = 12'h000;
	assign des_io_out[96+:12] = 12'h000;
	assign des_io_out[84+:12] = 12'h000;
	assign des_io_out[72+:12] = 12'h000;
	assign des_io_out[60+:12] = 12'h000;
	assign des_io_out[48+:12] = 12'h000;
	assign des_io_out[36+:12] = 12'h000;
	assign des_io_out[24+:12] = 12'h000;
	assign des_io_out[12+:12] = 12'h000;
	assign des_io_out[0+:12] = 12'h000;
endmodule
