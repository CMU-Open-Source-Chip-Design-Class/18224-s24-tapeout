module d01_example_adder (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire _07_;
	wire _08_;
	wire _09_;
	wire _10_;
	wire _11_;
	wire _12_;
	wire _13_;
	wire _14_;
	wire _15_;
	wire _16_;
	wire _17_;
	wire _18_;
	wire _19_;
	wire _20_;
	wire _21_;
	wire _22_;
	wire _23_;
	wire _24_;
	wire _25_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _00_ = io_in[5] ^ io_in[11];
	assign _01_ = ~(io_in[4] ^ io_in[10]);
	assign _02_ = _00_ & ~_01_;
	assign _03_ = ~(io_in[3] & io_in[9]);
	assign _04_ = io_in[3] ^ io_in[9];
	assign _05_ = ~(io_in[2] & io_in[8]);
	assign _06_ = _04_ & ~_05_;
	assign _07_ = _03_ & ~_06_;
	assign _08_ = ~(io_in[2] ^ io_in[8]);
	assign _09_ = _04_ & ~_08_;
	assign _10_ = ~(io_in[1] & io_in[7]);
	assign _11_ = io_in[1] ^ io_in[7];
	assign _12_ = ~(io_in[0] & io_in[6]);
	assign _13_ = _11_ & ~_12_;
	assign _14_ = _10_ & ~_13_;
	assign _15_ = _09_ & ~_14_;
	assign _16_ = _07_ & ~_15_;
	assign _17_ = _02_ & ~_16_;
	assign _18_ = ~(io_in[4] & io_in[10]);
	assign _19_ = _00_ & ~_18_;
	assign _20_ = io_in[5] & io_in[11];
	assign _21_ = _20_ | _19_;
	assign io_out[6] = _21_ | _17_;
	assign io_out[1] = ~(_12_ ^ _11_);
	assign io_out[2] = _14_ ^ _08_;
	assign _22_ = ~(_14_ | _08_);
	assign _23_ = _22_ | ~_05_;
	assign io_out[3] = _23_ ^ _04_;
	assign io_out[4] = _16_ ^ _01_;
	assign _24_ = ~(_16_ | _01_);
	assign _25_ = _24_ | ~_18_;
	assign io_out[5] = _25_ ^ _00_;
	assign io_out[0] = io_in[0] ^ io_in[6];
	assign io_out[13:7] = 7'h00;
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {5'h00, io_out[6:0]};
	assign \mchip.reset  = io_in[13];
endmodule
module d02_example_counter (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire [11:0] _059_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire \mchip.enable ;
	wire [11:0] \mchip.io_in ;
	reg [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire \mchip.updown ;
	assign _059_[0] = ~\mchip.io_out [0];
	assign _001_ = ~(io_in[1] & io_in[0]);
	assign _002_ = io_in[1] | ~io_in[0];
	assign _000_ = ~(_002_ & _001_);
	assign _003_ = _001_ ^ \mchip.io_out [1];
	assign _059_[1] = _003_ ^ _059_[0];
	assign _004_ = \mchip.io_out [1] & ~_001_;
	assign _005_ = \mchip.io_out [0] & ~_003_;
	assign _006_ = _005_ | _004_;
	assign _007_ = _001_ ^ \mchip.io_out [2];
	assign _059_[2] = ~(_007_ ^ _006_);
	assign _008_ = \mchip.io_out [2] & ~_001_;
	assign _009_ = _006_ & ~_007_;
	assign _010_ = ~(_009_ | _008_);
	assign _011_ = _001_ ^ \mchip.io_out [3];
	assign _059_[3] = _011_ ^ _010_;
	assign _012_ = _011_ | _007_;
	assign _013_ = _006_ & ~_012_;
	assign _014_ = \mchip.io_out [3] & ~_001_;
	assign _015_ = _008_ & ~_011_;
	assign _016_ = _015_ | _014_;
	assign _017_ = _016_ | _013_;
	assign _018_ = _001_ ^ \mchip.io_out [4];
	assign _059_[4] = ~(_018_ ^ _017_);
	assign _019_ = \mchip.io_out [4] & ~_001_;
	assign _020_ = _017_ & ~_018_;
	assign _021_ = ~(_020_ | _019_);
	assign _022_ = _001_ ^ \mchip.io_out [5];
	assign _059_[5] = _022_ ^ _021_;
	assign _023_ = _022_ | _018_;
	assign _024_ = _017_ & ~_023_;
	assign _025_ = \mchip.io_out [5] & ~_001_;
	assign _026_ = _019_ & ~_022_;
	assign _027_ = _026_ | _025_;
	assign _028_ = _027_ | _024_;
	assign _029_ = _001_ ^ \mchip.io_out [6];
	assign _059_[6] = ~(_029_ ^ _028_);
	assign _030_ = \mchip.io_out [6] & ~_001_;
	assign _031_ = _028_ & ~_029_;
	assign _032_ = ~(_031_ | _030_);
	assign _033_ = _001_ ^ \mchip.io_out [7];
	assign _059_[7] = _033_ ^ _032_;
	assign _034_ = \mchip.io_out [7] & ~_001_;
	assign _035_ = _030_ & ~_033_;
	assign _036_ = _035_ | _034_;
	assign _037_ = _033_ | _029_;
	assign _038_ = _027_ & ~_037_;
	assign _039_ = _038_ | _036_;
	assign _040_ = _037_ | _023_;
	assign _041_ = _017_ & ~_040_;
	assign _042_ = _041_ | _039_;
	assign _043_ = ~(_001_ ^ \mchip.io_out [8]);
	assign _059_[8] = _043_ ^ _042_;
	assign _044_ = \mchip.io_out [8] & ~_001_;
	assign _045_ = _043_ & _042_;
	assign _046_ = _045_ | _044_;
	assign _047_ = ~(_001_ ^ \mchip.io_out [9]);
	assign _059_[9] = _047_ ^ _046_;
	assign _048_ = \mchip.io_out [9] & ~_001_;
	assign _049_ = _047_ & _044_;
	assign _050_ = _049_ | _048_;
	assign _051_ = ~(_047_ & _043_);
	assign _052_ = _042_ & ~_051_;
	assign _053_ = _052_ | _050_;
	assign _054_ = ~(_001_ ^ \mchip.io_out [10]);
	assign _059_[10] = _054_ ^ _053_;
	assign _055_ = \mchip.io_out [10] & ~_001_;
	assign _056_ = _054_ & _053_;
	assign _057_ = _056_ | _055_;
	assign _058_ = ~(_001_ ^ \mchip.io_out [11]);
	assign _059_[11] = _058_ ^ _057_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [0] <= 1'h0;
		else if (_000_)
			\mchip.io_out [0] <= _059_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [1] <= 1'h0;
		else if (_000_)
			\mchip.io_out [1] <= _059_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [2] <= 1'h0;
		else if (_000_)
			\mchip.io_out [2] <= _059_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [3] <= 1'h0;
		else if (_000_)
			\mchip.io_out [3] <= _059_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [4] <= 1'h0;
		else if (_000_)
			\mchip.io_out [4] <= _059_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [5] <= 1'h0;
		else if (_000_)
			\mchip.io_out [5] <= _059_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [6] <= 1'h0;
		else if (_000_)
			\mchip.io_out [6] <= _059_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [7] <= 1'h0;
		else if (_000_)
			\mchip.io_out [7] <= _059_[7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [8] <= 1'h0;
		else if (_000_)
			\mchip.io_out [8] <= _059_[8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [9] <= 1'h0;
		else if (_000_)
			\mchip.io_out [9] <= _059_[9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [10] <= 1'h0;
		else if (_000_)
			\mchip.io_out [10] <= _059_[10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [11] <= 1'h0;
		else if (_000_)
			\mchip.io_out [11] <= _059_[11];
	assign io_out = {2'h0, \mchip.io_out };
	assign \mchip.clock  = io_in[12];
	assign \mchip.enable  = io_in[0];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.reset  = io_in[13];
	assign \mchip.updown  = io_in[1];
endmodule
module d05_meta_info (
	io_in,
	io_out
);
	wire _00000_;
	wire _00001_;
	wire _00002_;
	wire _00003_;
	wire _00004_;
	wire _00005_;
	wire _00006_;
	wire _00007_;
	wire _00008_;
	wire _00009_;
	wire _00010_;
	wire _00011_;
	wire _00012_;
	wire _00013_;
	wire _00014_;
	wire _00015_;
	wire _00016_;
	wire _00017_;
	wire _00018_;
	wire _00019_;
	wire _00020_;
	wire _00021_;
	wire _00022_;
	wire _00023_;
	wire _00024_;
	wire _00025_;
	wire _00026_;
	wire _00027_;
	wire _00028_;
	wire _00029_;
	wire _00030_;
	wire _00031_;
	wire _00032_;
	wire _00033_;
	wire _00034_;
	wire _00035_;
	wire _00036_;
	wire _00037_;
	wire _00038_;
	wire _00039_;
	wire _00040_;
	wire _00041_;
	wire _00042_;
	wire _00043_;
	wire _00044_;
	wire _00045_;
	wire _00046_;
	wire _00047_;
	wire _00048_;
	wire _00049_;
	wire _00050_;
	wire _00051_;
	wire _00052_;
	wire _00053_;
	wire _00054_;
	wire _00055_;
	wire _00056_;
	wire _00057_;
	wire _00058_;
	wire _00059_;
	wire _00060_;
	wire _00061_;
	wire _00062_;
	wire _00063_;
	wire _00064_;
	wire _00065_;
	wire _00066_;
	wire _00067_;
	wire _00068_;
	wire _00069_;
	wire _00070_;
	wire _00071_;
	wire _00072_;
	wire _00073_;
	wire _00074_;
	wire _00075_;
	wire _00076_;
	wire _00077_;
	wire _00078_;
	wire _00079_;
	wire _00080_;
	wire _00081_;
	wire _00082_;
	wire _00083_;
	wire _00084_;
	wire _00085_;
	wire _00086_;
	wire _00087_;
	wire _00088_;
	wire _00089_;
	wire _00090_;
	wire _00091_;
	wire _00092_;
	wire _00093_;
	wire _00094_;
	wire _00095_;
	wire _00096_;
	wire _00097_;
	wire _00098_;
	wire _00099_;
	wire _00100_;
	wire _00101_;
	wire _00102_;
	wire _00103_;
	wire _00104_;
	wire _00105_;
	wire _00106_;
	wire _00107_;
	wire _00108_;
	wire _00109_;
	wire _00110_;
	wire _00111_;
	wire _00112_;
	wire _00113_;
	wire _00114_;
	wire _00115_;
	wire _00116_;
	wire _00117_;
	wire _00118_;
	wire _00119_;
	wire _00120_;
	wire _00121_;
	wire _00122_;
	wire _00123_;
	wire _00124_;
	wire _00125_;
	wire _00126_;
	wire _00127_;
	wire _00128_;
	wire _00129_;
	wire _00130_;
	wire _00131_;
	wire _00132_;
	wire _00133_;
	wire _00134_;
	wire _00135_;
	wire _00136_;
	wire _00137_;
	wire _00138_;
	wire _00139_;
	wire _00140_;
	wire _00141_;
	wire _00142_;
	wire _00143_;
	wire _00144_;
	wire _00145_;
	wire _00146_;
	wire _00147_;
	wire _00148_;
	wire _00149_;
	wire _00150_;
	wire _00151_;
	wire _00152_;
	wire _00153_;
	wire _00154_;
	wire _00155_;
	wire _00156_;
	wire _00157_;
	wire _00158_;
	wire _00159_;
	wire _00160_;
	wire _00161_;
	wire _00162_;
	wire _00163_;
	wire _00164_;
	wire _00165_;
	wire _00166_;
	wire _00167_;
	wire _00168_;
	wire _00169_;
	wire _00170_;
	wire _00171_;
	wire _00172_;
	wire _00173_;
	wire _00174_;
	wire _00175_;
	wire _00176_;
	wire _00177_;
	wire _00178_;
	wire _00179_;
	wire _00180_;
	wire _00181_;
	wire _00182_;
	wire _00183_;
	wire _00184_;
	wire _00185_;
	wire _00186_;
	wire _00187_;
	wire _00188_;
	wire _00189_;
	wire _00190_;
	wire _00191_;
	wire _00192_;
	wire _00193_;
	wire _00194_;
	wire _00195_;
	wire _00196_;
	wire _00197_;
	wire _00198_;
	wire _00199_;
	wire _00200_;
	wire _00201_;
	wire _00202_;
	wire _00203_;
	wire _00204_;
	wire _00205_;
	wire _00206_;
	wire _00207_;
	wire _00208_;
	wire _00209_;
	wire _00210_;
	wire _00211_;
	wire _00212_;
	wire _00213_;
	wire _00214_;
	wire _00215_;
	wire _00216_;
	wire _00217_;
	wire _00218_;
	wire _00219_;
	wire _00220_;
	wire _00221_;
	wire _00222_;
	wire _00223_;
	wire _00224_;
	wire _00225_;
	wire _00226_;
	wire _00227_;
	wire _00228_;
	wire _00229_;
	wire _00230_;
	wire _00231_;
	wire _00232_;
	wire _00233_;
	wire _00234_;
	wire _00235_;
	wire _00236_;
	wire _00237_;
	wire _00238_;
	wire _00239_;
	wire _00240_;
	wire _00241_;
	wire _00242_;
	wire _00243_;
	wire _00244_;
	wire _00245_;
	wire _00246_;
	wire _00247_;
	wire _00248_;
	wire _00249_;
	wire _00250_;
	wire _00251_;
	wire _00252_;
	wire _00253_;
	wire _00254_;
	wire _00255_;
	wire _00256_;
	wire _00257_;
	wire _00258_;
	wire _00259_;
	wire _00260_;
	wire _00261_;
	wire _00262_;
	wire _00263_;
	wire _00264_;
	wire _00265_;
	wire _00266_;
	wire _00267_;
	wire _00268_;
	wire _00269_;
	wire _00270_;
	wire _00271_;
	wire _00272_;
	wire _00273_;
	wire _00274_;
	wire _00275_;
	wire _00276_;
	wire _00277_;
	wire _00278_;
	wire _00279_;
	wire _00280_;
	wire _00281_;
	wire _00282_;
	wire _00283_;
	wire _00284_;
	wire _00285_;
	wire _00286_;
	wire _00287_;
	wire _00288_;
	wire _00289_;
	wire _00290_;
	wire _00291_;
	wire _00292_;
	wire _00293_;
	wire _00294_;
	wire _00295_;
	wire _00296_;
	wire _00297_;
	wire _00298_;
	wire _00299_;
	wire _00300_;
	wire _00301_;
	wire _00302_;
	wire _00303_;
	wire _00304_;
	wire _00305_;
	wire _00306_;
	wire _00307_;
	wire _00308_;
	wire _00309_;
	wire _00310_;
	wire _00311_;
	wire _00312_;
	wire _00313_;
	wire _00314_;
	wire _00315_;
	wire _00316_;
	wire _00317_;
	wire _00318_;
	wire _00319_;
	wire _00320_;
	wire _00321_;
	wire _00322_;
	wire _00323_;
	wire _00324_;
	wire _00325_;
	wire _00326_;
	wire _00327_;
	wire _00328_;
	wire _00329_;
	wire _00330_;
	wire _00331_;
	wire _00332_;
	wire _00333_;
	wire _00334_;
	wire _00335_;
	wire _00336_;
	wire _00337_;
	wire _00338_;
	wire _00339_;
	wire _00340_;
	wire _00341_;
	wire _00342_;
	wire _00343_;
	wire _00344_;
	wire _00345_;
	wire _00346_;
	wire _00347_;
	wire _00348_;
	wire _00349_;
	wire _00350_;
	wire _00351_;
	wire _00352_;
	wire _00353_;
	wire _00354_;
	wire _00355_;
	wire _00356_;
	wire _00357_;
	wire _00358_;
	wire _00359_;
	wire _00360_;
	wire _00361_;
	wire _00362_;
	wire _00363_;
	wire _00364_;
	wire _00365_;
	wire _00366_;
	wire _00367_;
	wire _00368_;
	wire _00369_;
	wire _00370_;
	wire _00371_;
	wire _00372_;
	wire _00373_;
	wire _00374_;
	wire _00375_;
	wire _00376_;
	wire _00377_;
	wire _00378_;
	wire _00379_;
	wire _00380_;
	wire _00381_;
	wire _00382_;
	wire _00383_;
	wire _00384_;
	wire _00385_;
	wire _00386_;
	wire _00387_;
	wire _00388_;
	wire _00389_;
	wire _00390_;
	wire _00391_;
	wire _00392_;
	wire _00393_;
	wire _00394_;
	wire _00395_;
	wire _00396_;
	wire _00397_;
	wire _00398_;
	wire _00399_;
	wire _00400_;
	wire _00401_;
	wire _00402_;
	wire _00403_;
	wire _00404_;
	wire _00405_;
	wire _00406_;
	wire _00407_;
	wire _00408_;
	wire _00409_;
	wire _00410_;
	wire _00411_;
	wire _00412_;
	wire _00413_;
	wire _00414_;
	wire _00415_;
	wire _00416_;
	wire _00417_;
	wire _00418_;
	wire _00419_;
	wire _00420_;
	wire _00421_;
	wire _00422_;
	wire _00423_;
	wire _00424_;
	wire _00425_;
	wire _00426_;
	wire _00427_;
	wire _00428_;
	wire _00429_;
	wire _00430_;
	wire _00431_;
	wire _00432_;
	wire _00433_;
	wire _00434_;
	wire _00435_;
	wire _00436_;
	wire _00437_;
	wire _00438_;
	wire _00439_;
	wire _00440_;
	wire _00441_;
	wire _00442_;
	wire _00443_;
	wire _00444_;
	wire _00445_;
	wire _00446_;
	wire _00447_;
	wire _00448_;
	wire _00449_;
	wire _00450_;
	wire _00451_;
	wire _00452_;
	wire _00453_;
	wire _00454_;
	wire _00455_;
	wire _00456_;
	wire _00457_;
	wire _00458_;
	wire _00459_;
	wire _00460_;
	wire _00461_;
	wire _00462_;
	wire _00463_;
	wire _00464_;
	wire _00465_;
	wire _00466_;
	wire _00467_;
	wire _00468_;
	wire _00469_;
	wire _00470_;
	wire _00471_;
	wire _00472_;
	wire _00473_;
	wire _00474_;
	wire _00475_;
	wire _00476_;
	wire _00477_;
	wire _00478_;
	wire _00479_;
	wire _00480_;
	wire _00481_;
	wire _00482_;
	wire _00483_;
	wire _00484_;
	wire _00485_;
	wire _00486_;
	wire _00487_;
	wire _00488_;
	wire _00489_;
	wire _00490_;
	wire _00491_;
	wire _00492_;
	wire _00493_;
	wire _00494_;
	wire _00495_;
	wire _00496_;
	wire _00497_;
	wire _00498_;
	wire _00499_;
	wire _00500_;
	wire _00501_;
	wire _00502_;
	wire _00503_;
	wire _00504_;
	wire _00505_;
	wire _00506_;
	wire _00507_;
	wire _00508_;
	wire _00509_;
	wire _00510_;
	wire _00511_;
	wire _00512_;
	wire _00513_;
	wire _00514_;
	wire _00515_;
	wire _00516_;
	wire _00517_;
	wire _00518_;
	wire _00519_;
	wire _00520_;
	wire _00521_;
	wire _00522_;
	wire _00523_;
	wire _00524_;
	wire _00525_;
	wire _00526_;
	wire _00527_;
	wire _00528_;
	wire _00529_;
	wire _00530_;
	wire _00531_;
	wire _00532_;
	wire _00533_;
	wire _00534_;
	wire _00535_;
	wire _00536_;
	wire _00537_;
	wire _00538_;
	wire _00539_;
	wire _00540_;
	wire _00541_;
	wire _00542_;
	wire _00543_;
	wire _00544_;
	wire _00545_;
	wire _00546_;
	wire _00547_;
	wire _00548_;
	wire _00549_;
	wire _00550_;
	wire _00551_;
	wire _00552_;
	wire _00553_;
	wire _00554_;
	wire _00555_;
	wire _00556_;
	wire _00557_;
	wire _00558_;
	wire _00559_;
	wire _00560_;
	wire _00561_;
	wire _00562_;
	wire _00563_;
	wire _00564_;
	wire _00565_;
	wire _00566_;
	wire _00567_;
	wire _00568_;
	wire _00569_;
	wire _00570_;
	wire _00571_;
	wire _00572_;
	wire _00573_;
	wire _00574_;
	wire _00575_;
	wire _00576_;
	wire _00577_;
	wire _00578_;
	wire _00579_;
	wire _00580_;
	wire _00581_;
	wire _00582_;
	wire _00583_;
	wire _00584_;
	wire _00585_;
	wire _00586_;
	wire _00587_;
	wire _00588_;
	wire _00589_;
	wire _00590_;
	wire _00591_;
	wire _00592_;
	wire _00593_;
	wire _00594_;
	wire _00595_;
	wire _00596_;
	wire _00597_;
	wire _00598_;
	wire _00599_;
	wire _00600_;
	wire _00601_;
	wire _00602_;
	wire _00603_;
	wire _00604_;
	wire _00605_;
	wire _00606_;
	wire _00607_;
	wire _00608_;
	wire _00609_;
	wire _00610_;
	wire _00611_;
	wire _00612_;
	wire _00613_;
	wire _00614_;
	wire _00615_;
	wire _00616_;
	wire _00617_;
	wire _00618_;
	wire _00619_;
	wire _00620_;
	wire _00621_;
	wire _00622_;
	wire _00623_;
	wire _00624_;
	wire _00625_;
	wire _00626_;
	wire _00627_;
	wire _00628_;
	wire _00629_;
	wire _00630_;
	wire _00631_;
	wire _00632_;
	wire _00633_;
	wire _00634_;
	wire _00635_;
	wire _00636_;
	wire _00637_;
	wire _00638_;
	wire _00639_;
	wire _00640_;
	wire _00641_;
	wire _00642_;
	wire _00643_;
	wire _00644_;
	wire _00645_;
	wire _00646_;
	wire _00647_;
	wire _00648_;
	wire _00649_;
	wire _00650_;
	wire _00651_;
	wire _00652_;
	wire _00653_;
	wire _00654_;
	wire _00655_;
	wire _00656_;
	wire _00657_;
	wire _00658_;
	wire _00659_;
	wire _00660_;
	wire _00661_;
	wire _00662_;
	wire _00663_;
	wire _00664_;
	wire _00665_;
	wire _00666_;
	wire _00667_;
	wire _00668_;
	wire _00669_;
	wire _00670_;
	wire _00671_;
	wire _00672_;
	wire _00673_;
	wire _00674_;
	wire _00675_;
	wire _00676_;
	wire _00677_;
	wire _00678_;
	wire _00679_;
	wire _00680_;
	wire _00681_;
	wire _00682_;
	wire _00683_;
	wire _00684_;
	wire _00685_;
	wire _00686_;
	wire _00687_;
	wire _00688_;
	wire _00689_;
	wire _00690_;
	wire _00691_;
	wire _00692_;
	wire _00693_;
	wire _00694_;
	wire _00695_;
	wire _00696_;
	wire _00697_;
	wire _00698_;
	wire _00699_;
	wire _00700_;
	wire _00701_;
	wire _00702_;
	wire _00703_;
	wire _00704_;
	wire _00705_;
	wire _00706_;
	wire _00707_;
	wire _00708_;
	wire _00709_;
	wire _00710_;
	wire _00711_;
	wire _00712_;
	wire _00713_;
	wire _00714_;
	wire _00715_;
	wire _00716_;
	wire _00717_;
	wire _00718_;
	wire _00719_;
	wire _00720_;
	wire _00721_;
	wire _00722_;
	wire _00723_;
	wire _00724_;
	wire _00725_;
	wire _00726_;
	wire _00727_;
	wire _00728_;
	wire _00729_;
	wire _00730_;
	wire _00731_;
	wire _00732_;
	wire _00733_;
	wire _00734_;
	wire _00735_;
	wire _00736_;
	wire _00737_;
	wire _00738_;
	wire _00739_;
	wire _00740_;
	wire _00741_;
	wire _00742_;
	wire _00743_;
	wire _00744_;
	wire _00745_;
	wire _00746_;
	wire _00747_;
	wire _00748_;
	wire _00749_;
	wire _00750_;
	wire _00751_;
	wire _00752_;
	wire _00753_;
	wire _00754_;
	wire _00755_;
	wire _00756_;
	wire _00757_;
	wire _00758_;
	wire _00759_;
	wire _00760_;
	wire _00761_;
	wire _00762_;
	wire _00763_;
	wire _00764_;
	wire _00765_;
	wire _00766_;
	wire _00767_;
	wire _00768_;
	wire _00769_;
	wire _00770_;
	wire _00771_;
	wire _00772_;
	wire _00773_;
	wire _00774_;
	wire _00775_;
	wire _00776_;
	wire _00777_;
	wire _00778_;
	wire _00779_;
	wire _00780_;
	wire _00781_;
	wire _00782_;
	wire _00783_;
	wire _00784_;
	wire _00785_;
	wire _00786_;
	wire _00787_;
	wire _00788_;
	wire _00789_;
	wire _00790_;
	wire _00791_;
	wire _00792_;
	wire _00793_;
	wire _00794_;
	wire _00795_;
	wire _00796_;
	wire _00797_;
	wire _00798_;
	wire _00799_;
	wire _00800_;
	wire _00801_;
	wire _00802_;
	wire _00803_;
	wire _00804_;
	wire _00805_;
	wire _00806_;
	wire _00807_;
	wire _00808_;
	wire _00809_;
	wire _00810_;
	wire _00811_;
	wire _00812_;
	wire _00813_;
	wire _00814_;
	wire _00815_;
	wire _00816_;
	wire _00817_;
	wire _00818_;
	wire _00819_;
	wire _00820_;
	wire _00821_;
	wire _00822_;
	wire _00823_;
	wire _00824_;
	wire _00825_;
	wire _00826_;
	wire _00827_;
	wire _00828_;
	wire _00829_;
	wire _00830_;
	wire _00831_;
	wire _00832_;
	wire _00833_;
	wire _00834_;
	wire _00835_;
	wire _00836_;
	wire _00837_;
	wire _00838_;
	wire _00839_;
	wire _00840_;
	wire _00841_;
	wire _00842_;
	wire _00843_;
	wire _00844_;
	wire _00845_;
	wire _00846_;
	wire _00847_;
	wire _00848_;
	wire _00849_;
	wire _00850_;
	wire _00851_;
	wire _00852_;
	wire _00853_;
	wire _00854_;
	wire _00855_;
	wire _00856_;
	wire _00857_;
	wire _00858_;
	wire _00859_;
	wire _00860_;
	wire _00861_;
	wire _00862_;
	wire _00863_;
	wire _00864_;
	wire _00865_;
	wire _00866_;
	wire _00867_;
	wire _00868_;
	wire _00869_;
	wire _00870_;
	wire _00871_;
	wire _00872_;
	wire _00873_;
	wire _00874_;
	wire _00875_;
	wire _00876_;
	wire _00877_;
	wire _00878_;
	wire _00879_;
	wire _00880_;
	wire _00881_;
	wire _00882_;
	wire _00883_;
	wire _00884_;
	wire _00885_;
	wire _00886_;
	wire _00887_;
	wire _00888_;
	wire _00889_;
	wire _00890_;
	wire _00891_;
	wire _00892_;
	wire _00893_;
	wire _00894_;
	wire _00895_;
	wire _00896_;
	wire _00897_;
	wire _00898_;
	wire _00899_;
	wire _00900_;
	wire _00901_;
	wire _00902_;
	wire _00903_;
	wire _00904_;
	wire _00905_;
	wire _00906_;
	wire _00907_;
	wire _00908_;
	wire _00909_;
	wire _00910_;
	wire _00911_;
	wire _00912_;
	wire _00913_;
	wire _00914_;
	wire _00915_;
	wire _00916_;
	wire _00917_;
	wire _00918_;
	wire _00919_;
	wire _00920_;
	wire _00921_;
	wire _00922_;
	wire _00923_;
	wire _00924_;
	wire _00925_;
	wire _00926_;
	wire _00927_;
	wire _00928_;
	wire _00929_;
	wire _00930_;
	wire _00931_;
	wire _00932_;
	wire _00933_;
	wire _00934_;
	wire _00935_;
	wire _00936_;
	wire _00937_;
	wire _00938_;
	wire _00939_;
	wire _00940_;
	wire _00941_;
	wire _00942_;
	wire _00943_;
	wire _00944_;
	wire _00945_;
	wire _00946_;
	wire _00947_;
	wire _00948_;
	wire _00949_;
	wire _00950_;
	wire _00951_;
	wire _00952_;
	wire _00953_;
	wire _00954_;
	wire _00955_;
	wire _00956_;
	wire _00957_;
	wire _00958_;
	wire _00959_;
	wire _00960_;
	wire _00961_;
	wire _00962_;
	wire _00963_;
	wire _00964_;
	wire _00965_;
	wire _00966_;
	wire _00967_;
	wire _00968_;
	wire _00969_;
	wire _00970_;
	wire _00971_;
	wire _00972_;
	wire _00973_;
	wire _00974_;
	wire _00975_;
	wire _00976_;
	wire _00977_;
	wire _00978_;
	wire _00979_;
	wire _00980_;
	wire _00981_;
	wire _00982_;
	wire _00983_;
	wire _00984_;
	wire _00985_;
	wire _00986_;
	wire _00987_;
	wire _00988_;
	wire _00989_;
	wire _00990_;
	wire _00991_;
	wire _00992_;
	wire _00993_;
	wire _00994_;
	wire _00995_;
	wire _00996_;
	wire _00997_;
	wire _00998_;
	wire _00999_;
	wire _01000_;
	wire _01001_;
	wire _01002_;
	wire _01003_;
	wire _01004_;
	wire _01005_;
	wire _01006_;
	wire _01007_;
	wire _01008_;
	wire _01009_;
	wire _01010_;
	wire _01011_;
	wire _01012_;
	wire _01013_;
	wire _01014_;
	wire _01015_;
	wire _01016_;
	wire _01017_;
	wire _01018_;
	wire _01019_;
	wire _01020_;
	wire _01021_;
	wire _01022_;
	wire _01023_;
	wire _01024_;
	wire _01025_;
	wire _01026_;
	wire _01027_;
	wire _01028_;
	wire _01029_;
	wire _01030_;
	wire _01031_;
	wire _01032_;
	wire _01033_;
	wire _01034_;
	wire _01035_;
	wire _01036_;
	wire _01037_;
	wire _01038_;
	wire _01039_;
	wire _01040_;
	wire _01041_;
	wire _01042_;
	wire _01043_;
	wire _01044_;
	wire _01045_;
	wire _01046_;
	wire _01047_;
	wire _01048_;
	wire _01049_;
	wire _01050_;
	wire _01051_;
	wire _01052_;
	wire _01053_;
	wire _01054_;
	wire _01055_;
	wire _01056_;
	wire _01057_;
	wire _01058_;
	wire _01059_;
	wire _01060_;
	wire _01061_;
	wire _01062_;
	wire _01063_;
	wire _01064_;
	wire _01065_;
	wire _01066_;
	wire _01067_;
	wire _01068_;
	wire _01069_;
	wire _01070_;
	wire _01071_;
	wire _01072_;
	wire _01073_;
	wire _01074_;
	wire _01075_;
	wire _01076_;
	wire _01077_;
	wire _01078_;
	wire _01079_;
	wire _01080_;
	wire _01081_;
	wire _01082_;
	wire _01083_;
	wire _01084_;
	wire _01085_;
	wire _01086_;
	wire _01087_;
	wire _01088_;
	wire _01089_;
	wire _01090_;
	wire _01091_;
	wire _01092_;
	wire _01093_;
	wire _01094_;
	wire _01095_;
	wire _01096_;
	wire _01097_;
	wire _01098_;
	wire _01099_;
	wire _01100_;
	wire _01101_;
	wire _01102_;
	wire _01103_;
	wire _01104_;
	wire _01105_;
	wire _01106_;
	wire _01107_;
	wire _01108_;
	wire _01109_;
	wire _01110_;
	wire _01111_;
	wire _01112_;
	wire _01113_;
	wire _01114_;
	wire _01115_;
	wire _01116_;
	wire _01117_;
	wire _01118_;
	wire _01119_;
	wire _01120_;
	wire _01121_;
	wire _01122_;
	wire _01123_;
	wire _01124_;
	wire _01125_;
	wire _01126_;
	wire _01127_;
	wire _01128_;
	wire _01129_;
	wire _01130_;
	wire _01131_;
	wire _01132_;
	wire _01133_;
	wire _01134_;
	wire _01135_;
	wire _01136_;
	wire _01137_;
	wire _01138_;
	wire _01139_;
	wire _01140_;
	wire _01141_;
	wire _01142_;
	wire _01143_;
	wire _01144_;
	wire _01145_;
	wire _01146_;
	wire _01147_;
	wire _01148_;
	wire _01149_;
	wire _01150_;
	wire _01151_;
	wire _01152_;
	wire _01153_;
	wire _01154_;
	wire _01155_;
	wire _01156_;
	wire _01157_;
	wire _01158_;
	wire _01159_;
	wire _01160_;
	wire _01161_;
	wire _01162_;
	wire _01163_;
	wire _01164_;
	wire _01165_;
	wire _01166_;
	wire _01167_;
	wire _01168_;
	wire _01169_;
	wire _01170_;
	wire _01171_;
	wire _01172_;
	wire _01173_;
	wire _01174_;
	wire _01175_;
	wire _01176_;
	wire _01177_;
	wire _01178_;
	wire _01179_;
	wire _01180_;
	wire _01181_;
	wire _01182_;
	wire _01183_;
	wire _01184_;
	wire _01185_;
	wire _01186_;
	wire _01187_;
	wire _01188_;
	wire _01189_;
	wire _01190_;
	wire _01191_;
	wire _01192_;
	wire _01193_;
	wire _01194_;
	wire _01195_;
	wire _01196_;
	wire _01197_;
	wire _01198_;
	wire _01199_;
	wire _01200_;
	wire _01201_;
	wire _01202_;
	wire _01203_;
	wire _01204_;
	wire _01205_;
	wire _01206_;
	wire _01207_;
	wire _01208_;
	wire _01209_;
	wire _01210_;
	wire _01211_;
	wire _01212_;
	wire _01213_;
	wire _01214_;
	wire _01215_;
	wire _01216_;
	wire _01217_;
	wire _01218_;
	wire _01219_;
	wire _01220_;
	wire _01221_;
	wire _01222_;
	wire _01223_;
	wire _01224_;
	wire _01225_;
	wire _01226_;
	wire _01227_;
	wire _01228_;
	wire _01229_;
	wire _01230_;
	wire _01231_;
	wire _01232_;
	wire _01233_;
	wire _01234_;
	wire _01235_;
	wire _01236_;
	wire _01237_;
	wire _01238_;
	wire _01239_;
	wire _01240_;
	wire _01241_;
	wire _01242_;
	wire _01243_;
	wire _01244_;
	wire _01245_;
	wire _01246_;
	wire _01247_;
	wire _01248_;
	wire _01249_;
	wire _01250_;
	wire _01251_;
	wire _01252_;
	wire _01253_;
	wire _01254_;
	wire _01255_;
	wire _01256_;
	wire _01257_;
	wire _01258_;
	wire _01259_;
	wire _01260_;
	wire _01261_;
	wire _01262_;
	wire _01263_;
	wire _01264_;
	wire _01265_;
	wire _01266_;
	wire _01267_;
	wire _01268_;
	wire _01269_;
	wire _01270_;
	wire _01271_;
	wire _01272_;
	wire _01273_;
	wire _01274_;
	wire _01275_;
	wire _01276_;
	wire _01277_;
	wire _01278_;
	wire _01279_;
	wire _01280_;
	wire _01281_;
	wire _01282_;
	wire _01283_;
	wire _01284_;
	wire _01285_;
	wire _01286_;
	wire _01287_;
	wire _01288_;
	wire _01289_;
	wire _01290_;
	wire _01291_;
	wire _01292_;
	wire _01293_;
	wire _01294_;
	wire _01295_;
	wire _01296_;
	wire _01297_;
	wire _01298_;
	wire _01299_;
	wire _01300_;
	wire _01301_;
	wire _01302_;
	wire _01303_;
	wire _01304_;
	wire _01305_;
	wire _01306_;
	wire _01307_;
	wire _01308_;
	wire _01309_;
	wire _01310_;
	wire _01311_;
	wire _01312_;
	wire _01313_;
	wire _01314_;
	wire _01315_;
	wire _01316_;
	wire _01317_;
	wire _01318_;
	wire _01319_;
	wire _01320_;
	wire _01321_;
	wire _01322_;
	wire _01323_;
	wire _01324_;
	wire _01325_;
	wire _01326_;
	wire _01327_;
	wire _01328_;
	wire _01329_;
	wire _01330_;
	wire _01331_;
	wire _01332_;
	wire _01333_;
	wire _01334_;
	wire _01335_;
	wire _01336_;
	wire _01337_;
	wire _01338_;
	wire _01339_;
	wire _01340_;
	wire _01341_;
	wire _01342_;
	wire _01343_;
	wire _01344_;
	wire _01345_;
	wire _01346_;
	wire _01347_;
	wire _01348_;
	wire _01349_;
	wire _01350_;
	wire _01351_;
	wire _01352_;
	wire _01353_;
	wire _01354_;
	wire _01355_;
	wire _01356_;
	wire _01357_;
	wire _01358_;
	wire _01359_;
	wire _01360_;
	wire _01361_;
	wire _01362_;
	wire _01363_;
	wire _01364_;
	wire _01365_;
	wire _01366_;
	wire _01367_;
	wire _01368_;
	wire _01369_;
	wire _01370_;
	wire _01371_;
	wire _01372_;
	wire _01373_;
	wire _01374_;
	wire _01375_;
	wire _01376_;
	wire _01377_;
	wire _01378_;
	wire _01379_;
	wire _01380_;
	wire _01381_;
	wire _01382_;
	wire _01383_;
	wire _01384_;
	wire _01385_;
	wire _01386_;
	wire _01387_;
	wire _01388_;
	wire _01389_;
	wire _01390_;
	wire _01391_;
	wire _01392_;
	wire _01393_;
	wire _01394_;
	wire _01395_;
	wire _01396_;
	wire _01397_;
	wire _01398_;
	wire _01399_;
	wire _01400_;
	wire _01401_;
	wire _01402_;
	wire _01403_;
	wire _01404_;
	wire _01405_;
	wire _01406_;
	wire _01407_;
	wire _01408_;
	wire _01409_;
	wire _01410_;
	wire _01411_;
	wire _01412_;
	wire _01413_;
	wire _01414_;
	wire _01415_;
	wire _01416_;
	wire _01417_;
	wire _01418_;
	wire _01419_;
	wire _01420_;
	wire _01421_;
	wire _01422_;
	wire _01423_;
	wire _01424_;
	wire _01425_;
	wire _01426_;
	wire _01427_;
	wire _01428_;
	wire _01429_;
	wire _01430_;
	wire _01431_;
	wire _01432_;
	wire _01433_;
	wire _01434_;
	wire _01435_;
	wire _01436_;
	wire _01437_;
	wire _01438_;
	wire _01439_;
	wire _01440_;
	wire _01441_;
	wire _01442_;
	wire _01443_;
	wire _01444_;
	wire _01445_;
	wire _01446_;
	wire _01447_;
	wire _01448_;
	wire _01449_;
	wire _01450_;
	wire _01451_;
	wire _01452_;
	wire _01453_;
	wire _01454_;
	wire _01455_;
	wire _01456_;
	wire _01457_;
	wire _01458_;
	wire _01459_;
	wire _01460_;
	wire _01461_;
	wire _01462_;
	wire _01463_;
	wire _01464_;
	wire _01465_;
	wire _01466_;
	wire _01467_;
	wire _01468_;
	wire _01469_;
	wire _01470_;
	wire _01471_;
	wire _01472_;
	wire _01473_;
	wire _01474_;
	wire _01475_;
	wire _01476_;
	wire _01477_;
	wire _01478_;
	wire _01479_;
	wire _01480_;
	wire _01481_;
	wire _01482_;
	wire _01483_;
	wire _01484_;
	wire _01485_;
	wire _01486_;
	wire _01487_;
	wire _01488_;
	wire _01489_;
	wire _01490_;
	wire _01491_;
	wire _01492_;
	wire _01493_;
	wire _01494_;
	wire _01495_;
	wire _01496_;
	wire _01497_;
	wire _01498_;
	wire _01499_;
	wire _01500_;
	wire _01501_;
	wire _01502_;
	wire _01503_;
	wire _01504_;
	wire _01505_;
	wire _01506_;
	wire _01507_;
	wire _01508_;
	wire _01509_;
	wire _01510_;
	wire _01511_;
	wire _01512_;
	wire _01513_;
	wire _01514_;
	wire _01515_;
	wire _01516_;
	wire _01517_;
	wire _01518_;
	wire _01519_;
	wire _01520_;
	wire _01521_;
	wire _01522_;
	wire _01523_;
	wire _01524_;
	wire _01525_;
	wire _01526_;
	wire _01527_;
	wire _01528_;
	wire _01529_;
	wire _01530_;
	wire _01531_;
	wire _01532_;
	wire _01533_;
	wire _01534_;
	wire _01535_;
	wire _01536_;
	wire _01537_;
	wire _01538_;
	wire _01539_;
	wire _01540_;
	wire _01541_;
	wire _01542_;
	wire _01543_;
	wire _01544_;
	wire _01545_;
	wire _01546_;
	wire _01547_;
	wire _01548_;
	wire _01549_;
	wire _01550_;
	wire _01551_;
	wire _01552_;
	wire _01553_;
	wire _01554_;
	wire _01555_;
	wire _01556_;
	wire _01557_;
	wire _01558_;
	wire _01559_;
	wire _01560_;
	wire _01561_;
	wire _01562_;
	wire _01563_;
	wire _01564_;
	wire _01565_;
	wire _01566_;
	wire _01567_;
	wire _01568_;
	wire _01569_;
	wire _01570_;
	wire _01571_;
	wire _01572_;
	wire _01573_;
	wire _01574_;
	wire _01575_;
	wire _01576_;
	wire _01577_;
	wire _01578_;
	wire _01579_;
	wire _01580_;
	wire _01581_;
	wire _01582_;
	wire _01583_;
	wire _01584_;
	wire _01585_;
	wire _01586_;
	wire _01587_;
	wire _01588_;
	wire _01589_;
	wire _01590_;
	wire _01591_;
	wire _01592_;
	wire _01593_;
	wire _01594_;
	wire _01595_;
	wire _01596_;
	wire _01597_;
	wire _01598_;
	wire _01599_;
	wire _01600_;
	wire _01601_;
	wire _01602_;
	wire _01603_;
	wire _01604_;
	wire _01605_;
	wire _01606_;
	wire _01607_;
	wire _01608_;
	wire _01609_;
	wire _01610_;
	wire _01611_;
	wire _01612_;
	wire _01613_;
	wire _01614_;
	wire _01615_;
	wire _01616_;
	wire _01617_;
	wire _01618_;
	wire _01619_;
	wire _01620_;
	wire _01621_;
	wire _01622_;
	wire _01623_;
	wire _01624_;
	wire _01625_;
	wire _01626_;
	wire _01627_;
	wire _01628_;
	wire _01629_;
	wire _01630_;
	wire _01631_;
	wire _01632_;
	wire _01633_;
	wire _01634_;
	wire _01635_;
	wire _01636_;
	wire _01637_;
	wire _01638_;
	wire _01639_;
	wire _01640_;
	wire _01641_;
	wire _01642_;
	wire _01643_;
	wire _01644_;
	wire _01645_;
	wire _01646_;
	wire _01647_;
	wire _01648_;
	wire _01649_;
	wire _01650_;
	wire _01651_;
	wire _01652_;
	wire _01653_;
	wire _01654_;
	wire _01655_;
	wire _01656_;
	wire _01657_;
	wire _01658_;
	wire _01659_;
	wire _01660_;
	wire _01661_;
	wire _01662_;
	wire _01663_;
	wire _01664_;
	wire _01665_;
	wire _01666_;
	wire _01667_;
	wire _01668_;
	wire _01669_;
	wire _01670_;
	wire _01671_;
	wire _01672_;
	wire _01673_;
	wire _01674_;
	wire _01675_;
	wire _01676_;
	wire _01677_;
	wire _01678_;
	wire _01679_;
	wire _01680_;
	wire _01681_;
	wire _01682_;
	wire _01683_;
	wire _01684_;
	wire _01685_;
	wire _01686_;
	wire _01687_;
	wire _01688_;
	wire _01689_;
	wire _01690_;
	wire _01691_;
	wire _01692_;
	wire _01693_;
	wire _01694_;
	wire _01695_;
	wire _01696_;
	wire _01697_;
	wire _01698_;
	wire _01699_;
	wire _01700_;
	wire _01701_;
	wire _01702_;
	wire _01703_;
	wire _01704_;
	wire _01705_;
	wire _01706_;
	wire _01707_;
	wire _01708_;
	wire _01709_;
	wire _01710_;
	wire _01711_;
	wire _01712_;
	wire _01713_;
	wire _01714_;
	wire _01715_;
	wire _01716_;
	wire _01717_;
	wire _01718_;
	wire _01719_;
	wire _01720_;
	wire _01721_;
	wire _01722_;
	wire _01723_;
	wire _01724_;
	wire _01725_;
	wire _01726_;
	wire _01727_;
	wire _01728_;
	wire _01729_;
	wire _01730_;
	wire _01731_;
	wire _01732_;
	wire _01733_;
	wire _01734_;
	wire _01735_;
	wire _01736_;
	wire _01737_;
	wire _01738_;
	wire _01739_;
	wire _01740_;
	wire _01741_;
	wire _01742_;
	wire _01743_;
	wire _01744_;
	wire _01745_;
	wire _01746_;
	wire _01747_;
	wire _01748_;
	wire _01749_;
	wire _01750_;
	wire _01751_;
	wire _01752_;
	wire _01753_;
	wire _01754_;
	wire _01755_;
	wire _01756_;
	wire _01757_;
	wire _01758_;
	wire _01759_;
	wire _01760_;
	wire _01761_;
	wire _01762_;
	wire _01763_;
	wire _01764_;
	wire _01765_;
	wire _01766_;
	wire _01767_;
	wire _01768_;
	wire _01769_;
	wire _01770_;
	wire _01771_;
	wire _01772_;
	wire _01773_;
	wire _01774_;
	wire _01775_;
	wire _01776_;
	wire _01777_;
	wire _01778_;
	wire _01779_;
	wire _01780_;
	wire _01781_;
	wire _01782_;
	wire _01783_;
	wire _01784_;
	wire _01785_;
	wire _01786_;
	wire _01787_;
	wire _01788_;
	wire _01789_;
	wire _01790_;
	wire _01791_;
	wire _01792_;
	wire _01793_;
	wire _01794_;
	wire _01795_;
	wire _01796_;
	wire _01797_;
	wire _01798_;
	wire _01799_;
	wire _01800_;
	wire _01801_;
	wire _01802_;
	wire _01803_;
	wire _01804_;
	wire _01805_;
	wire _01806_;
	wire _01807_;
	wire _01808_;
	wire _01809_;
	wire _01810_;
	wire _01811_;
	wire _01812_;
	wire _01813_;
	wire _01814_;
	wire _01815_;
	wire _01816_;
	wire _01817_;
	wire _01818_;
	wire _01819_;
	wire _01820_;
	wire _01821_;
	wire _01822_;
	wire _01823_;
	wire _01824_;
	wire _01825_;
	wire _01826_;
	wire _01827_;
	wire _01828_;
	wire _01829_;
	wire _01830_;
	wire _01831_;
	wire _01832_;
	wire _01833_;
	wire _01834_;
	wire _01835_;
	wire _01836_;
	wire _01837_;
	wire _01838_;
	wire _01839_;
	wire _01840_;
	wire _01841_;
	wire _01842_;
	wire _01843_;
	wire _01844_;
	wire _01845_;
	wire _01846_;
	wire _01847_;
	wire _01848_;
	wire _01849_;
	wire _01850_;
	wire _01851_;
	wire _01852_;
	wire _01853_;
	wire _01854_;
	wire _01855_;
	wire _01856_;
	wire _01857_;
	wire _01858_;
	wire _01859_;
	wire _01860_;
	wire _01861_;
	wire _01862_;
	wire _01863_;
	wire _01864_;
	wire _01865_;
	wire _01866_;
	wire _01867_;
	wire _01868_;
	wire _01869_;
	wire _01870_;
	wire _01871_;
	wire _01872_;
	wire _01873_;
	wire _01874_;
	wire _01875_;
	wire _01876_;
	wire _01877_;
	wire _01878_;
	wire _01879_;
	wire _01880_;
	wire _01881_;
	wire _01882_;
	wire _01883_;
	wire _01884_;
	wire _01885_;
	wire _01886_;
	wire _01887_;
	wire _01888_;
	wire _01889_;
	wire _01890_;
	wire _01891_;
	wire _01892_;
	wire _01893_;
	wire _01894_;
	wire _01895_;
	wire _01896_;
	wire _01897_;
	wire _01898_;
	wire _01899_;
	wire _01900_;
	wire _01901_;
	wire _01902_;
	wire _01903_;
	wire _01904_;
	wire _01905_;
	wire _01906_;
	wire _01907_;
	wire _01908_;
	wire _01909_;
	wire _01910_;
	wire _01911_;
	wire _01912_;
	wire _01913_;
	wire _01914_;
	wire _01915_;
	wire _01916_;
	wire _01917_;
	wire _01918_;
	wire _01919_;
	wire _01920_;
	wire _01921_;
	wire _01922_;
	wire _01923_;
	wire _01924_;
	wire _01925_;
	wire _01926_;
	wire _01927_;
	wire _01928_;
	wire _01929_;
	wire _01930_;
	wire _01931_;
	wire _01932_;
	wire _01933_;
	wire _01934_;
	wire _01935_;
	wire _01936_;
	wire _01937_;
	wire _01938_;
	wire _01939_;
	wire _01940_;
	wire _01941_;
	wire _01942_;
	wire _01943_;
	wire _01944_;
	wire _01945_;
	wire _01946_;
	wire _01947_;
	wire _01948_;
	wire _01949_;
	wire _01950_;
	wire _01951_;
	wire _01952_;
	wire _01953_;
	wire _01954_;
	wire _01955_;
	wire _01956_;
	wire _01957_;
	wire _01958_;
	wire _01959_;
	wire _01960_;
	wire _01961_;
	wire _01962_;
	wire _01963_;
	wire _01964_;
	wire _01965_;
	wire _01966_;
	wire _01967_;
	wire _01968_;
	wire _01969_;
	wire _01970_;
	wire _01971_;
	wire _01972_;
	wire _01973_;
	wire _01974_;
	wire _01975_;
	wire _01976_;
	wire _01977_;
	wire _01978_;
	wire _01979_;
	wire _01980_;
	wire _01981_;
	wire _01982_;
	wire _01983_;
	wire _01984_;
	wire _01985_;
	wire _01986_;
	wire _01987_;
	wire _01988_;
	wire _01989_;
	wire _01990_;
	wire _01991_;
	wire _01992_;
	wire _01993_;
	wire _01994_;
	wire _01995_;
	wire _01996_;
	wire _01997_;
	wire _01998_;
	wire _01999_;
	wire _02000_;
	wire _02001_;
	wire _02002_;
	wire _02003_;
	wire _02004_;
	wire _02005_;
	wire _02006_;
	wire _02007_;
	wire _02008_;
	wire _02009_;
	wire _02010_;
	wire _02011_;
	wire _02012_;
	wire _02013_;
	wire _02014_;
	wire _02015_;
	wire _02016_;
	wire _02017_;
	wire _02018_;
	wire _02019_;
	wire _02020_;
	wire _02021_;
	wire _02022_;
	wire _02023_;
	wire _02024_;
	wire _02025_;
	wire _02026_;
	wire _02027_;
	wire _02028_;
	wire _02029_;
	wire _02030_;
	wire _02031_;
	wire _02032_;
	wire _02033_;
	wire _02034_;
	wire _02035_;
	wire _02036_;
	wire _02037_;
	wire _02038_;
	wire _02039_;
	wire _02040_;
	wire _02041_;
	wire _02042_;
	wire _02043_;
	wire _02044_;
	wire _02045_;
	wire _02046_;
	wire _02047_;
	wire _02048_;
	wire _02049_;
	wire _02050_;
	wire _02051_;
	wire _02052_;
	wire _02053_;
	wire _02054_;
	wire _02055_;
	wire _02056_;
	wire _02057_;
	wire _02058_;
	wire _02059_;
	wire _02060_;
	wire _02061_;
	wire _02062_;
	wire _02063_;
	wire _02064_;
	wire _02065_;
	wire _02066_;
	wire _02067_;
	wire _02068_;
	wire _02069_;
	wire _02070_;
	wire _02071_;
	wire _02072_;
	wire _02073_;
	wire _02074_;
	wire _02075_;
	wire _02076_;
	wire _02077_;
	wire _02078_;
	wire _02079_;
	wire _02080_;
	wire _02081_;
	wire _02082_;
	wire _02083_;
	wire _02084_;
	wire _02085_;
	wire _02086_;
	wire _02087_;
	wire _02088_;
	wire _02089_;
	wire _02090_;
	wire _02091_;
	wire _02092_;
	wire _02093_;
	wire _02094_;
	wire _02095_;
	wire _02096_;
	wire _02097_;
	wire _02098_;
	wire _02099_;
	wire _02100_;
	wire _02101_;
	wire _02102_;
	wire _02103_;
	wire _02104_;
	wire _02105_;
	wire _02106_;
	wire _02107_;
	wire _02108_;
	wire _02109_;
	wire _02110_;
	wire _02111_;
	wire _02112_;
	wire _02113_;
	wire _02114_;
	wire _02115_;
	wire _02116_;
	wire _02117_;
	wire _02118_;
	wire _02119_;
	wire _02120_;
	wire _02121_;
	wire _02122_;
	wire _02123_;
	wire _02124_;
	wire _02125_;
	wire _02126_;
	wire _02127_;
	wire _02128_;
	wire _02129_;
	wire _02130_;
	wire _02131_;
	wire _02132_;
	wire _02133_;
	wire _02134_;
	wire _02135_;
	wire _02136_;
	wire _02137_;
	wire _02138_;
	wire _02139_;
	wire _02140_;
	wire _02141_;
	wire _02142_;
	wire _02143_;
	wire _02144_;
	wire _02145_;
	wire _02146_;
	wire _02147_;
	wire _02148_;
	wire _02149_;
	wire _02150_;
	wire _02151_;
	wire _02152_;
	wire _02153_;
	wire _02154_;
	wire _02155_;
	wire _02156_;
	wire _02157_;
	wire _02158_;
	wire _02159_;
	wire _02160_;
	wire _02161_;
	wire _02162_;
	wire _02163_;
	wire _02164_;
	wire _02165_;
	wire _02166_;
	wire _02167_;
	wire _02168_;
	wire _02169_;
	wire _02170_;
	wire _02171_;
	wire _02172_;
	wire _02173_;
	wire _02174_;
	wire _02175_;
	wire _02176_;
	wire _02177_;
	wire _02178_;
	wire _02179_;
	wire _02180_;
	wire _02181_;
	wire _02182_;
	wire _02183_;
	wire _02184_;
	wire _02185_;
	wire _02186_;
	wire _02187_;
	wire _02188_;
	wire _02189_;
	wire _02190_;
	wire _02191_;
	wire _02192_;
	wire _02193_;
	wire _02194_;
	wire _02195_;
	wire _02196_;
	wire _02197_;
	wire _02198_;
	wire _02199_;
	wire _02200_;
	wire _02201_;
	wire _02202_;
	wire _02203_;
	wire _02204_;
	wire _02205_;
	wire _02206_;
	wire _02207_;
	wire _02208_;
	wire _02209_;
	wire _02210_;
	wire _02211_;
	wire _02212_;
	wire _02213_;
	wire _02214_;
	wire _02215_;
	wire _02216_;
	wire _02217_;
	wire _02218_;
	wire _02219_;
	wire _02220_;
	wire _02221_;
	wire _02222_;
	wire _02223_;
	wire _02224_;
	wire _02225_;
	wire _02226_;
	wire _02227_;
	wire _02228_;
	wire _02229_;
	wire _02230_;
	wire _02231_;
	wire _02232_;
	wire _02233_;
	wire _02234_;
	wire _02235_;
	wire _02236_;
	wire _02237_;
	wire _02238_;
	wire _02239_;
	wire _02240_;
	wire _02241_;
	wire _02242_;
	wire _02243_;
	wire _02244_;
	wire _02245_;
	wire _02246_;
	wire _02247_;
	wire _02248_;
	wire _02249_;
	wire _02250_;
	wire _02251_;
	wire _02252_;
	wire _02253_;
	wire _02254_;
	wire _02255_;
	wire _02256_;
	wire _02257_;
	wire _02258_;
	wire _02259_;
	wire _02260_;
	wire _02261_;
	wire _02262_;
	wire _02263_;
	wire _02264_;
	wire _02265_;
	wire _02266_;
	wire _02267_;
	wire _02268_;
	wire _02269_;
	wire _02270_;
	wire _02271_;
	wire _02272_;
	wire _02273_;
	wire _02274_;
	wire _02275_;
	wire _02276_;
	wire _02277_;
	wire _02278_;
	wire _02279_;
	wire _02280_;
	wire _02281_;
	wire _02282_;
	wire _02283_;
	wire _02284_;
	wire _02285_;
	wire _02286_;
	wire _02287_;
	wire _02288_;
	wire _02289_;
	wire _02290_;
	wire _02291_;
	wire _02292_;
	wire _02293_;
	wire _02294_;
	wire _02295_;
	wire _02296_;
	wire _02297_;
	wire _02298_;
	wire _02299_;
	wire _02300_;
	wire _02301_;
	wire _02302_;
	wire _02303_;
	wire _02304_;
	wire _02305_;
	wire _02306_;
	wire _02307_;
	wire _02308_;
	wire _02309_;
	wire _02310_;
	wire _02311_;
	wire _02312_;
	wire _02313_;
	wire _02314_;
	wire _02315_;
	wire _02316_;
	wire _02317_;
	wire _02318_;
	wire _02319_;
	wire _02320_;
	wire _02321_;
	wire _02322_;
	wire _02323_;
	wire _02324_;
	wire _02325_;
	wire _02326_;
	wire _02327_;
	wire _02328_;
	wire _02329_;
	wire _02330_;
	wire _02331_;
	wire _02332_;
	wire _02333_;
	wire _02334_;
	wire _02335_;
	wire _02336_;
	wire _02337_;
	wire _02338_;
	wire _02339_;
	wire _02340_;
	wire _02341_;
	wire _02342_;
	wire _02343_;
	wire _02344_;
	wire _02345_;
	wire _02346_;
	wire _02347_;
	wire _02348_;
	wire _02349_;
	wire _02350_;
	wire _02351_;
	wire _02352_;
	wire _02353_;
	wire _02354_;
	wire _02355_;
	wire _02356_;
	wire _02357_;
	wire _02358_;
	wire _02359_;
	wire _02360_;
	wire _02361_;
	wire _02362_;
	wire _02363_;
	wire _02364_;
	wire _02365_;
	wire _02366_;
	wire _02367_;
	wire _02368_;
	wire _02369_;
	wire _02370_;
	wire _02371_;
	wire _02372_;
	wire _02373_;
	wire _02374_;
	wire _02375_;
	wire _02376_;
	wire _02377_;
	wire _02378_;
	wire _02379_;
	wire _02380_;
	wire _02381_;
	wire _02382_;
	wire _02383_;
	wire _02384_;
	wire _02385_;
	wire _02386_;
	wire _02387_;
	wire _02388_;
	wire _02389_;
	wire _02390_;
	wire _02391_;
	wire _02392_;
	wire _02393_;
	wire _02394_;
	wire _02395_;
	wire _02396_;
	wire _02397_;
	wire _02398_;
	wire _02399_;
	wire _02400_;
	wire _02401_;
	wire _02402_;
	wire _02403_;
	wire _02404_;
	wire _02405_;
	wire _02406_;
	wire _02407_;
	wire _02408_;
	wire _02409_;
	wire _02410_;
	wire _02411_;
	wire _02412_;
	wire _02413_;
	wire _02414_;
	wire _02415_;
	wire _02416_;
	wire _02417_;
	wire _02418_;
	wire _02419_;
	wire _02420_;
	wire _02421_;
	wire _02422_;
	wire _02423_;
	wire _02424_;
	wire _02425_;
	wire _02426_;
	wire _02427_;
	wire _02428_;
	wire _02429_;
	wire _02430_;
	wire _02431_;
	wire _02432_;
	wire _02433_;
	wire _02434_;
	wire _02435_;
	wire _02436_;
	wire _02437_;
	wire _02438_;
	wire _02439_;
	wire _02440_;
	wire _02441_;
	wire _02442_;
	wire _02443_;
	wire _02444_;
	wire _02445_;
	wire _02446_;
	wire _02447_;
	wire _02448_;
	wire _02449_;
	wire _02450_;
	wire _02451_;
	wire _02452_;
	wire _02453_;
	wire _02454_;
	wire _02455_;
	wire _02456_;
	wire _02457_;
	wire _02458_;
	wire _02459_;
	wire _02460_;
	wire _02461_;
	wire _02462_;
	wire _02463_;
	wire _02464_;
	wire _02465_;
	wire _02466_;
	wire _02467_;
	wire _02468_;
	wire _02469_;
	wire _02470_;
	wire _02471_;
	wire _02472_;
	wire _02473_;
	wire _02474_;
	wire _02475_;
	wire _02476_;
	wire _02477_;
	wire _02478_;
	wire _02479_;
	wire _02480_;
	wire _02481_;
	wire _02482_;
	wire _02483_;
	wire _02484_;
	wire _02485_;
	wire _02486_;
	wire _02487_;
	wire _02488_;
	wire _02489_;
	wire _02490_;
	wire _02491_;
	wire _02492_;
	wire _02493_;
	wire _02494_;
	wire _02495_;
	wire _02496_;
	wire _02497_;
	wire _02498_;
	wire _02499_;
	wire _02500_;
	wire _02501_;
	wire _02502_;
	wire _02503_;
	wire _02504_;
	wire _02505_;
	wire _02506_;
	wire _02507_;
	wire _02508_;
	wire _02509_;
	wire _02510_;
	wire _02511_;
	wire _02512_;
	wire _02513_;
	wire _02514_;
	wire _02515_;
	wire _02516_;
	wire _02517_;
	wire _02518_;
	wire _02519_;
	wire _02520_;
	wire _02521_;
	wire _02522_;
	wire _02523_;
	wire _02524_;
	wire _02525_;
	wire _02526_;
	wire _02527_;
	wire _02528_;
	wire _02529_;
	wire _02530_;
	wire _02531_;
	wire _02532_;
	wire _02533_;
	wire _02534_;
	wire _02535_;
	wire _02536_;
	wire _02537_;
	wire _02538_;
	wire _02539_;
	wire _02540_;
	wire _02541_;
	wire _02542_;
	wire _02543_;
	wire _02544_;
	wire _02545_;
	wire _02546_;
	wire _02547_;
	wire _02548_;
	wire _02549_;
	wire _02550_;
	wire _02551_;
	wire _02552_;
	wire _02553_;
	wire _02554_;
	wire _02555_;
	wire _02556_;
	wire _02557_;
	wire _02558_;
	wire _02559_;
	wire _02560_;
	wire _02561_;
	wire _02562_;
	wire _02563_;
	wire _02564_;
	wire _02565_;
	wire _02566_;
	wire _02567_;
	wire _02568_;
	wire _02569_;
	wire _02570_;
	wire _02571_;
	wire _02572_;
	wire _02573_;
	wire _02574_;
	wire _02575_;
	wire _02576_;
	wire _02577_;
	wire _02578_;
	wire _02579_;
	wire _02580_;
	wire _02581_;
	wire _02582_;
	wire _02583_;
	wire _02584_;
	wire _02585_;
	wire _02586_;
	wire _02587_;
	wire _02588_;
	wire _02589_;
	wire _02590_;
	wire _02591_;
	wire _02592_;
	wire _02593_;
	wire _02594_;
	wire _02595_;
	wire _02596_;
	wire _02597_;
	wire _02598_;
	wire _02599_;
	wire _02600_;
	wire _02601_;
	wire _02602_;
	wire _02603_;
	wire _02604_;
	wire _02605_;
	wire _02606_;
	wire _02607_;
	wire _02608_;
	wire _02609_;
	wire _02610_;
	wire _02611_;
	wire _02612_;
	wire _02613_;
	wire _02614_;
	wire _02615_;
	wire _02616_;
	wire _02617_;
	wire _02618_;
	wire _02619_;
	wire _02620_;
	wire _02621_;
	wire _02622_;
	wire _02623_;
	wire _02624_;
	wire _02625_;
	wire _02626_;
	wire _02627_;
	wire _02628_;
	wire _02629_;
	wire _02630_;
	wire _02631_;
	wire _02632_;
	wire _02633_;
	wire _02634_;
	wire _02635_;
	wire _02636_;
	wire _02637_;
	wire _02638_;
	wire _02639_;
	wire _02640_;
	wire _02641_;
	wire _02642_;
	wire _02643_;
	wire _02644_;
	wire _02645_;
	wire _02646_;
	wire _02647_;
	wire _02648_;
	wire _02649_;
	wire _02650_;
	wire _02651_;
	wire _02652_;
	wire _02653_;
	wire _02654_;
	wire _02655_;
	wire _02656_;
	wire _02657_;
	wire _02658_;
	wire _02659_;
	wire _02660_;
	wire _02661_;
	wire _02662_;
	wire _02663_;
	wire _02664_;
	wire _02665_;
	wire _02666_;
	wire _02667_;
	wire _02668_;
	wire _02669_;
	wire _02670_;
	wire _02671_;
	wire _02672_;
	wire _02673_;
	wire _02674_;
	wire _02675_;
	wire _02676_;
	wire _02677_;
	wire _02678_;
	wire _02679_;
	wire _02680_;
	wire _02681_;
	wire _02682_;
	wire _02683_;
	wire _02684_;
	wire _02685_;
	wire _02686_;
	wire _02687_;
	wire _02688_;
	wire _02689_;
	wire _02690_;
	wire _02691_;
	wire _02692_;
	wire _02693_;
	wire _02694_;
	wire _02695_;
	wire _02696_;
	wire _02697_;
	wire _02698_;
	wire _02699_;
	wire _02700_;
	wire _02701_;
	wire _02702_;
	wire _02703_;
	wire _02704_;
	wire _02705_;
	wire _02706_;
	wire _02707_;
	wire _02708_;
	wire _02709_;
	wire _02710_;
	wire _02711_;
	wire _02712_;
	wire _02713_;
	wire _02714_;
	wire _02715_;
	wire _02716_;
	wire _02717_;
	wire _02718_;
	wire _02719_;
	wire _02720_;
	wire _02721_;
	wire _02722_;
	wire _02723_;
	wire _02724_;
	wire _02725_;
	wire _02726_;
	wire _02727_;
	wire _02728_;
	wire _02729_;
	wire _02730_;
	wire _02731_;
	wire _02732_;
	wire _02733_;
	wire _02734_;
	wire _02735_;
	wire _02736_;
	wire _02737_;
	wire _02738_;
	wire _02739_;
	wire _02740_;
	wire _02741_;
	wire _02742_;
	wire _02743_;
	wire _02744_;
	wire _02745_;
	wire _02746_;
	wire _02747_;
	wire _02748_;
	wire _02749_;
	wire _02750_;
	wire _02751_;
	wire _02752_;
	wire _02753_;
	wire _02754_;
	wire _02755_;
	wire _02756_;
	wire _02757_;
	wire _02758_;
	wire _02759_;
	wire _02760_;
	wire _02761_;
	wire _02762_;
	wire _02763_;
	wire _02764_;
	wire _02765_;
	wire _02766_;
	wire _02767_;
	wire _02768_;
	wire _02769_;
	wire _02770_;
	wire _02771_;
	wire _02772_;
	wire _02773_;
	wire _02774_;
	wire _02775_;
	wire _02776_;
	wire _02777_;
	wire _02778_;
	wire _02779_;
	wire _02780_;
	wire _02781_;
	wire _02782_;
	wire _02783_;
	wire _02784_;
	wire _02785_;
	wire _02786_;
	wire _02787_;
	wire _02788_;
	wire _02789_;
	wire _02790_;
	wire _02791_;
	wire _02792_;
	wire _02793_;
	wire _02794_;
	wire _02795_;
	wire _02796_;
	wire _02797_;
	wire _02798_;
	wire _02799_;
	wire _02800_;
	wire _02801_;
	wire _02802_;
	wire _02803_;
	wire _02804_;
	wire _02805_;
	wire _02806_;
	wire _02807_;
	wire _02808_;
	wire _02809_;
	wire _02810_;
	wire _02811_;
	wire _02812_;
	wire _02813_;
	wire _02814_;
	wire _02815_;
	wire _02816_;
	wire _02817_;
	wire _02818_;
	wire _02819_;
	wire _02820_;
	wire _02821_;
	wire _02822_;
	wire _02823_;
	wire _02824_;
	wire _02825_;
	wire _02826_;
	wire _02827_;
	wire _02828_;
	wire _02829_;
	wire _02830_;
	wire _02831_;
	wire _02832_;
	wire _02833_;
	wire _02834_;
	wire _02835_;
	wire _02836_;
	wire _02837_;
	wire _02838_;
	wire _02839_;
	wire _02840_;
	wire _02841_;
	wire _02842_;
	wire _02843_;
	wire _02844_;
	wire _02845_;
	wire _02846_;
	wire _02847_;
	wire _02848_;
	wire _02849_;
	wire _02850_;
	wire _02851_;
	wire _02852_;
	wire _02853_;
	wire _02854_;
	wire _02855_;
	wire _02856_;
	wire _02857_;
	wire _02858_;
	wire _02859_;
	wire _02860_;
	wire _02861_;
	wire _02862_;
	wire _02863_;
	wire _02864_;
	wire _02865_;
	wire _02866_;
	wire _02867_;
	wire _02868_;
	wire _02869_;
	wire _02870_;
	wire _02871_;
	wire _02872_;
	wire _02873_;
	wire _02874_;
	wire _02875_;
	wire _02876_;
	wire _02877_;
	wire _02878_;
	wire _02879_;
	wire _02880_;
	wire _02881_;
	wire _02882_;
	wire _02883_;
	wire _02884_;
	wire _02885_;
	wire _02886_;
	wire _02887_;
	wire _02888_;
	wire _02889_;
	wire _02890_;
	wire _02891_;
	wire _02892_;
	wire _02893_;
	wire _02894_;
	wire _02895_;
	wire _02896_;
	wire _02897_;
	wire _02898_;
	wire _02899_;
	wire _02900_;
	wire _02901_;
	wire _02902_;
	wire _02903_;
	wire _02904_;
	wire _02905_;
	wire _02906_;
	wire _02907_;
	wire _02908_;
	wire _02909_;
	wire _02910_;
	wire _02911_;
	wire _02912_;
	wire _02913_;
	wire _02914_;
	wire _02915_;
	wire _02916_;
	wire _02917_;
	wire _02918_;
	wire _02919_;
	wire _02920_;
	wire _02921_;
	wire _02922_;
	wire _02923_;
	wire _02924_;
	wire _02925_;
	wire _02926_;
	wire _02927_;
	wire _02928_;
	wire _02929_;
	wire _02930_;
	wire _02931_;
	wire _02932_;
	wire _02933_;
	wire _02934_;
	wire _02935_;
	wire _02936_;
	wire _02937_;
	wire _02938_;
	wire _02939_;
	wire _02940_;
	wire _02941_;
	wire _02942_;
	wire _02943_;
	wire _02944_;
	wire _02945_;
	wire _02946_;
	wire _02947_;
	wire _02948_;
	wire _02949_;
	wire _02950_;
	wire _02951_;
	wire _02952_;
	wire _02953_;
	wire _02954_;
	wire _02955_;
	wire _02956_;
	wire _02957_;
	wire _02958_;
	wire _02959_;
	wire _02960_;
	wire _02961_;
	wire _02962_;
	wire _02963_;
	wire _02964_;
	wire _02965_;
	wire _02966_;
	wire _02967_;
	wire _02968_;
	wire _02969_;
	wire _02970_;
	wire _02971_;
	wire _02972_;
	wire _02973_;
	wire _02974_;
	wire _02975_;
	wire _02976_;
	wire _02977_;
	wire _02978_;
	wire _02979_;
	wire _02980_;
	wire _02981_;
	wire _02982_;
	wire _02983_;
	wire _02984_;
	wire _02985_;
	wire _02986_;
	wire _02987_;
	wire _02988_;
	wire _02989_;
	wire _02990_;
	wire _02991_;
	wire _02992_;
	wire _02993_;
	wire _02994_;
	wire _02995_;
	wire _02996_;
	wire _02997_;
	wire _02998_;
	wire _02999_;
	wire _03000_;
	wire _03001_;
	wire _03002_;
	wire _03003_;
	wire _03004_;
	wire _03005_;
	wire _03006_;
	wire _03007_;
	wire _03008_;
	wire _03009_;
	wire _03010_;
	wire _03011_;
	wire _03012_;
	wire _03013_;
	wire _03014_;
	wire _03015_;
	wire _03016_;
	wire _03017_;
	wire _03018_;
	wire _03019_;
	wire _03020_;
	wire _03021_;
	wire _03022_;
	wire _03023_;
	wire _03024_;
	wire _03025_;
	wire _03026_;
	wire _03027_;
	wire _03028_;
	wire _03029_;
	wire _03030_;
	wire _03031_;
	wire _03032_;
	wire _03033_;
	wire _03034_;
	wire _03035_;
	wire _03036_;
	wire _03037_;
	wire _03038_;
	wire _03039_;
	wire _03040_;
	wire _03041_;
	wire _03042_;
	wire _03043_;
	wire _03044_;
	wire _03045_;
	wire _03046_;
	wire _03047_;
	wire _03048_;
	wire _03049_;
	wire _03050_;
	wire _03051_;
	wire _03052_;
	wire _03053_;
	wire _03054_;
	wire _03055_;
	wire _03056_;
	wire _03057_;
	wire _03058_;
	wire _03059_;
	wire _03060_;
	wire _03061_;
	wire _03062_;
	wire _03063_;
	wire _03064_;
	wire _03065_;
	wire _03066_;
	wire _03067_;
	wire _03068_;
	wire _03069_;
	wire _03070_;
	wire _03071_;
	wire _03072_;
	wire _03073_;
	wire _03074_;
	wire _03075_;
	wire _03076_;
	wire _03077_;
	wire _03078_;
	wire _03079_;
	wire _03080_;
	wire _03081_;
	wire _03082_;
	wire _03083_;
	wire _03084_;
	wire _03085_;
	wire _03086_;
	wire _03087_;
	wire _03088_;
	wire _03089_;
	wire _03090_;
	wire _03091_;
	wire _03092_;
	wire _03093_;
	wire _03094_;
	wire _03095_;
	wire _03096_;
	wire _03097_;
	wire _03098_;
	wire _03099_;
	wire _03100_;
	wire _03101_;
	wire _03102_;
	wire _03103_;
	wire _03104_;
	wire _03105_;
	wire _03106_;
	wire _03107_;
	wire _03108_;
	wire _03109_;
	wire _03110_;
	wire _03111_;
	wire _03112_;
	wire _03113_;
	wire _03114_;
	wire _03115_;
	wire _03116_;
	wire _03117_;
	wire _03118_;
	wire _03119_;
	wire _03120_;
	wire _03121_;
	wire _03122_;
	wire _03123_;
	wire _03124_;
	wire _03125_;
	wire _03126_;
	wire _03127_;
	wire _03128_;
	wire _03129_;
	wire _03130_;
	wire _03131_;
	wire _03132_;
	wire _03133_;
	wire _03134_;
	wire _03135_;
	wire _03136_;
	wire _03137_;
	wire _03138_;
	wire _03139_;
	wire _03140_;
	wire _03141_;
	wire _03142_;
	wire _03143_;
	wire _03144_;
	wire _03145_;
	wire _03146_;
	wire _03147_;
	wire _03148_;
	wire _03149_;
	wire _03150_;
	wire _03151_;
	wire _03152_;
	wire _03153_;
	wire _03154_;
	wire _03155_;
	wire _03156_;
	wire _03157_;
	wire _03158_;
	wire _03159_;
	wire _03160_;
	wire _03161_;
	wire _03162_;
	wire _03163_;
	wire _03164_;
	wire _03165_;
	wire _03166_;
	wire _03167_;
	wire _03168_;
	wire _03169_;
	wire _03170_;
	wire _03171_;
	wire _03172_;
	wire _03173_;
	wire _03174_;
	wire _03175_;
	wire _03176_;
	wire _03177_;
	wire _03178_;
	wire _03179_;
	wire _03180_;
	wire _03181_;
	wire _03182_;
	wire _03183_;
	wire _03184_;
	wire _03185_;
	wire _03186_;
	wire _03187_;
	wire _03188_;
	wire _03189_;
	wire _03190_;
	wire _03191_;
	wire _03192_;
	wire _03193_;
	wire _03194_;
	wire _03195_;
	wire _03196_;
	wire _03197_;
	wire _03198_;
	wire _03199_;
	wire _03200_;
	wire _03201_;
	wire _03202_;
	wire _03203_;
	wire _03204_;
	wire _03205_;
	wire _03206_;
	wire _03207_;
	wire _03208_;
	wire _03209_;
	wire _03210_;
	wire _03211_;
	wire _03212_;
	wire _03213_;
	wire _03214_;
	wire _03215_;
	wire _03216_;
	wire _03217_;
	wire _03218_;
	wire _03219_;
	wire _03220_;
	wire _03221_;
	wire _03222_;
	wire _03223_;
	wire _03224_;
	wire _03225_;
	wire _03226_;
	wire _03227_;
	wire _03228_;
	wire _03229_;
	wire _03230_;
	wire _03231_;
	wire _03232_;
	wire _03233_;
	wire _03234_;
	wire _03235_;
	wire _03236_;
	wire _03237_;
	wire _03238_;
	wire _03239_;
	wire _03240_;
	wire _03241_;
	wire _03242_;
	wire _03243_;
	wire _03244_;
	wire _03245_;
	wire _03246_;
	wire _03247_;
	wire _03248_;
	wire _03249_;
	wire _03250_;
	wire _03251_;
	wire _03252_;
	wire _03253_;
	wire _03254_;
	wire _03255_;
	wire _03256_;
	wire _03257_;
	wire _03258_;
	wire _03259_;
	wire _03260_;
	wire _03261_;
	wire _03262_;
	wire _03263_;
	wire _03264_;
	wire _03265_;
	wire _03266_;
	wire _03267_;
	wire _03268_;
	wire _03269_;
	wire _03270_;
	wire _03271_;
	wire _03272_;
	wire _03273_;
	wire _03274_;
	wire _03275_;
	wire _03276_;
	wire _03277_;
	wire _03278_;
	wire _03279_;
	wire _03280_;
	wire _03281_;
	wire _03282_;
	wire _03283_;
	wire _03284_;
	wire _03285_;
	wire _03286_;
	wire _03287_;
	wire _03288_;
	wire _03289_;
	wire _03290_;
	wire _03291_;
	wire _03292_;
	wire _03293_;
	wire _03294_;
	wire _03295_;
	wire _03296_;
	wire _03297_;
	wire _03298_;
	wire _03299_;
	wire _03300_;
	wire _03301_;
	wire _03302_;
	wire _03303_;
	wire _03304_;
	wire _03305_;
	wire _03306_;
	wire _03307_;
	wire _03308_;
	wire _03309_;
	wire _03310_;
	wire _03311_;
	wire _03312_;
	wire _03313_;
	wire _03314_;
	wire _03315_;
	wire _03316_;
	wire _03317_;
	wire _03318_;
	wire _03319_;
	wire _03320_;
	wire _03321_;
	wire _03322_;
	wire _03323_;
	wire _03324_;
	wire _03325_;
	wire _03326_;
	wire _03327_;
	wire _03328_;
	wire _03329_;
	wire _03330_;
	wire _03331_;
	wire _03332_;
	wire _03333_;
	wire _03334_;
	wire _03335_;
	wire _03336_;
	wire _03337_;
	wire _03338_;
	wire _03339_;
	wire _03340_;
	wire _03341_;
	wire _03342_;
	wire _03343_;
	wire _03344_;
	wire _03345_;
	wire _03346_;
	wire _03347_;
	wire _03348_;
	wire _03349_;
	wire _03350_;
	wire _03351_;
	wire _03352_;
	wire _03353_;
	wire _03354_;
	wire _03355_;
	wire _03356_;
	wire _03357_;
	wire _03358_;
	wire _03359_;
	wire _03360_;
	wire _03361_;
	wire _03362_;
	wire _03363_;
	wire _03364_;
	wire _03365_;
	wire _03366_;
	wire _03367_;
	wire _03368_;
	wire _03369_;
	wire _03370_;
	wire _03371_;
	wire _03372_;
	wire _03373_;
	wire _03374_;
	wire _03375_;
	wire _03376_;
	wire _03377_;
	wire _03378_;
	wire _03379_;
	wire _03380_;
	wire _03381_;
	wire _03382_;
	wire _03383_;
	wire _03384_;
	wire _03385_;
	wire _03386_;
	wire _03387_;
	wire _03388_;
	wire _03389_;
	wire _03390_;
	wire _03391_;
	wire _03392_;
	wire _03393_;
	wire _03394_;
	wire _03395_;
	wire _03396_;
	wire _03397_;
	wire _03398_;
	wire _03399_;
	wire _03400_;
	wire _03401_;
	wire _03402_;
	wire _03403_;
	wire _03404_;
	wire _03405_;
	wire _03406_;
	wire _03407_;
	wire _03408_;
	wire _03409_;
	wire _03410_;
	wire _03411_;
	wire _03412_;
	wire _03413_;
	wire _03414_;
	wire _03415_;
	wire _03416_;
	wire _03417_;
	wire _03418_;
	wire _03419_;
	wire _03420_;
	wire _03421_;
	wire _03422_;
	wire _03423_;
	wire _03424_;
	wire _03425_;
	wire _03426_;
	wire _03427_;
	wire _03428_;
	wire _03429_;
	wire _03430_;
	wire _03431_;
	wire _03432_;
	wire _03433_;
	wire _03434_;
	wire _03435_;
	wire _03436_;
	wire _03437_;
	wire _03438_;
	wire _03439_;
	wire _03440_;
	wire _03441_;
	wire _03442_;
	wire _03443_;
	wire _03444_;
	wire _03445_;
	wire _03446_;
	wire _03447_;
	wire _03448_;
	wire _03449_;
	wire _03450_;
	wire _03451_;
	wire _03452_;
	wire _03453_;
	wire _03454_;
	wire _03455_;
	wire _03456_;
	wire _03457_;
	wire _03458_;
	wire _03459_;
	wire _03460_;
	wire _03461_;
	wire _03462_;
	wire _03463_;
	wire _03464_;
	wire _03465_;
	wire _03466_;
	wire _03467_;
	wire _03468_;
	wire _03469_;
	wire _03470_;
	wire _03471_;
	wire _03472_;
	wire _03473_;
	wire _03474_;
	wire _03475_;
	wire _03476_;
	wire _03477_;
	wire _03478_;
	wire _03479_;
	wire _03480_;
	wire _03481_;
	wire _03482_;
	wire _03483_;
	wire _03484_;
	wire _03485_;
	wire _03486_;
	wire _03487_;
	wire _03488_;
	wire _03489_;
	wire _03490_;
	wire _03491_;
	wire _03492_;
	wire _03493_;
	wire _03494_;
	wire _03495_;
	wire _03496_;
	wire _03497_;
	wire _03498_;
	wire _03499_;
	wire _03500_;
	wire _03501_;
	wire _03502_;
	wire _03503_;
	wire _03504_;
	wire _03505_;
	wire _03506_;
	wire _03507_;
	wire _03508_;
	wire _03509_;
	wire _03510_;
	wire _03511_;
	wire _03512_;
	wire _03513_;
	wire _03514_;
	wire _03515_;
	wire _03516_;
	wire _03517_;
	wire _03518_;
	wire _03519_;
	wire _03520_;
	wire _03521_;
	wire _03522_;
	wire _03523_;
	wire _03524_;
	wire _03525_;
	wire _03526_;
	wire _03527_;
	wire _03528_;
	wire _03529_;
	wire _03530_;
	wire _03531_;
	wire _03532_;
	wire _03533_;
	wire _03534_;
	wire _03535_;
	wire _03536_;
	wire _03537_;
	wire _03538_;
	wire _03539_;
	wire _03540_;
	wire _03541_;
	wire _03542_;
	wire _03543_;
	wire _03544_;
	wire _03545_;
	wire _03546_;
	wire _03547_;
	wire _03548_;
	wire _03549_;
	wire _03550_;
	wire _03551_;
	wire _03552_;
	wire _03553_;
	wire _03554_;
	wire _03555_;
	wire _03556_;
	wire _03557_;
	wire _03558_;
	wire _03559_;
	wire _03560_;
	wire _03561_;
	wire _03562_;
	wire _03563_;
	wire _03564_;
	wire _03565_;
	wire _03566_;
	wire _03567_;
	wire _03568_;
	wire _03569_;
	wire _03570_;
	wire _03571_;
	wire _03572_;
	wire _03573_;
	wire _03574_;
	wire _03575_;
	wire _03576_;
	wire _03577_;
	wire _03578_;
	wire _03579_;
	wire _03580_;
	wire _03581_;
	wire _03582_;
	wire _03583_;
	wire _03584_;
	wire _03585_;
	wire _03586_;
	wire _03587_;
	wire _03588_;
	wire _03589_;
	wire _03590_;
	wire _03591_;
	wire _03592_;
	wire _03593_;
	wire _03594_;
	wire _03595_;
	wire _03596_;
	wire _03597_;
	wire _03598_;
	wire _03599_;
	wire _03600_;
	wire _03601_;
	wire _03602_;
	wire _03603_;
	wire _03604_;
	wire _03605_;
	wire _03606_;
	wire _03607_;
	wire _03608_;
	wire _03609_;
	wire _03610_;
	wire _03611_;
	wire _03612_;
	wire _03613_;
	wire _03614_;
	wire _03615_;
	wire _03616_;
	wire _03617_;
	wire _03618_;
	wire _03619_;
	wire _03620_;
	wire _03621_;
	wire _03622_;
	wire _03623_;
	wire _03624_;
	wire _03625_;
	wire _03626_;
	wire _03627_;
	wire _03628_;
	wire _03629_;
	wire _03630_;
	wire _03631_;
	wire _03632_;
	wire _03633_;
	wire _03634_;
	wire _03635_;
	wire _03636_;
	wire _03637_;
	wire _03638_;
	wire _03639_;
	wire _03640_;
	wire _03641_;
	wire _03642_;
	wire _03643_;
	wire _03644_;
	wire _03645_;
	wire _03646_;
	wire _03647_;
	wire _03648_;
	wire _03649_;
	wire _03650_;
	wire _03651_;
	wire _03652_;
	wire _03653_;
	wire _03654_;
	wire _03655_;
	wire _03656_;
	wire _03657_;
	wire _03658_;
	wire _03659_;
	wire _03660_;
	wire _03661_;
	wire _03662_;
	wire _03663_;
	wire _03664_;
	wire _03665_;
	wire _03666_;
	wire _03667_;
	wire _03668_;
	wire _03669_;
	wire _03670_;
	wire _03671_;
	wire _03672_;
	wire _03673_;
	wire _03674_;
	wire _03675_;
	wire _03676_;
	wire _03677_;
	wire _03678_;
	wire _03679_;
	wire _03680_;
	wire _03681_;
	wire _03682_;
	wire _03683_;
	wire _03684_;
	wire _03685_;
	wire _03686_;
	wire _03687_;
	wire _03688_;
	wire _03689_;
	wire _03690_;
	wire _03691_;
	wire _03692_;
	wire _03693_;
	wire _03694_;
	wire _03695_;
	wire _03696_;
	wire _03697_;
	wire _03698_;
	wire _03699_;
	wire _03700_;
	wire _03701_;
	wire _03702_;
	wire _03703_;
	wire _03704_;
	wire _03705_;
	wire _03706_;
	wire _03707_;
	wire _03708_;
	wire _03709_;
	wire _03710_;
	wire _03711_;
	wire _03712_;
	wire _03713_;
	wire _03714_;
	wire _03715_;
	wire _03716_;
	wire _03717_;
	wire _03718_;
	wire _03719_;
	wire _03720_;
	wire _03721_;
	wire _03722_;
	wire _03723_;
	wire _03724_;
	wire _03725_;
	wire _03726_;
	wire _03727_;
	wire _03728_;
	wire _03729_;
	wire _03730_;
	wire _03731_;
	wire _03732_;
	wire _03733_;
	wire _03734_;
	wire _03735_;
	wire _03736_;
	wire _03737_;
	wire _03738_;
	wire _03739_;
	wire _03740_;
	wire _03741_;
	wire _03742_;
	wire _03743_;
	wire _03744_;
	wire _03745_;
	wire _03746_;
	wire _03747_;
	wire _03748_;
	wire _03749_;
	wire _03750_;
	wire _03751_;
	wire _03752_;
	wire _03753_;
	wire _03754_;
	wire _03755_;
	wire _03756_;
	wire _03757_;
	wire _03758_;
	wire _03759_;
	wire _03760_;
	wire _03761_;
	wire _03762_;
	wire _03763_;
	wire _03764_;
	wire _03765_;
	wire _03766_;
	wire _03767_;
	wire _03768_;
	wire _03769_;
	wire _03770_;
	wire _03771_;
	wire _03772_;
	wire _03773_;
	wire _03774_;
	wire _03775_;
	wire _03776_;
	wire _03777_;
	wire _03778_;
	wire _03779_;
	wire _03780_;
	wire _03781_;
	wire _03782_;
	wire _03783_;
	wire _03784_;
	wire _03785_;
	wire _03786_;
	wire _03787_;
	wire _03788_;
	wire _03789_;
	wire _03790_;
	wire _03791_;
	wire _03792_;
	wire _03793_;
	wire _03794_;
	wire _03795_;
	wire _03796_;
	wire _03797_;
	wire _03798_;
	wire _03799_;
	wire _03800_;
	wire _03801_;
	wire _03802_;
	wire _03803_;
	wire _03804_;
	wire _03805_;
	wire _03806_;
	wire _03807_;
	wire _03808_;
	wire _03809_;
	wire _03810_;
	wire _03811_;
	wire _03812_;
	wire _03813_;
	wire _03814_;
	wire _03815_;
	wire _03816_;
	wire _03817_;
	wire _03818_;
	wire _03819_;
	wire _03820_;
	wire _03821_;
	wire _03822_;
	wire _03823_;
	wire _03824_;
	wire _03825_;
	wire _03826_;
	wire _03827_;
	wire _03828_;
	wire _03829_;
	wire _03830_;
	wire _03831_;
	wire _03832_;
	wire _03833_;
	wire _03834_;
	wire _03835_;
	wire _03836_;
	wire _03837_;
	wire _03838_;
	wire _03839_;
	wire _03840_;
	wire _03841_;
	wire _03842_;
	wire _03843_;
	wire _03844_;
	wire _03845_;
	wire _03846_;
	wire _03847_;
	wire _03848_;
	wire _03849_;
	wire _03850_;
	wire _03851_;
	wire _03852_;
	wire _03853_;
	wire _03854_;
	wire _03855_;
	wire _03856_;
	wire _03857_;
	wire _03858_;
	wire _03859_;
	wire _03860_;
	wire _03861_;
	wire _03862_;
	wire _03863_;
	wire _03864_;
	wire _03865_;
	wire _03866_;
	wire _03867_;
	wire _03868_;
	wire _03869_;
	wire _03870_;
	wire _03871_;
	wire _03872_;
	wire _03873_;
	wire _03874_;
	wire _03875_;
	wire _03876_;
	wire _03877_;
	wire _03878_;
	wire _03879_;
	wire _03880_;
	wire _03881_;
	wire _03882_;
	wire _03883_;
	wire _03884_;
	wire _03885_;
	wire _03886_;
	wire _03887_;
	wire _03888_;
	wire _03889_;
	wire _03890_;
	wire _03891_;
	wire _03892_;
	wire _03893_;
	wire _03894_;
	wire _03895_;
	wire _03896_;
	wire _03897_;
	wire _03898_;
	wire _03899_;
	wire _03900_;
	wire _03901_;
	wire _03902_;
	wire _03903_;
	wire _03904_;
	wire _03905_;
	wire _03906_;
	wire _03907_;
	wire _03908_;
	wire _03909_;
	wire _03910_;
	wire _03911_;
	wire _03912_;
	wire _03913_;
	wire _03914_;
	wire _03915_;
	wire _03916_;
	wire _03917_;
	wire _03918_;
	wire _03919_;
	wire _03920_;
	wire _03921_;
	wire _03922_;
	wire _03923_;
	wire _03924_;
	wire _03925_;
	wire _03926_;
	wire _03927_;
	wire _03928_;
	wire _03929_;
	wire _03930_;
	wire _03931_;
	wire _03932_;
	wire _03933_;
	wire _03934_;
	wire _03935_;
	wire _03936_;
	wire _03937_;
	wire _03938_;
	wire _03939_;
	wire _03940_;
	wire _03941_;
	wire _03942_;
	wire _03943_;
	wire _03944_;
	wire _03945_;
	wire _03946_;
	wire _03947_;
	wire _03948_;
	wire _03949_;
	wire _03950_;
	wire _03951_;
	wire _03952_;
	wire _03953_;
	wire _03954_;
	wire _03955_;
	wire _03956_;
	wire _03957_;
	wire _03958_;
	wire _03959_;
	wire _03960_;
	wire _03961_;
	wire _03962_;
	wire _03963_;
	wire _03964_;
	wire _03965_;
	wire _03966_;
	wire _03967_;
	wire _03968_;
	wire _03969_;
	wire _03970_;
	wire _03971_;
	wire _03972_;
	wire _03973_;
	wire _03974_;
	wire _03975_;
	wire _03976_;
	wire _03977_;
	wire _03978_;
	wire _03979_;
	wire _03980_;
	wire _03981_;
	wire _03982_;
	wire _03983_;
	wire _03984_;
	wire _03985_;
	wire _03986_;
	wire _03987_;
	wire _03988_;
	wire _03989_;
	wire _03990_;
	wire _03991_;
	wire _03992_;
	wire _03993_;
	wire _03994_;
	wire _03995_;
	wire _03996_;
	wire _03997_;
	wire _03998_;
	wire _03999_;
	wire _04000_;
	wire _04001_;
	wire _04002_;
	wire _04003_;
	wire _04004_;
	wire _04005_;
	wire _04006_;
	wire _04007_;
	wire _04008_;
	wire _04009_;
	wire _04010_;
	wire _04011_;
	wire _04012_;
	wire _04013_;
	wire _04014_;
	wire _04015_;
	wire _04016_;
	wire _04017_;
	wire _04018_;
	wire _04019_;
	wire _04020_;
	wire _04021_;
	wire _04022_;
	wire _04023_;
	wire _04024_;
	wire _04025_;
	wire _04026_;
	wire _04027_;
	wire _04028_;
	wire _04029_;
	wire _04030_;
	wire _04031_;
	wire _04032_;
	wire _04033_;
	wire _04034_;
	wire _04035_;
	wire _04036_;
	wire _04037_;
	wire _04038_;
	wire _04039_;
	wire _04040_;
	wire _04041_;
	wire _04042_;
	wire _04043_;
	wire _04044_;
	wire _04045_;
	wire _04046_;
	wire _04047_;
	wire _04048_;
	wire _04049_;
	wire _04050_;
	wire _04051_;
	wire _04052_;
	wire _04053_;
	wire _04054_;
	wire _04055_;
	wire _04056_;
	wire _04057_;
	wire _04058_;
	wire _04059_;
	wire _04060_;
	wire _04061_;
	wire _04062_;
	wire _04063_;
	wire _04064_;
	wire _04065_;
	wire _04066_;
	wire _04067_;
	wire _04068_;
	wire _04069_;
	wire _04070_;
	wire _04071_;
	wire _04072_;
	wire _04073_;
	wire _04074_;
	wire _04075_;
	wire _04076_;
	wire _04077_;
	wire _04078_;
	wire _04079_;
	wire _04080_;
	wire _04081_;
	wire _04082_;
	wire _04083_;
	wire _04084_;
	wire _04085_;
	wire _04086_;
	wire _04087_;
	wire _04088_;
	wire _04089_;
	wire _04090_;
	wire _04091_;
	wire _04092_;
	wire _04093_;
	wire _04094_;
	wire _04095_;
	wire _04096_;
	wire _04097_;
	wire _04098_;
	wire _04099_;
	wire _04100_;
	wire _04101_;
	wire _04102_;
	wire _04103_;
	wire _04104_;
	wire _04105_;
	wire _04106_;
	wire _04107_;
	wire _04108_;
	wire _04109_;
	wire _04110_;
	wire _04111_;
	wire _04112_;
	wire _04113_;
	wire _04114_;
	wire _04115_;
	wire _04116_;
	wire _04117_;
	wire _04118_;
	wire _04119_;
	wire _04120_;
	wire _04121_;
	wire _04122_;
	wire _04123_;
	wire _04124_;
	wire _04125_;
	wire _04126_;
	wire _04127_;
	wire _04128_;
	wire _04129_;
	wire _04130_;
	wire _04131_;
	wire _04132_;
	wire _04133_;
	wire _04134_;
	wire _04135_;
	wire _04136_;
	wire _04137_;
	wire _04138_;
	wire _04139_;
	wire _04140_;
	wire _04141_;
	wire _04142_;
	wire _04143_;
	wire _04144_;
	wire _04145_;
	wire _04146_;
	wire _04147_;
	wire _04148_;
	wire _04149_;
	wire _04150_;
	wire _04151_;
	wire _04152_;
	wire _04153_;
	wire _04154_;
	wire _04155_;
	wire _04156_;
	wire _04157_;
	wire _04158_;
	wire _04159_;
	wire _04160_;
	wire _04161_;
	wire _04162_;
	wire _04163_;
	wire _04164_;
	wire _04165_;
	wire _04166_;
	wire _04167_;
	wire _04168_;
	wire _04169_;
	wire _04170_;
	wire _04171_;
	wire _04172_;
	wire _04173_;
	wire _04174_;
	wire _04175_;
	wire _04176_;
	wire _04177_;
	wire _04178_;
	wire _04179_;
	wire _04180_;
	wire _04181_;
	wire _04182_;
	wire _04183_;
	wire _04184_;
	wire _04185_;
	wire _04186_;
	wire _04187_;
	wire _04188_;
	wire _04189_;
	wire _04190_;
	wire _04191_;
	wire _04192_;
	wire _04193_;
	wire _04194_;
	wire _04195_;
	wire _04196_;
	wire _04197_;
	wire _04198_;
	wire _04199_;
	wire _04200_;
	wire _04201_;
	wire _04202_;
	wire _04203_;
	wire _04204_;
	wire _04205_;
	wire _04206_;
	wire _04207_;
	wire _04208_;
	wire _04209_;
	wire _04210_;
	wire _04211_;
	wire _04212_;
	wire _04213_;
	wire _04214_;
	wire _04215_;
	wire _04216_;
	wire _04217_;
	wire _04218_;
	wire _04219_;
	wire _04220_;
	wire _04221_;
	wire _04222_;
	wire _04223_;
	wire _04224_;
	wire _04225_;
	wire _04226_;
	wire _04227_;
	wire _04228_;
	wire _04229_;
	wire _04230_;
	wire _04231_;
	wire _04232_;
	wire _04233_;
	wire _04234_;
	wire _04235_;
	wire _04236_;
	wire _04237_;
	wire _04238_;
	wire _04239_;
	wire _04240_;
	wire _04241_;
	wire _04242_;
	wire _04243_;
	wire _04244_;
	wire _04245_;
	wire _04246_;
	wire _04247_;
	wire _04248_;
	wire _04249_;
	wire _04250_;
	wire _04251_;
	wire _04252_;
	wire _04253_;
	wire _04254_;
	wire _04255_;
	wire _04256_;
	wire _04257_;
	wire _04258_;
	wire _04259_;
	wire _04260_;
	wire _04261_;
	wire _04262_;
	wire _04263_;
	wire _04264_;
	wire _04265_;
	wire _04266_;
	wire _04267_;
	wire _04268_;
	wire _04269_;
	wire _04270_;
	wire _04271_;
	wire _04272_;
	wire _04273_;
	wire _04274_;
	wire _04275_;
	wire _04276_;
	wire _04277_;
	wire _04278_;
	wire _04279_;
	wire _04280_;
	wire _04281_;
	wire _04282_;
	wire _04283_;
	wire _04284_;
	wire _04285_;
	wire _04286_;
	wire _04287_;
	wire _04288_;
	wire _04289_;
	wire _04290_;
	wire _04291_;
	wire _04292_;
	wire _04293_;
	wire _04294_;
	wire _04295_;
	wire _04296_;
	wire _04297_;
	wire _04298_;
	wire _04299_;
	wire _04300_;
	wire _04301_;
	wire _04302_;
	wire _04303_;
	wire _04304_;
	wire _04305_;
	wire _04306_;
	wire _04307_;
	wire _04308_;
	wire _04309_;
	wire _04310_;
	wire _04311_;
	wire _04312_;
	wire _04313_;
	wire _04314_;
	wire _04315_;
	wire _04316_;
	wire _04317_;
	wire _04318_;
	wire _04319_;
	wire _04320_;
	wire _04321_;
	wire _04322_;
	wire _04323_;
	wire _04324_;
	wire _04325_;
	wire _04326_;
	wire _04327_;
	wire _04328_;
	wire _04329_;
	wire _04330_;
	wire _04331_;
	wire _04332_;
	wire _04333_;
	wire _04334_;
	wire _04335_;
	wire _04336_;
	wire _04337_;
	wire _04338_;
	wire _04339_;
	wire _04340_;
	wire _04341_;
	wire _04342_;
	wire _04343_;
	wire _04344_;
	wire _04345_;
	wire _04346_;
	wire _04347_;
	wire _04348_;
	wire _04349_;
	wire _04350_;
	wire _04351_;
	wire _04352_;
	wire _04353_;
	wire _04354_;
	wire _04355_;
	wire _04356_;
	wire _04357_;
	wire _04358_;
	wire _04359_;
	wire _04360_;
	wire _04361_;
	wire _04362_;
	wire _04363_;
	wire _04364_;
	wire _04365_;
	wire _04366_;
	wire _04367_;
	wire _04368_;
	wire _04369_;
	wire _04370_;
	wire _04371_;
	wire _04372_;
	wire _04373_;
	wire _04374_;
	wire _04375_;
	wire _04376_;
	wire _04377_;
	wire _04378_;
	wire _04379_;
	wire _04380_;
	wire _04381_;
	wire _04382_;
	wire _04383_;
	wire _04384_;
	wire _04385_;
	wire _04386_;
	wire _04387_;
	wire _04388_;
	wire _04389_;
	wire _04390_;
	wire _04391_;
	wire _04392_;
	wire _04393_;
	wire _04394_;
	wire _04395_;
	wire _04396_;
	wire _04397_;
	wire _04398_;
	wire _04399_;
	wire _04400_;
	wire _04401_;
	wire _04402_;
	wire _04403_;
	wire _04404_;
	wire _04405_;
	wire _04406_;
	wire _04407_;
	wire _04408_;
	wire _04409_;
	wire _04410_;
	wire _04411_;
	wire _04412_;
	wire _04413_;
	wire _04414_;
	wire _04415_;
	wire _04416_;
	wire _04417_;
	wire _04418_;
	wire _04419_;
	wire _04420_;
	wire _04421_;
	wire _04422_;
	wire _04423_;
	wire _04424_;
	wire _04425_;
	wire _04426_;
	wire _04427_;
	wire _04428_;
	wire _04429_;
	wire _04430_;
	wire _04431_;
	wire _04432_;
	wire _04433_;
	wire _04434_;
	wire _04435_;
	wire _04436_;
	wire _04437_;
	wire _04438_;
	wire _04439_;
	wire _04440_;
	wire _04441_;
	wire _04442_;
	wire _04443_;
	wire _04444_;
	wire _04445_;
	wire _04446_;
	wire _04447_;
	wire _04448_;
	wire _04449_;
	wire _04450_;
	wire _04451_;
	wire _04452_;
	wire _04453_;
	wire _04454_;
	wire _04455_;
	wire _04456_;
	wire _04457_;
	wire _04458_;
	wire _04459_;
	wire _04460_;
	wire _04461_;
	wire _04462_;
	wire _04463_;
	wire _04464_;
	wire _04465_;
	wire _04466_;
	wire _04467_;
	wire _04468_;
	wire _04469_;
	wire _04470_;
	wire _04471_;
	wire _04472_;
	wire _04473_;
	wire _04474_;
	wire _04475_;
	wire _04476_;
	wire _04477_;
	wire _04478_;
	wire _04479_;
	wire _04480_;
	wire _04481_;
	wire _04482_;
	wire _04483_;
	wire _04484_;
	wire _04485_;
	wire _04486_;
	wire _04487_;
	wire _04488_;
	wire _04489_;
	wire _04490_;
	wire _04491_;
	wire _04492_;
	wire _04493_;
	wire _04494_;
	wire _04495_;
	wire _04496_;
	wire _04497_;
	wire _04498_;
	wire _04499_;
	wire _04500_;
	wire _04501_;
	wire _04502_;
	wire _04503_;
	wire _04504_;
	wire _04505_;
	wire _04506_;
	wire _04507_;
	wire _04508_;
	wire _04509_;
	wire _04510_;
	wire _04511_;
	wire _04512_;
	wire _04513_;
	wire _04514_;
	wire _04515_;
	wire _04516_;
	wire _04517_;
	wire _04518_;
	wire _04519_;
	wire _04520_;
	wire _04521_;
	wire _04522_;
	wire _04523_;
	wire _04524_;
	wire _04525_;
	wire _04526_;
	wire _04527_;
	wire _04528_;
	wire _04529_;
	wire _04530_;
	wire _04531_;
	wire _04532_;
	wire _04533_;
	wire _04534_;
	wire _04535_;
	wire _04536_;
	wire _04537_;
	wire _04538_;
	wire _04539_;
	wire _04540_;
	wire _04541_;
	wire _04542_;
	wire _04543_;
	wire _04544_;
	wire _04545_;
	wire _04546_;
	wire _04547_;
	wire _04548_;
	wire _04549_;
	wire _04550_;
	wire _04551_;
	wire _04552_;
	wire _04553_;
	wire _04554_;
	wire _04555_;
	wire _04556_;
	wire _04557_;
	wire _04558_;
	wire _04559_;
	wire _04560_;
	wire _04561_;
	wire _04562_;
	wire _04563_;
	wire _04564_;
	wire _04565_;
	wire _04566_;
	wire _04567_;
	wire _04568_;
	wire _04569_;
	wire _04570_;
	wire _04571_;
	wire _04572_;
	wire _04573_;
	wire _04574_;
	wire _04575_;
	wire _04576_;
	wire _04577_;
	wire _04578_;
	wire _04579_;
	wire _04580_;
	wire _04581_;
	wire _04582_;
	wire _04583_;
	wire _04584_;
	wire _04585_;
	wire _04586_;
	wire _04587_;
	wire _04588_;
	wire _04589_;
	wire _04590_;
	wire _04591_;
	wire _04592_;
	wire _04593_;
	wire _04594_;
	wire _04595_;
	wire _04596_;
	wire _04597_;
	wire _04598_;
	wire _04599_;
	wire _04600_;
	wire _04601_;
	wire _04602_;
	wire _04603_;
	wire _04604_;
	wire _04605_;
	wire _04606_;
	wire _04607_;
	wire _04608_;
	wire _04609_;
	wire _04610_;
	wire _04611_;
	wire _04612_;
	wire _04613_;
	wire _04614_;
	wire _04615_;
	wire _04616_;
	wire _04617_;
	wire _04618_;
	wire _04619_;
	wire _04620_;
	wire _04621_;
	wire _04622_;
	wire _04623_;
	wire _04624_;
	wire _04625_;
	wire _04626_;
	wire _04627_;
	wire _04628_;
	wire _04629_;
	wire _04630_;
	wire _04631_;
	wire _04632_;
	wire _04633_;
	wire _04634_;
	wire _04635_;
	wire _04636_;
	wire _04637_;
	wire _04638_;
	wire _04639_;
	wire _04640_;
	wire _04641_;
	wire _04642_;
	wire _04643_;
	wire _04644_;
	wire _04645_;
	wire _04646_;
	wire _04647_;
	wire _04648_;
	wire _04649_;
	wire _04650_;
	wire _04651_;
	wire _04652_;
	wire _04653_;
	wire _04654_;
	wire _04655_;
	wire _04656_;
	wire _04657_;
	wire _04658_;
	wire _04659_;
	wire _04660_;
	wire _04661_;
	wire _04662_;
	wire _04663_;
	wire _04664_;
	wire _04665_;
	wire _04666_;
	wire _04667_;
	wire _04668_;
	wire _04669_;
	wire _04670_;
	wire _04671_;
	wire _04672_;
	wire _04673_;
	wire _04674_;
	wire _04675_;
	wire _04676_;
	wire _04677_;
	wire _04678_;
	wire _04679_;
	wire _04680_;
	wire _04681_;
	wire _04682_;
	wire _04683_;
	wire _04684_;
	wire _04685_;
	wire _04686_;
	wire _04687_;
	wire _04688_;
	wire _04689_;
	wire _04690_;
	wire _04691_;
	wire _04692_;
	wire _04693_;
	wire _04694_;
	wire _04695_;
	wire _04696_;
	wire _04697_;
	wire _04698_;
	wire _04699_;
	wire _04700_;
	wire _04701_;
	wire _04702_;
	wire _04703_;
	wire _04704_;
	wire _04705_;
	wire _04706_;
	wire _04707_;
	wire _04708_;
	wire _04709_;
	wire _04710_;
	wire _04711_;
	wire _04712_;
	wire _04713_;
	wire _04714_;
	wire _04715_;
	wire _04716_;
	wire _04717_;
	wire _04718_;
	wire _04719_;
	wire _04720_;
	wire _04721_;
	wire _04722_;
	wire _04723_;
	wire _04724_;
	wire _04725_;
	wire _04726_;
	wire _04727_;
	wire _04728_;
	wire _04729_;
	wire _04730_;
	wire _04731_;
	wire _04732_;
	wire _04733_;
	wire _04734_;
	wire _04735_;
	wire _04736_;
	wire _04737_;
	wire _04738_;
	wire _04739_;
	wire _04740_;
	wire _04741_;
	wire _04742_;
	wire _04743_;
	wire _04744_;
	wire _04745_;
	wire _04746_;
	wire _04747_;
	wire _04748_;
	wire _04749_;
	wire _04750_;
	wire _04751_;
	wire _04752_;
	wire _04753_;
	wire _04754_;
	wire _04755_;
	wire _04756_;
	wire _04757_;
	wire _04758_;
	wire _04759_;
	wire _04760_;
	wire _04761_;
	wire _04762_;
	wire _04763_;
	wire _04764_;
	wire _04765_;
	wire _04766_;
	wire _04767_;
	wire _04768_;
	wire _04769_;
	wire _04770_;
	wire _04771_;
	wire _04772_;
	wire _04773_;
	wire _04774_;
	wire _04775_;
	wire _04776_;
	wire _04777_;
	wire _04778_;
	wire _04779_;
	wire _04780_;
	wire _04781_;
	wire _04782_;
	wire _04783_;
	wire _04784_;
	wire _04785_;
	wire _04786_;
	wire _04787_;
	wire _04788_;
	wire _04789_;
	wire _04790_;
	wire _04791_;
	wire _04792_;
	wire _04793_;
	wire _04794_;
	wire _04795_;
	wire _04796_;
	wire _04797_;
	wire _04798_;
	wire _04799_;
	wire _04800_;
	wire _04801_;
	wire _04802_;
	wire _04803_;
	wire _04804_;
	wire _04805_;
	wire _04806_;
	wire _04807_;
	wire _04808_;
	wire _04809_;
	wire _04810_;
	wire _04811_;
	wire _04812_;
	wire _04813_;
	wire _04814_;
	wire _04815_;
	wire _04816_;
	wire _04817_;
	wire _04818_;
	wire _04819_;
	wire _04820_;
	wire _04821_;
	wire _04822_;
	wire _04823_;
	wire _04824_;
	wire _04825_;
	wire _04826_;
	wire _04827_;
	wire _04828_;
	wire _04829_;
	wire _04830_;
	wire _04831_;
	wire _04832_;
	wire _04833_;
	wire _04834_;
	wire _04835_;
	wire _04836_;
	wire _04837_;
	wire _04838_;
	wire _04839_;
	wire _04840_;
	wire _04841_;
	wire _04842_;
	wire _04843_;
	wire _04844_;
	wire _04845_;
	wire _04846_;
	wire _04847_;
	wire _04848_;
	wire _04849_;
	wire _04850_;
	wire _04851_;
	wire _04852_;
	wire _04853_;
	wire _04854_;
	wire _04855_;
	wire _04856_;
	wire _04857_;
	wire _04858_;
	wire _04859_;
	wire _04860_;
	wire _04861_;
	wire _04862_;
	wire _04863_;
	wire _04864_;
	wire _04865_;
	wire _04866_;
	wire _04867_;
	wire _04868_;
	wire _04869_;
	wire _04870_;
	wire _04871_;
	wire _04872_;
	wire _04873_;
	wire _04874_;
	wire _04875_;
	wire _04876_;
	wire _04877_;
	wire _04878_;
	wire _04879_;
	wire _04880_;
	wire _04881_;
	wire _04882_;
	wire _04883_;
	wire _04884_;
	wire _04885_;
	wire _04886_;
	wire _04887_;
	wire _04888_;
	wire _04889_;
	wire _04890_;
	wire _04891_;
	wire _04892_;
	wire _04893_;
	wire _04894_;
	wire _04895_;
	wire _04896_;
	wire _04897_;
	wire _04898_;
	wire _04899_;
	wire _04900_;
	wire _04901_;
	wire _04902_;
	wire _04903_;
	wire _04904_;
	wire _04905_;
	wire _04906_;
	wire _04907_;
	wire _04908_;
	wire _04909_;
	wire _04910_;
	wire _04911_;
	wire _04912_;
	wire _04913_;
	wire _04914_;
	wire _04915_;
	wire _04916_;
	wire _04917_;
	wire _04918_;
	wire _04919_;
	wire _04920_;
	wire _04921_;
	wire _04922_;
	wire _04923_;
	wire _04924_;
	wire _04925_;
	wire _04926_;
	wire _04927_;
	wire _04928_;
	wire _04929_;
	wire _04930_;
	wire _04931_;
	wire _04932_;
	wire _04933_;
	wire _04934_;
	wire _04935_;
	wire _04936_;
	wire _04937_;
	wire _04938_;
	wire _04939_;
	wire _04940_;
	wire _04941_;
	wire _04942_;
	wire _04943_;
	wire _04944_;
	wire _04945_;
	wire _04946_;
	wire _04947_;
	wire _04948_;
	wire _04949_;
	wire _04950_;
	wire _04951_;
	wire _04952_;
	wire _04953_;
	wire _04954_;
	wire _04955_;
	wire _04956_;
	wire _04957_;
	wire _04958_;
	wire _04959_;
	wire _04960_;
	wire _04961_;
	wire _04962_;
	wire _04963_;
	wire _04964_;
	wire _04965_;
	wire _04966_;
	wire _04967_;
	wire _04968_;
	wire _04969_;
	wire _04970_;
	wire _04971_;
	wire _04972_;
	wire _04973_;
	wire _04974_;
	wire _04975_;
	wire _04976_;
	wire _04977_;
	wire _04978_;
	wire _04979_;
	wire _04980_;
	wire _04981_;
	wire _04982_;
	wire _04983_;
	wire _04984_;
	wire _04985_;
	wire _04986_;
	wire _04987_;
	wire _04988_;
	wire _04989_;
	wire _04990_;
	wire _04991_;
	wire _04992_;
	wire _04993_;
	wire _04994_;
	wire _04995_;
	wire _04996_;
	wire _04997_;
	wire _04998_;
	wire _04999_;
	wire _05000_;
	wire _05001_;
	wire _05002_;
	wire _05003_;
	wire _05004_;
	wire _05005_;
	wire _05006_;
	wire _05007_;
	wire _05008_;
	wire _05009_;
	wire _05010_;
	wire _05011_;
	wire _05012_;
	wire _05013_;
	wire _05014_;
	wire _05015_;
	wire _05016_;
	wire _05017_;
	wire _05018_;
	wire _05019_;
	wire _05020_;
	wire _05021_;
	wire _05022_;
	wire _05023_;
	wire _05024_;
	wire _05025_;
	wire _05026_;
	wire _05027_;
	wire _05028_;
	wire _05029_;
	wire _05030_;
	wire _05031_;
	wire _05032_;
	wire _05033_;
	wire _05034_;
	wire _05035_;
	wire _05036_;
	wire _05037_;
	wire _05038_;
	wire _05039_;
	wire _05040_;
	wire _05041_;
	wire _05042_;
	wire _05043_;
	wire _05044_;
	wire _05045_;
	wire _05046_;
	wire _05047_;
	wire _05048_;
	wire _05049_;
	wire _05050_;
	wire _05051_;
	wire _05052_;
	wire _05053_;
	wire _05054_;
	wire _05055_;
	wire _05056_;
	wire _05057_;
	wire _05058_;
	wire _05059_;
	wire _05060_;
	wire _05061_;
	wire _05062_;
	wire _05063_;
	wire _05064_;
	wire _05065_;
	wire _05066_;
	wire _05067_;
	wire _05068_;
	wire _05069_;
	wire _05070_;
	wire _05071_;
	wire _05072_;
	wire _05073_;
	wire _05074_;
	wire _05075_;
	wire _05076_;
	wire _05077_;
	wire _05078_;
	wire _05079_;
	wire _05080_;
	wire _05081_;
	wire _05082_;
	wire _05083_;
	wire _05084_;
	wire _05085_;
	wire _05086_;
	wire _05087_;
	wire _05088_;
	wire _05089_;
	wire _05090_;
	wire _05091_;
	wire _05092_;
	wire _05093_;
	wire _05094_;
	wire _05095_;
	wire _05096_;
	wire _05097_;
	wire _05098_;
	wire _05099_;
	wire _05100_;
	wire _05101_;
	wire _05102_;
	wire _05103_;
	wire _05104_;
	wire _05105_;
	wire _05106_;
	wire _05107_;
	wire _05108_;
	wire _05109_;
	wire _05110_;
	wire _05111_;
	wire _05112_;
	wire _05113_;
	wire _05114_;
	wire _05115_;
	wire _05116_;
	wire _05117_;
	wire _05118_;
	wire _05119_;
	wire _05120_;
	wire _05121_;
	wire _05122_;
	wire _05123_;
	wire _05124_;
	wire _05125_;
	wire _05126_;
	wire _05127_;
	wire _05128_;
	wire _05129_;
	wire _05130_;
	wire _05131_;
	wire _05132_;
	wire _05133_;
	wire _05134_;
	wire _05135_;
	wire _05136_;
	wire _05137_;
	wire _05138_;
	wire _05139_;
	wire _05140_;
	wire _05141_;
	wire _05142_;
	wire _05143_;
	wire _05144_;
	wire _05145_;
	wire _05146_;
	wire _05147_;
	wire _05148_;
	wire _05149_;
	wire _05150_;
	wire _05151_;
	wire _05152_;
	wire _05153_;
	wire _05154_;
	wire _05155_;
	wire _05156_;
	wire _05157_;
	wire _05158_;
	wire _05159_;
	wire _05160_;
	wire _05161_;
	wire _05162_;
	wire _05163_;
	wire _05164_;
	wire _05165_;
	wire _05166_;
	wire _05167_;
	wire _05168_;
	wire _05169_;
	wire _05170_;
	wire _05171_;
	wire _05172_;
	wire _05173_;
	wire _05174_;
	wire _05175_;
	wire _05176_;
	wire _05177_;
	wire _05178_;
	wire _05179_;
	wire _05180_;
	wire _05181_;
	wire _05182_;
	wire _05183_;
	wire _05184_;
	wire _05185_;
	wire _05186_;
	wire _05187_;
	wire _05188_;
	wire _05189_;
	wire _05190_;
	wire _05191_;
	wire _05192_;
	wire _05193_;
	wire _05194_;
	wire _05195_;
	wire _05196_;
	wire _05197_;
	wire _05198_;
	wire _05199_;
	wire _05200_;
	wire _05201_;
	wire _05202_;
	wire _05203_;
	wire _05204_;
	wire _05205_;
	wire _05206_;
	wire _05207_;
	wire _05208_;
	wire _05209_;
	wire _05210_;
	wire _05211_;
	wire _05212_;
	wire _05213_;
	wire _05214_;
	wire _05215_;
	wire _05216_;
	wire _05217_;
	wire _05218_;
	wire _05219_;
	wire _05220_;
	wire _05221_;
	wire _05222_;
	wire _05223_;
	wire _05224_;
	wire _05225_;
	wire _05226_;
	wire _05227_;
	wire _05228_;
	wire _05229_;
	wire _05230_;
	wire _05231_;
	wire _05232_;
	wire _05233_;
	wire _05234_;
	wire _05235_;
	wire _05236_;
	wire _05237_;
	wire _05238_;
	wire _05239_;
	wire _05240_;
	wire _05241_;
	wire _05242_;
	wire _05243_;
	wire _05244_;
	wire _05245_;
	wire _05246_;
	wire _05247_;
	wire _05248_;
	wire _05249_;
	wire _05250_;
	wire _05251_;
	wire _05252_;
	wire _05253_;
	wire _05254_;
	wire _05255_;
	wire _05256_;
	wire _05257_;
	wire _05258_;
	wire _05259_;
	wire _05260_;
	wire _05261_;
	wire _05262_;
	wire _05263_;
	wire _05264_;
	wire _05265_;
	wire _05266_;
	wire _05267_;
	wire _05268_;
	wire _05269_;
	wire _05270_;
	wire _05271_;
	wire _05272_;
	wire _05273_;
	wire _05274_;
	wire _05275_;
	wire _05276_;
	wire _05277_;
	wire _05278_;
	wire _05279_;
	wire _05280_;
	wire _05281_;
	wire _05282_;
	wire _05283_;
	wire _05284_;
	wire _05285_;
	wire _05286_;
	wire _05287_;
	wire _05288_;
	wire _05289_;
	wire _05290_;
	wire _05291_;
	wire _05292_;
	wire _05293_;
	wire _05294_;
	wire _05295_;
	wire _05296_;
	wire _05297_;
	wire _05298_;
	wire _05299_;
	wire _05300_;
	wire _05301_;
	wire _05302_;
	wire _05303_;
	wire _05304_;
	wire _05305_;
	wire _05306_;
	wire _05307_;
	wire _05308_;
	wire _05309_;
	wire _05310_;
	wire _05311_;
	wire _05312_;
	wire _05313_;
	wire _05314_;
	wire _05315_;
	wire _05316_;
	wire _05317_;
	wire _05318_;
	wire _05319_;
	wire _05320_;
	wire _05321_;
	wire _05322_;
	wire _05323_;
	wire _05324_;
	wire _05325_;
	wire _05326_;
	wire _05327_;
	wire _05328_;
	wire _05329_;
	wire _05330_;
	wire _05331_;
	wire _05332_;
	wire _05333_;
	wire _05334_;
	wire _05335_;
	wire _05336_;
	wire _05337_;
	wire _05338_;
	wire _05339_;
	wire _05340_;
	wire _05341_;
	wire _05342_;
	wire _05343_;
	wire _05344_;
	wire _05345_;
	wire _05346_;
	wire _05347_;
	wire _05348_;
	wire _05349_;
	wire _05350_;
	wire _05351_;
	wire _05352_;
	wire _05353_;
	wire _05354_;
	wire _05355_;
	wire _05356_;
	wire _05357_;
	wire _05358_;
	wire _05359_;
	wire _05360_;
	wire _05361_;
	wire _05362_;
	wire _05363_;
	wire _05364_;
	wire _05365_;
	wire _05366_;
	wire _05367_;
	wire _05368_;
	wire _05369_;
	wire _05370_;
	wire _05371_;
	wire _05372_;
	wire _05373_;
	wire _05374_;
	wire _05375_;
	wire _05376_;
	wire _05377_;
	wire _05378_;
	wire _05379_;
	wire _05380_;
	wire _05381_;
	wire _05382_;
	wire _05383_;
	wire _05384_;
	wire _05385_;
	wire _05386_;
	wire _05387_;
	wire _05388_;
	wire _05389_;
	wire _05390_;
	wire _05391_;
	wire _05392_;
	wire _05393_;
	wire _05394_;
	wire _05395_;
	wire _05396_;
	wire _05397_;
	wire _05398_;
	wire _05399_;
	wire _05400_;
	wire _05401_;
	wire _05402_;
	wire _05403_;
	wire _05404_;
	wire _05405_;
	wire _05406_;
	wire _05407_;
	wire _05408_;
	wire _05409_;
	wire _05410_;
	wire _05411_;
	wire _05412_;
	wire _05413_;
	wire _05414_;
	wire _05415_;
	wire _05416_;
	wire _05417_;
	wire _05418_;
	wire _05419_;
	wire _05420_;
	wire _05421_;
	wire _05422_;
	wire _05423_;
	wire _05424_;
	wire _05425_;
	wire _05426_;
	wire _05427_;
	wire _05428_;
	wire _05429_;
	wire _05430_;
	wire _05431_;
	wire _05432_;
	wire _05433_;
	wire _05434_;
	wire _05435_;
	wire _05436_;
	wire _05437_;
	wire _05438_;
	wire _05439_;
	wire _05440_;
	wire _05441_;
	wire _05442_;
	wire _05443_;
	wire _05444_;
	wire _05445_;
	wire _05446_;
	wire _05447_;
	wire _05448_;
	wire _05449_;
	wire _05450_;
	wire _05451_;
	wire _05452_;
	wire _05453_;
	wire _05454_;
	wire _05455_;
	wire _05456_;
	wire _05457_;
	wire _05458_;
	wire _05459_;
	wire _05460_;
	wire _05461_;
	wire _05462_;
	wire _05463_;
	wire _05464_;
	wire _05465_;
	wire _05466_;
	wire _05467_;
	wire _05468_;
	wire _05469_;
	wire _05470_;
	wire _05471_;
	wire _05472_;
	wire _05473_;
	wire _05474_;
	wire _05475_;
	wire _05476_;
	wire _05477_;
	wire _05478_;
	wire _05479_;
	wire _05480_;
	wire _05481_;
	wire _05482_;
	wire _05483_;
	wire _05484_;
	wire _05485_;
	wire _05486_;
	wire _05487_;
	wire _05488_;
	wire _05489_;
	wire _05490_;
	wire _05491_;
	wire _05492_;
	wire _05493_;
	wire _05494_;
	wire _05495_;
	wire _05496_;
	wire _05497_;
	wire _05498_;
	wire _05499_;
	wire _05500_;
	wire _05501_;
	wire _05502_;
	wire _05503_;
	wire _05504_;
	wire _05505_;
	wire _05506_;
	wire _05507_;
	wire _05508_;
	wire _05509_;
	wire _05510_;
	wire _05511_;
	wire _05512_;
	wire _05513_;
	wire _05514_;
	wire _05515_;
	wire _05516_;
	wire _05517_;
	wire _05518_;
	wire _05519_;
	wire _05520_;
	wire _05521_;
	wire _05522_;
	wire _05523_;
	wire _05524_;
	wire _05525_;
	wire _05526_;
	wire _05527_;
	wire _05528_;
	wire _05529_;
	wire _05530_;
	wire _05531_;
	wire _05532_;
	wire _05533_;
	wire _05534_;
	wire _05535_;
	wire _05536_;
	wire _05537_;
	wire _05538_;
	wire _05539_;
	wire _05540_;
	wire _05541_;
	wire _05542_;
	wire _05543_;
	wire _05544_;
	wire _05545_;
	wire _05546_;
	wire _05547_;
	wire _05548_;
	wire _05549_;
	wire _05550_;
	wire _05551_;
	wire _05552_;
	wire _05553_;
	wire _05554_;
	wire _05555_;
	wire _05556_;
	wire _05557_;
	wire _05558_;
	wire _05559_;
	wire _05560_;
	wire _05561_;
	wire _05562_;
	wire _05563_;
	wire _05564_;
	wire _05565_;
	wire _05566_;
	wire _05567_;
	wire _05568_;
	wire _05569_;
	wire _05570_;
	wire _05571_;
	wire _05572_;
	wire _05573_;
	wire _05574_;
	wire _05575_;
	wire _05576_;
	wire _05577_;
	wire _05578_;
	wire _05579_;
	wire _05580_;
	wire _05581_;
	wire _05582_;
	wire _05583_;
	wire _05584_;
	wire _05585_;
	wire _05586_;
	wire _05587_;
	wire _05588_;
	wire _05589_;
	wire _05590_;
	wire _05591_;
	wire _05592_;
	wire _05593_;
	wire _05594_;
	wire _05595_;
	wire _05596_;
	wire _05597_;
	wire _05598_;
	wire _05599_;
	wire _05600_;
	wire _05601_;
	wire _05602_;
	wire _05603_;
	wire _05604_;
	wire _05605_;
	wire _05606_;
	wire _05607_;
	wire _05608_;
	wire _05609_;
	wire _05610_;
	wire _05611_;
	wire _05612_;
	wire _05613_;
	wire _05614_;
	wire _05615_;
	wire _05616_;
	wire _05617_;
	wire _05618_;
	wire _05619_;
	wire _05620_;
	wire _05621_;
	wire _05622_;
	wire _05623_;
	wire _05624_;
	wire _05625_;
	wire _05626_;
	wire _05627_;
	wire _05628_;
	wire _05629_;
	wire _05630_;
	wire _05631_;
	wire _05632_;
	wire _05633_;
	wire _05634_;
	wire _05635_;
	wire _05636_;
	wire _05637_;
	wire _05638_;
	wire _05639_;
	wire _05640_;
	wire _05641_;
	wire _05642_;
	wire _05643_;
	wire _05644_;
	wire _05645_;
	wire _05646_;
	wire _05647_;
	wire _05648_;
	wire _05649_;
	wire _05650_;
	wire _05651_;
	wire _05652_;
	wire _05653_;
	wire _05654_;
	wire _05655_;
	wire _05656_;
	wire _05657_;
	wire _05658_;
	wire _05659_;
	wire _05660_;
	wire _05661_;
	wire _05662_;
	wire _05663_;
	wire _05664_;
	wire _05665_;
	wire _05666_;
	wire _05667_;
	wire _05668_;
	wire _05669_;
	wire _05670_;
	wire _05671_;
	wire _05672_;
	wire _05673_;
	wire _05674_;
	wire _05675_;
	wire _05676_;
	wire _05677_;
	wire _05678_;
	wire _05679_;
	wire _05680_;
	wire _05681_;
	wire _05682_;
	wire _05683_;
	wire _05684_;
	wire _05685_;
	wire _05686_;
	wire _05687_;
	wire _05688_;
	wire _05689_;
	wire _05690_;
	wire _05691_;
	wire _05692_;
	wire _05693_;
	wire _05694_;
	wire _05695_;
	wire _05696_;
	wire _05697_;
	wire _05698_;
	wire _05699_;
	wire _05700_;
	wire _05701_;
	wire _05702_;
	wire _05703_;
	wire _05704_;
	wire _05705_;
	wire _05706_;
	wire _05707_;
	wire _05708_;
	wire _05709_;
	wire _05710_;
	wire _05711_;
	wire _05712_;
	wire _05713_;
	wire _05714_;
	wire _05715_;
	wire _05716_;
	wire _05717_;
	wire _05718_;
	wire _05719_;
	wire _05720_;
	wire _05721_;
	wire _05722_;
	wire _05723_;
	wire _05724_;
	wire _05725_;
	wire _05726_;
	wire _05727_;
	wire _05728_;
	wire _05729_;
	wire _05730_;
	wire _05731_;
	wire _05732_;
	wire _05733_;
	wire _05734_;
	wire _05735_;
	wire _05736_;
	wire _05737_;
	wire _05738_;
	wire _05739_;
	wire _05740_;
	wire _05741_;
	wire _05742_;
	wire _05743_;
	wire _05744_;
	wire _05745_;
	wire _05746_;
	wire _05747_;
	wire _05748_;
	wire _05749_;
	wire _05750_;
	wire _05751_;
	wire _05752_;
	wire _05753_;
	wire _05754_;
	wire _05755_;
	wire _05756_;
	wire _05757_;
	wire _05758_;
	wire _05759_;
	wire _05760_;
	wire _05761_;
	wire _05762_;
	wire _05763_;
	wire _05764_;
	wire _05765_;
	wire _05766_;
	wire _05767_;
	wire _05768_;
	wire _05769_;
	wire _05770_;
	wire _05771_;
	wire _05772_;
	wire _05773_;
	wire _05774_;
	wire _05775_;
	wire _05776_;
	wire _05777_;
	wire _05778_;
	wire _05779_;
	wire _05780_;
	wire _05781_;
	wire _05782_;
	wire _05783_;
	wire _05784_;
	wire _05785_;
	wire _05786_;
	wire _05787_;
	wire _05788_;
	wire _05789_;
	wire _05790_;
	wire _05791_;
	wire _05792_;
	wire _05793_;
	wire _05794_;
	wire _05795_;
	wire _05796_;
	wire _05797_;
	wire _05798_;
	wire _05799_;
	wire _05800_;
	wire _05801_;
	wire _05802_;
	wire _05803_;
	wire _05804_;
	wire _05805_;
	wire _05806_;
	wire _05807_;
	wire _05808_;
	wire _05809_;
	wire _05810_;
	wire _05811_;
	wire _05812_;
	wire _05813_;
	wire _05814_;
	wire _05815_;
	wire _05816_;
	wire _05817_;
	wire _05818_;
	wire _05819_;
	wire _05820_;
	wire _05821_;
	wire _05822_;
	wire _05823_;
	wire _05824_;
	wire _05825_;
	wire _05826_;
	wire _05827_;
	wire _05828_;
	wire _05829_;
	wire _05830_;
	wire _05831_;
	wire _05832_;
	wire _05833_;
	wire _05834_;
	wire _05835_;
	wire _05836_;
	wire _05837_;
	wire _05838_;
	wire _05839_;
	wire _05840_;
	wire _05841_;
	wire _05842_;
	wire _05843_;
	wire _05844_;
	wire _05845_;
	wire _05846_;
	wire _05847_;
	wire _05848_;
	wire _05849_;
	wire _05850_;
	wire _05851_;
	wire _05852_;
	wire _05853_;
	wire _05854_;
	wire _05855_;
	wire _05856_;
	wire _05857_;
	wire _05858_;
	wire _05859_;
	wire _05860_;
	wire _05861_;
	wire _05862_;
	wire _05863_;
	wire _05864_;
	wire _05865_;
	wire _05866_;
	wire _05867_;
	wire _05868_;
	wire _05869_;
	wire _05870_;
	wire _05871_;
	wire _05872_;
	wire _05873_;
	wire _05874_;
	wire _05875_;
	wire _05876_;
	wire _05877_;
	wire _05878_;
	wire _05879_;
	wire _05880_;
	wire _05881_;
	wire _05882_;
	wire _05883_;
	wire _05884_;
	wire _05885_;
	wire _05886_;
	wire _05887_;
	wire _05888_;
	wire _05889_;
	wire _05890_;
	wire _05891_;
	wire _05892_;
	wire _05893_;
	wire _05894_;
	wire _05895_;
	wire _05896_;
	wire _05897_;
	wire _05898_;
	wire _05899_;
	wire _05900_;
	wire _05901_;
	wire _05902_;
	wire _05903_;
	wire _05904_;
	wire _05905_;
	wire _05906_;
	wire _05907_;
	wire _05908_;
	wire _05909_;
	wire _05910_;
	wire _05911_;
	wire _05912_;
	wire _05913_;
	wire _05914_;
	wire _05915_;
	wire _05916_;
	wire _05917_;
	wire _05918_;
	wire _05919_;
	wire _05920_;
	wire _05921_;
	wire _05922_;
	wire _05923_;
	wire _05924_;
	wire _05925_;
	wire _05926_;
	wire _05927_;
	wire _05928_;
	wire _05929_;
	wire _05930_;
	wire _05931_;
	wire _05932_;
	wire _05933_;
	wire _05934_;
	wire _05935_;
	wire _05936_;
	wire _05937_;
	wire _05938_;
	wire _05939_;
	wire _05940_;
	wire _05941_;
	wire _05942_;
	wire _05943_;
	wire _05944_;
	wire _05945_;
	wire _05946_;
	wire _05947_;
	wire _05948_;
	wire _05949_;
	wire _05950_;
	wire _05951_;
	wire _05952_;
	wire _05953_;
	wire _05954_;
	wire _05955_;
	wire _05956_;
	wire _05957_;
	wire _05958_;
	wire _05959_;
	wire _05960_;
	wire _05961_;
	wire _05962_;
	wire _05963_;
	wire _05964_;
	wire _05965_;
	wire _05966_;
	wire _05967_;
	wire _05968_;
	wire _05969_;
	wire _05970_;
	wire _05971_;
	wire _05972_;
	wire _05973_;
	wire _05974_;
	wire _05975_;
	wire _05976_;
	wire _05977_;
	wire _05978_;
	wire _05979_;
	wire _05980_;
	wire _05981_;
	wire _05982_;
	wire _05983_;
	wire _05984_;
	wire _05985_;
	wire _05986_;
	wire _05987_;
	wire _05988_;
	wire _05989_;
	wire _05990_;
	wire _05991_;
	wire _05992_;
	wire _05993_;
	wire _05994_;
	wire _05995_;
	wire _05996_;
	wire _05997_;
	wire _05998_;
	wire _05999_;
	wire _06000_;
	wire _06001_;
	wire _06002_;
	wire _06003_;
	wire _06004_;
	wire _06005_;
	wire _06006_;
	wire _06007_;
	wire _06008_;
	wire _06009_;
	wire _06010_;
	wire _06011_;
	wire _06012_;
	wire _06013_;
	wire _06014_;
	wire _06015_;
	wire _06016_;
	wire _06017_;
	wire _06018_;
	wire _06019_;
	wire _06020_;
	wire _06021_;
	wire _06022_;
	wire _06023_;
	wire _06024_;
	wire _06025_;
	wire _06026_;
	wire _06027_;
	wire _06028_;
	wire _06029_;
	wire _06030_;
	wire _06031_;
	wire _06032_;
	wire _06033_;
	wire _06034_;
	wire _06035_;
	wire _06036_;
	wire _06037_;
	wire _06038_;
	wire _06039_;
	wire _06040_;
	wire _06041_;
	wire _06042_;
	wire _06043_;
	wire _06044_;
	wire _06045_;
	wire _06046_;
	wire _06047_;
	wire _06048_;
	wire _06049_;
	wire _06050_;
	wire _06051_;
	wire _06052_;
	wire _06053_;
	wire _06054_;
	wire _06055_;
	wire _06056_;
	wire _06057_;
	wire _06058_;
	wire _06059_;
	wire _06060_;
	wire _06061_;
	wire _06062_;
	wire _06063_;
	wire _06064_;
	wire _06065_;
	wire _06066_;
	wire _06067_;
	wire _06068_;
	wire _06069_;
	wire _06070_;
	wire _06071_;
	wire _06072_;
	wire _06073_;
	wire _06074_;
	wire _06075_;
	wire _06076_;
	wire _06077_;
	wire _06078_;
	wire _06079_;
	wire _06080_;
	wire _06081_;
	wire _06082_;
	wire _06083_;
	wire _06084_;
	wire _06085_;
	wire _06086_;
	wire _06087_;
	wire _06088_;
	wire _06089_;
	wire _06090_;
	wire _06091_;
	wire _06092_;
	wire _06093_;
	wire _06094_;
	wire _06095_;
	wire _06096_;
	wire _06097_;
	wire _06098_;
	wire _06099_;
	wire _06100_;
	wire _06101_;
	wire _06102_;
	wire _06103_;
	wire _06104_;
	wire _06105_;
	wire _06106_;
	wire _06107_;
	wire _06108_;
	wire _06109_;
	wire _06110_;
	wire _06111_;
	wire _06112_;
	wire _06113_;
	wire _06114_;
	wire _06115_;
	wire _06116_;
	wire _06117_;
	wire _06118_;
	wire _06119_;
	wire _06120_;
	wire _06121_;
	wire _06122_;
	wire _06123_;
	wire _06124_;
	wire _06125_;
	wire _06126_;
	wire _06127_;
	wire _06128_;
	wire _06129_;
	wire _06130_;
	wire _06131_;
	wire _06132_;
	wire _06133_;
	wire _06134_;
	wire _06135_;
	wire _06136_;
	wire _06137_;
	wire _06138_;
	wire _06139_;
	wire _06140_;
	wire _06141_;
	wire _06142_;
	wire _06143_;
	wire _06144_;
	wire _06145_;
	wire _06146_;
	wire _06147_;
	wire _06148_;
	wire _06149_;
	wire _06150_;
	wire _06151_;
	wire _06152_;
	wire _06153_;
	wire _06154_;
	wire _06155_;
	wire _06156_;
	wire _06157_;
	wire _06158_;
	wire _06159_;
	wire _06160_;
	wire _06161_;
	wire _06162_;
	wire _06163_;
	wire _06164_;
	wire _06165_;
	wire _06166_;
	wire _06167_;
	wire _06168_;
	wire _06169_;
	wire _06170_;
	wire _06171_;
	wire _06172_;
	wire _06173_;
	wire _06174_;
	wire _06175_;
	wire _06176_;
	wire _06177_;
	wire _06178_;
	wire _06179_;
	wire _06180_;
	wire _06181_;
	wire _06182_;
	wire _06183_;
	wire _06184_;
	wire _06185_;
	wire _06186_;
	wire _06187_;
	wire _06188_;
	wire _06189_;
	wire _06190_;
	wire _06191_;
	wire _06192_;
	wire _06193_;
	wire _06194_;
	wire _06195_;
	wire _06196_;
	wire _06197_;
	wire _06198_;
	wire _06199_;
	wire _06200_;
	wire _06201_;
	wire _06202_;
	wire _06203_;
	wire _06204_;
	wire _06205_;
	wire _06206_;
	wire _06207_;
	wire _06208_;
	wire _06209_;
	wire _06210_;
	wire _06211_;
	wire _06212_;
	wire _06213_;
	wire _06214_;
	wire _06215_;
	wire _06216_;
	wire _06217_;
	wire _06218_;
	wire _06219_;
	wire _06220_;
	wire _06221_;
	wire _06222_;
	wire _06223_;
	wire _06224_;
	wire _06225_;
	wire _06226_;
	wire _06227_;
	wire _06228_;
	wire _06229_;
	wire _06230_;
	wire _06231_;
	wire _06232_;
	wire _06233_;
	wire _06234_;
	wire _06235_;
	wire _06236_;
	wire _06237_;
	wire _06238_;
	wire _06239_;
	wire _06240_;
	wire _06241_;
	wire _06242_;
	wire _06243_;
	wire _06244_;
	wire _06245_;
	wire _06246_;
	wire _06247_;
	wire _06248_;
	wire _06249_;
	wire _06250_;
	wire _06251_;
	wire _06252_;
	wire _06253_;
	wire _06254_;
	wire _06255_;
	wire _06256_;
	wire _06257_;
	wire _06258_;
	wire _06259_;
	wire _06260_;
	wire _06261_;
	wire _06262_;
	wire _06263_;
	wire _06264_;
	wire _06265_;
	wire _06266_;
	wire _06267_;
	wire _06268_;
	wire _06269_;
	wire _06270_;
	wire _06271_;
	wire _06272_;
	wire _06273_;
	wire _06274_;
	wire _06275_;
	wire _06276_;
	wire _06277_;
	wire _06278_;
	wire _06279_;
	wire _06280_;
	wire _06281_;
	wire _06282_;
	wire _06283_;
	wire _06284_;
	wire _06285_;
	wire _06286_;
	wire _06287_;
	wire _06288_;
	wire _06289_;
	wire _06290_;
	wire _06291_;
	wire _06292_;
	wire _06293_;
	wire _06294_;
	wire _06295_;
	wire _06296_;
	wire _06297_;
	wire _06298_;
	wire _06299_;
	wire _06300_;
	wire _06301_;
	wire _06302_;
	wire _06303_;
	wire _06304_;
	wire _06305_;
	wire _06306_;
	wire _06307_;
	wire _06308_;
	wire _06309_;
	wire _06310_;
	wire _06311_;
	wire _06312_;
	wire _06313_;
	wire _06314_;
	wire _06315_;
	wire _06316_;
	wire _06317_;
	wire _06318_;
	wire _06319_;
	wire _06320_;
	wire _06321_;
	wire _06322_;
	wire _06323_;
	wire _06324_;
	wire _06325_;
	wire _06326_;
	wire _06327_;
	wire _06328_;
	wire _06329_;
	wire _06330_;
	wire _06331_;
	wire _06332_;
	wire _06333_;
	wire _06334_;
	wire _06335_;
	wire _06336_;
	wire _06337_;
	wire _06338_;
	wire _06339_;
	wire _06340_;
	wire _06341_;
	wire _06342_;
	wire _06343_;
	wire _06344_;
	wire _06345_;
	wire _06346_;
	wire _06347_;
	wire _06348_;
	wire _06349_;
	wire _06350_;
	wire _06351_;
	wire _06352_;
	wire _06353_;
	wire _06354_;
	wire _06355_;
	wire _06356_;
	wire _06357_;
	wire _06358_;
	wire _06359_;
	wire _06360_;
	wire _06361_;
	wire _06362_;
	wire _06363_;
	wire _06364_;
	wire _06365_;
	wire _06366_;
	wire _06367_;
	wire _06368_;
	wire _06369_;
	wire _06370_;
	wire _06371_;
	wire _06372_;
	wire _06373_;
	wire _06374_;
	wire _06375_;
	wire _06376_;
	wire _06377_;
	wire _06378_;
	wire _06379_;
	wire _06380_;
	wire _06381_;
	wire _06382_;
	wire _06383_;
	wire _06384_;
	wire _06385_;
	wire _06386_;
	wire _06387_;
	wire _06388_;
	wire _06389_;
	wire _06390_;
	wire _06391_;
	wire _06392_;
	wire _06393_;
	wire _06394_;
	wire _06395_;
	wire _06396_;
	wire _06397_;
	wire _06398_;
	wire _06399_;
	wire _06400_;
	wire _06401_;
	wire _06402_;
	wire _06403_;
	wire _06404_;
	wire _06405_;
	wire _06406_;
	wire _06407_;
	wire _06408_;
	wire _06409_;
	wire _06410_;
	wire _06411_;
	wire _06412_;
	wire _06413_;
	wire _06414_;
	wire _06415_;
	wire _06416_;
	wire _06417_;
	wire _06418_;
	wire _06419_;
	wire _06420_;
	wire _06421_;
	wire _06422_;
	wire _06423_;
	wire _06424_;
	wire _06425_;
	wire _06426_;
	wire _06427_;
	wire _06428_;
	wire _06429_;
	wire _06430_;
	wire _06431_;
	wire _06432_;
	wire _06433_;
	wire _06434_;
	wire _06435_;
	wire _06436_;
	wire _06437_;
	wire _06438_;
	wire _06439_;
	wire _06440_;
	wire _06441_;
	wire _06442_;
	wire _06443_;
	wire _06444_;
	wire _06445_;
	wire _06446_;
	wire _06447_;
	wire _06448_;
	wire _06449_;
	wire _06450_;
	wire _06451_;
	wire _06452_;
	wire _06453_;
	wire _06454_;
	wire _06455_;
	wire _06456_;
	wire _06457_;
	wire _06458_;
	wire _06459_;
	wire _06460_;
	wire _06461_;
	wire _06462_;
	wire _06463_;
	wire _06464_;
	wire _06465_;
	wire _06466_;
	wire _06467_;
	wire _06468_;
	wire _06469_;
	wire _06470_;
	wire _06471_;
	wire _06472_;
	wire _06473_;
	wire _06474_;
	wire _06475_;
	wire _06476_;
	wire _06477_;
	wire _06478_;
	wire _06479_;
	wire _06480_;
	wire _06481_;
	wire _06482_;
	wire _06483_;
	wire _06484_;
	wire _06485_;
	wire _06486_;
	wire _06487_;
	wire _06488_;
	wire _06489_;
	wire _06490_;
	wire _06491_;
	wire _06492_;
	wire _06493_;
	wire _06494_;
	wire _06495_;
	wire _06496_;
	wire _06497_;
	wire _06498_;
	wire _06499_;
	wire _06500_;
	wire _06501_;
	wire _06502_;
	wire _06503_;
	wire _06504_;
	wire _06505_;
	wire _06506_;
	wire _06507_;
	wire _06508_;
	wire _06509_;
	wire _06510_;
	wire _06511_;
	wire _06512_;
	wire _06513_;
	wire _06514_;
	wire _06515_;
	wire _06516_;
	wire _06517_;
	wire _06518_;
	wire _06519_;
	wire _06520_;
	wire _06521_;
	wire _06522_;
	wire _06523_;
	wire _06524_;
	wire _06525_;
	wire _06526_;
	wire _06527_;
	wire _06528_;
	wire _06529_;
	wire _06530_;
	wire _06531_;
	wire _06532_;
	wire _06533_;
	wire _06534_;
	wire _06535_;
	wire _06536_;
	wire _06537_;
	wire _06538_;
	wire _06539_;
	wire _06540_;
	wire _06541_;
	wire _06542_;
	wire _06543_;
	wire _06544_;
	wire _06545_;
	wire _06546_;
	wire _06547_;
	wire _06548_;
	wire _06549_;
	wire _06550_;
	wire _06551_;
	wire _06552_;
	wire _06553_;
	wire _06554_;
	wire _06555_;
	wire _06556_;
	wire _06557_;
	wire _06558_;
	wire _06559_;
	wire _06560_;
	wire _06561_;
	wire _06562_;
	wire _06563_;
	wire _06564_;
	wire _06565_;
	wire _06566_;
	wire _06567_;
	wire _06568_;
	wire _06569_;
	wire _06570_;
	wire _06571_;
	wire _06572_;
	wire _06573_;
	wire _06574_;
	wire _06575_;
	wire _06576_;
	wire _06577_;
	wire _06578_;
	wire _06579_;
	wire _06580_;
	wire _06581_;
	wire _06582_;
	wire _06583_;
	wire _06584_;
	wire _06585_;
	wire _06586_;
	wire _06587_;
	wire _06588_;
	wire _06589_;
	wire _06590_;
	wire _06591_;
	wire _06592_;
	wire _06593_;
	wire _06594_;
	wire _06595_;
	wire _06596_;
	wire _06597_;
	wire _06598_;
	wire _06599_;
	wire _06600_;
	wire _06601_;
	wire _06602_;
	wire _06603_;
	wire _06604_;
	wire _06605_;
	wire _06606_;
	wire _06607_;
	wire _06608_;
	wire _06609_;
	wire _06610_;
	wire _06611_;
	wire _06612_;
	wire _06613_;
	wire _06614_;
	wire _06615_;
	wire _06616_;
	wire _06617_;
	wire _06618_;
	wire _06619_;
	wire _06620_;
	wire _06621_;
	wire _06622_;
	wire _06623_;
	wire _06624_;
	wire _06625_;
	wire _06626_;
	wire _06627_;
	wire _06628_;
	wire _06629_;
	wire _06630_;
	wire _06631_;
	wire _06632_;
	wire _06633_;
	wire _06634_;
	wire _06635_;
	wire _06636_;
	wire _06637_;
	wire _06638_;
	wire _06639_;
	wire _06640_;
	wire _06641_;
	wire _06642_;
	wire _06643_;
	wire _06644_;
	wire _06645_;
	wire _06646_;
	wire _06647_;
	wire _06648_;
	wire _06649_;
	wire _06650_;
	wire _06651_;
	wire _06652_;
	wire _06653_;
	wire _06654_;
	wire _06655_;
	wire _06656_;
	wire _06657_;
	wire _06658_;
	wire _06659_;
	wire _06660_;
	wire _06661_;
	wire _06662_;
	wire _06663_;
	wire _06664_;
	wire _06665_;
	wire _06666_;
	wire _06667_;
	wire _06668_;
	wire _06669_;
	wire _06670_;
	wire _06671_;
	wire _06672_;
	wire _06673_;
	wire _06674_;
	wire _06675_;
	wire _06676_;
	wire _06677_;
	wire _06678_;
	wire _06679_;
	wire _06680_;
	wire _06681_;
	wire _06682_;
	wire _06683_;
	wire _06684_;
	wire _06685_;
	wire _06686_;
	wire _06687_;
	wire _06688_;
	wire _06689_;
	wire _06690_;
	wire _06691_;
	wire _06692_;
	wire _06693_;
	wire _06694_;
	wire _06695_;
	wire _06696_;
	wire _06697_;
	wire _06698_;
	wire _06699_;
	wire _06700_;
	wire _06701_;
	wire _06702_;
	wire _06703_;
	wire _06704_;
	wire _06705_;
	wire _06706_;
	wire _06707_;
	wire _06708_;
	wire _06709_;
	wire _06710_;
	wire _06711_;
	wire _06712_;
	wire _06713_;
	wire _06714_;
	wire _06715_;
	wire _06716_;
	wire _06717_;
	wire _06718_;
	wire _06719_;
	wire _06720_;
	wire _06721_;
	wire _06722_;
	wire _06723_;
	wire _06724_;
	wire _06725_;
	wire _06726_;
	wire _06727_;
	wire _06728_;
	wire _06729_;
	wire _06730_;
	wire _06731_;
	wire _06732_;
	wire _06733_;
	wire _06734_;
	wire _06735_;
	wire _06736_;
	wire _06737_;
	wire _06738_;
	wire _06739_;
	wire _06740_;
	wire _06741_;
	wire _06742_;
	wire _06743_;
	wire _06744_;
	wire _06745_;
	wire _06746_;
	wire _06747_;
	wire _06748_;
	wire _06749_;
	wire _06750_;
	wire _06751_;
	wire _06752_;
	wire _06753_;
	wire _06754_;
	wire _06755_;
	wire _06756_;
	wire _06757_;
	wire _06758_;
	wire _06759_;
	wire _06760_;
	wire _06761_;
	wire _06762_;
	wire _06763_;
	wire _06764_;
	wire _06765_;
	wire _06766_;
	wire _06767_;
	wire _06768_;
	wire _06769_;
	wire _06770_;
	wire _06771_;
	wire _06772_;
	wire _06773_;
	wire _06774_;
	wire _06775_;
	wire _06776_;
	wire _06777_;
	wire _06778_;
	wire _06779_;
	wire _06780_;
	wire _06781_;
	wire _06782_;
	wire _06783_;
	wire _06784_;
	wire _06785_;
	wire _06786_;
	wire _06787_;
	wire _06788_;
	wire _06789_;
	wire _06790_;
	wire _06791_;
	wire _06792_;
	wire _06793_;
	wire _06794_;
	wire _06795_;
	wire _06796_;
	wire _06797_;
	wire _06798_;
	wire _06799_;
	wire _06800_;
	wire _06801_;
	wire _06802_;
	wire _06803_;
	wire _06804_;
	wire _06805_;
	wire _06806_;
	wire _06807_;
	wire _06808_;
	wire _06809_;
	wire _06810_;
	wire _06811_;
	wire _06812_;
	wire _06813_;
	wire _06814_;
	wire _06815_;
	wire _06816_;
	wire _06817_;
	wire _06818_;
	wire _06819_;
	wire _06820_;
	wire _06821_;
	wire _06822_;
	wire _06823_;
	wire _06824_;
	wire _06825_;
	wire _06826_;
	wire _06827_;
	wire _06828_;
	wire _06829_;
	wire _06830_;
	wire _06831_;
	wire _06832_;
	wire _06833_;
	wire _06834_;
	wire _06835_;
	wire _06836_;
	wire _06837_;
	wire _06838_;
	wire _06839_;
	wire _06840_;
	wire _06841_;
	wire _06842_;
	wire _06843_;
	wire _06844_;
	wire _06845_;
	wire _06846_;
	wire _06847_;
	wire _06848_;
	wire _06849_;
	wire _06850_;
	wire _06851_;
	wire _06852_;
	wire _06853_;
	wire _06854_;
	wire _06855_;
	wire _06856_;
	wire _06857_;
	wire _06858_;
	wire _06859_;
	wire _06860_;
	wire _06861_;
	wire _06862_;
	wire _06863_;
	wire _06864_;
	wire _06865_;
	wire _06866_;
	wire _06867_;
	wire _06868_;
	wire _06869_;
	wire _06870_;
	wire _06871_;
	wire _06872_;
	wire _06873_;
	wire _06874_;
	wire _06875_;
	wire _06876_;
	wire _06877_;
	wire _06878_;
	wire _06879_;
	wire _06880_;
	wire _06881_;
	wire _06882_;
	wire _06883_;
	wire _06884_;
	wire _06885_;
	wire _06886_;
	wire _06887_;
	wire _06888_;
	wire _06889_;
	wire _06890_;
	wire _06891_;
	wire _06892_;
	wire _06893_;
	wire _06894_;
	wire _06895_;
	wire _06896_;
	wire _06897_;
	wire _06898_;
	wire _06899_;
	wire _06900_;
	wire _06901_;
	wire _06902_;
	wire _06903_;
	wire _06904_;
	wire _06905_;
	wire _06906_;
	wire _06907_;
	wire _06908_;
	wire _06909_;
	wire _06910_;
	wire _06911_;
	wire _06912_;
	wire _06913_;
	wire _06914_;
	wire _06915_;
	wire _06916_;
	wire _06917_;
	wire _06918_;
	wire _06919_;
	wire _06920_;
	wire _06921_;
	wire _06922_;
	wire _06923_;
	wire _06924_;
	wire _06925_;
	wire _06926_;
	wire _06927_;
	wire _06928_;
	wire _06929_;
	wire _06930_;
	wire _06931_;
	wire _06932_;
	wire _06933_;
	wire _06934_;
	wire _06935_;
	wire _06936_;
	wire _06937_;
	wire _06938_;
	wire _06939_;
	wire _06940_;
	wire _06941_;
	wire _06942_;
	wire _06943_;
	wire _06944_;
	wire _06945_;
	wire _06946_;
	wire _06947_;
	wire _06948_;
	wire _06949_;
	wire _06950_;
	wire _06951_;
	wire _06952_;
	wire _06953_;
	wire _06954_;
	wire _06955_;
	wire _06956_;
	wire _06957_;
	wire _06958_;
	wire _06959_;
	wire _06960_;
	wire _06961_;
	wire _06962_;
	wire _06963_;
	wire _06964_;
	wire _06965_;
	wire _06966_;
	wire _06967_;
	wire _06968_;
	wire _06969_;
	wire _06970_;
	wire _06971_;
	wire _06972_;
	wire _06973_;
	wire _06974_;
	wire _06975_;
	wire _06976_;
	wire _06977_;
	wire _06978_;
	wire _06979_;
	wire _06980_;
	wire _06981_;
	wire _06982_;
	wire _06983_;
	wire _06984_;
	wire _06985_;
	wire _06986_;
	wire _06987_;
	wire _06988_;
	wire _06989_;
	wire _06990_;
	wire _06991_;
	wire _06992_;
	wire _06993_;
	wire _06994_;
	wire _06995_;
	wire _06996_;
	wire _06997_;
	wire _06998_;
	wire _06999_;
	wire _07000_;
	wire _07001_;
	wire _07002_;
	wire _07003_;
	wire _07004_;
	wire _07005_;
	wire _07006_;
	wire _07007_;
	wire _07008_;
	wire _07009_;
	wire _07010_;
	wire _07011_;
	wire _07012_;
	wire _07013_;
	wire _07014_;
	wire _07015_;
	wire _07016_;
	wire _07017_;
	wire _07018_;
	wire _07019_;
	wire _07020_;
	wire _07021_;
	wire _07022_;
	wire _07023_;
	wire _07024_;
	wire _07025_;
	wire _07026_;
	wire _07027_;
	wire _07028_;
	wire _07029_;
	wire _07030_;
	wire _07031_;
	wire _07032_;
	wire _07033_;
	wire _07034_;
	wire _07035_;
	wire _07036_;
	wire _07037_;
	wire _07038_;
	wire _07039_;
	wire _07040_;
	wire _07041_;
	wire _07042_;
	wire _07043_;
	wire _07044_;
	wire _07045_;
	wire _07046_;
	wire _07047_;
	wire _07048_;
	wire _07049_;
	wire _07050_;
	wire _07051_;
	wire _07052_;
	wire _07053_;
	wire _07054_;
	wire _07055_;
	wire _07056_;
	wire _07057_;
	wire _07058_;
	wire _07059_;
	wire _07060_;
	wire _07061_;
	wire _07062_;
	wire _07063_;
	wire _07064_;
	wire _07065_;
	wire _07066_;
	wire _07067_;
	wire _07068_;
	wire _07069_;
	wire _07070_;
	wire _07071_;
	wire _07072_;
	wire _07073_;
	wire _07074_;
	wire _07075_;
	wire _07076_;
	wire _07077_;
	wire _07078_;
	wire _07079_;
	wire _07080_;
	wire _07081_;
	wire _07082_;
	wire _07083_;
	wire _07084_;
	wire _07085_;
	wire _07086_;
	wire _07087_;
	wire _07088_;
	wire _07089_;
	wire _07090_;
	wire _07091_;
	wire _07092_;
	wire _07093_;
	wire _07094_;
	wire _07095_;
	wire _07096_;
	wire _07097_;
	wire _07098_;
	wire _07099_;
	wire _07100_;
	wire _07101_;
	wire _07102_;
	wire _07103_;
	wire _07104_;
	wire _07105_;
	wire _07106_;
	wire _07107_;
	wire _07108_;
	wire _07109_;
	wire _07110_;
	wire _07111_;
	wire _07112_;
	wire _07113_;
	wire _07114_;
	wire _07115_;
	wire _07116_;
	wire _07117_;
	wire _07118_;
	wire _07119_;
	wire _07120_;
	wire _07121_;
	wire _07122_;
	wire _07123_;
	wire _07124_;
	wire _07125_;
	wire _07126_;
	wire _07127_;
	wire _07128_;
	wire _07129_;
	wire _07130_;
	wire _07131_;
	wire _07132_;
	wire _07133_;
	wire _07134_;
	wire _07135_;
	wire _07136_;
	wire _07137_;
	wire _07138_;
	wire _07139_;
	wire _07140_;
	wire _07141_;
	wire _07142_;
	wire _07143_;
	wire _07144_;
	wire _07145_;
	wire _07146_;
	wire _07147_;
	wire _07148_;
	wire _07149_;
	wire _07150_;
	wire _07151_;
	wire _07152_;
	wire _07153_;
	wire _07154_;
	wire _07155_;
	wire _07156_;
	wire _07157_;
	wire _07158_;
	wire _07159_;
	wire _07160_;
	wire _07161_;
	wire _07162_;
	wire _07163_;
	wire _07164_;
	wire _07165_;
	wire _07166_;
	wire _07167_;
	wire _07168_;
	wire _07169_;
	wire _07170_;
	wire _07171_;
	wire _07172_;
	wire _07173_;
	wire _07174_;
	wire _07175_;
	wire _07176_;
	wire _07177_;
	wire _07178_;
	wire _07179_;
	wire _07180_;
	wire _07181_;
	wire _07182_;
	wire _07183_;
	wire _07184_;
	wire _07185_;
	wire _07186_;
	wire _07187_;
	wire _07188_;
	wire _07189_;
	wire _07190_;
	wire _07191_;
	wire _07192_;
	wire _07193_;
	wire _07194_;
	wire _07195_;
	wire _07196_;
	wire _07197_;
	wire _07198_;
	wire _07199_;
	wire _07200_;
	wire _07201_;
	wire _07202_;
	wire _07203_;
	wire _07204_;
	wire _07205_;
	wire _07206_;
	wire _07207_;
	wire _07208_;
	wire _07209_;
	wire _07210_;
	wire _07211_;
	wire _07212_;
	wire _07213_;
	wire _07214_;
	wire _07215_;
	wire _07216_;
	wire _07217_;
	wire _07218_;
	wire _07219_;
	wire _07220_;
	wire _07221_;
	wire _07222_;
	wire _07223_;
	wire _07224_;
	wire _07225_;
	wire _07226_;
	wire _07227_;
	wire _07228_;
	wire _07229_;
	wire _07230_;
	wire _07231_;
	wire _07232_;
	wire _07233_;
	wire _07234_;
	wire _07235_;
	wire _07236_;
	wire _07237_;
	wire _07238_;
	wire _07239_;
	wire _07240_;
	wire _07241_;
	wire _07242_;
	wire _07243_;
	wire _07244_;
	wire _07245_;
	wire _07246_;
	wire _07247_;
	wire _07248_;
	wire _07249_;
	wire _07250_;
	wire _07251_;
	wire _07252_;
	wire _07253_;
	wire _07254_;
	wire _07255_;
	wire _07256_;
	wire _07257_;
	wire _07258_;
	wire _07259_;
	wire _07260_;
	wire _07261_;
	wire _07262_;
	wire _07263_;
	wire _07264_;
	wire _07265_;
	wire _07266_;
	wire _07267_;
	wire _07268_;
	wire _07269_;
	wire _07270_;
	wire _07271_;
	wire _07272_;
	wire _07273_;
	wire _07274_;
	wire _07275_;
	wire _07276_;
	wire _07277_;
	wire _07278_;
	wire _07279_;
	wire _07280_;
	wire _07281_;
	wire _07282_;
	wire _07283_;
	wire _07284_;
	wire _07285_;
	wire _07286_;
	wire _07287_;
	wire _07288_;
	wire _07289_;
	wire _07290_;
	wire _07291_;
	wire _07292_;
	wire _07293_;
	wire _07294_;
	wire _07295_;
	wire _07296_;
	wire _07297_;
	wire _07298_;
	wire _07299_;
	wire _07300_;
	wire _07301_;
	wire _07302_;
	wire _07303_;
	wire _07304_;
	wire _07305_;
	wire _07306_;
	wire _07307_;
	wire _07308_;
	wire _07309_;
	wire _07310_;
	wire _07311_;
	wire _07312_;
	wire _07313_;
	wire _07314_;
	wire _07315_;
	wire _07316_;
	wire _07317_;
	wire _07318_;
	wire _07319_;
	wire _07320_;
	wire _07321_;
	wire _07322_;
	wire _07323_;
	wire _07324_;
	wire _07325_;
	wire _07326_;
	wire _07327_;
	wire _07328_;
	wire _07329_;
	wire _07330_;
	wire _07331_;
	wire _07332_;
	wire _07333_;
	wire _07334_;
	wire _07335_;
	wire _07336_;
	wire _07337_;
	wire _07338_;
	wire _07339_;
	wire _07340_;
	wire _07341_;
	wire _07342_;
	wire _07343_;
	wire _07344_;
	wire _07345_;
	wire _07346_;
	wire _07347_;
	wire _07348_;
	wire _07349_;
	wire _07350_;
	wire _07351_;
	wire _07352_;
	wire _07353_;
	wire _07354_;
	wire _07355_;
	wire _07356_;
	wire _07357_;
	wire _07358_;
	wire _07359_;
	wire _07360_;
	wire _07361_;
	wire _07362_;
	wire _07363_;
	wire _07364_;
	wire _07365_;
	wire _07366_;
	wire _07367_;
	wire _07368_;
	wire _07369_;
	wire _07370_;
	wire _07371_;
	wire _07372_;
	wire _07373_;
	wire _07374_;
	wire _07375_;
	wire _07376_;
	wire _07377_;
	wire _07378_;
	wire _07379_;
	wire _07380_;
	wire _07381_;
	wire _07382_;
	wire _07383_;
	wire _07384_;
	wire _07385_;
	wire _07386_;
	wire _07387_;
	wire _07388_;
	wire _07389_;
	wire _07390_;
	wire _07391_;
	wire _07392_;
	wire _07393_;
	wire _07394_;
	wire _07395_;
	wire _07396_;
	wire _07397_;
	wire _07398_;
	wire _07399_;
	wire _07400_;
	wire _07401_;
	wire _07402_;
	wire _07403_;
	wire _07404_;
	wire _07405_;
	wire _07406_;
	wire _07407_;
	wire _07408_;
	wire _07409_;
	wire _07410_;
	wire _07411_;
	wire _07412_;
	wire _07413_;
	wire _07414_;
	wire _07415_;
	wire _07416_;
	wire _07417_;
	wire _07418_;
	wire _07419_;
	wire _07420_;
	wire _07421_;
	wire _07422_;
	wire _07423_;
	wire _07424_;
	wire _07425_;
	wire _07426_;
	wire _07427_;
	wire _07428_;
	wire _07429_;
	wire _07430_;
	wire _07431_;
	wire _07432_;
	wire _07433_;
	wire _07434_;
	wire _07435_;
	wire _07436_;
	wire _07437_;
	wire _07438_;
	wire _07439_;
	wire _07440_;
	wire _07441_;
	wire _07442_;
	wire _07443_;
	wire _07444_;
	wire _07445_;
	wire _07446_;
	wire _07447_;
	wire _07448_;
	wire _07449_;
	wire _07450_;
	wire _07451_;
	wire _07452_;
	wire _07453_;
	wire _07454_;
	wire _07455_;
	wire _07456_;
	wire _07457_;
	wire _07458_;
	wire _07459_;
	wire _07460_;
	wire _07461_;
	wire _07462_;
	wire _07463_;
	wire _07464_;
	wire _07465_;
	wire _07466_;
	wire _07467_;
	wire _07468_;
	wire _07469_;
	wire _07470_;
	wire _07471_;
	wire _07472_;
	wire _07473_;
	wire _07474_;
	wire _07475_;
	wire _07476_;
	wire _07477_;
	wire _07478_;
	wire _07479_;
	wire _07480_;
	wire _07481_;
	wire _07482_;
	wire _07483_;
	wire _07484_;
	wire _07485_;
	wire _07486_;
	wire _07487_;
	wire _07488_;
	wire _07489_;
	wire _07490_;
	wire _07491_;
	wire _07492_;
	wire _07493_;
	wire _07494_;
	wire _07495_;
	wire _07496_;
	wire _07497_;
	wire _07498_;
	wire _07499_;
	wire _07500_;
	wire _07501_;
	wire _07502_;
	wire _07503_;
	wire _07504_;
	wire _07505_;
	wire _07506_;
	wire _07507_;
	wire _07508_;
	wire _07509_;
	wire _07510_;
	wire _07511_;
	wire _07512_;
	wire _07513_;
	wire _07514_;
	wire _07515_;
	wire _07516_;
	wire _07517_;
	wire _07518_;
	wire _07519_;
	wire _07520_;
	wire _07521_;
	wire _07522_;
	wire _07523_;
	wire _07524_;
	wire _07525_;
	wire _07526_;
	wire _07527_;
	wire _07528_;
	wire _07529_;
	wire _07530_;
	wire _07531_;
	wire _07532_;
	wire _07533_;
	wire _07534_;
	wire _07535_;
	wire _07536_;
	wire _07537_;
	wire _07538_;
	wire _07539_;
	wire _07540_;
	wire _07541_;
	wire _07542_;
	wire _07543_;
	wire _07544_;
	wire _07545_;
	wire _07546_;
	wire _07547_;
	wire _07548_;
	wire _07549_;
	wire _07550_;
	wire _07551_;
	wire _07552_;
	wire _07553_;
	wire _07554_;
	wire _07555_;
	wire _07556_;
	wire _07557_;
	wire _07558_;
	wire _07559_;
	wire _07560_;
	wire _07561_;
	wire _07562_;
	wire _07563_;
	wire _07564_;
	wire _07565_;
	wire _07566_;
	wire _07567_;
	wire _07568_;
	wire _07569_;
	wire _07570_;
	wire _07571_;
	wire _07572_;
	wire _07573_;
	wire _07574_;
	wire _07575_;
	wire _07576_;
	wire _07577_;
	wire _07578_;
	wire _07579_;
	wire _07580_;
	wire _07581_;
	wire _07582_;
	wire _07583_;
	wire _07584_;
	wire _07585_;
	wire _07586_;
	wire _07587_;
	wire _07588_;
	wire _07589_;
	wire _07590_;
	wire _07591_;
	wire _07592_;
	wire _07593_;
	wire _07594_;
	wire _07595_;
	wire _07596_;
	wire _07597_;
	wire _07598_;
	wire _07599_;
	wire _07600_;
	wire _07601_;
	wire _07602_;
	wire _07603_;
	wire _07604_;
	wire _07605_;
	wire _07606_;
	wire _07607_;
	wire _07608_;
	wire _07609_;
	wire _07610_;
	wire _07611_;
	wire _07612_;
	wire _07613_;
	wire _07614_;
	wire _07615_;
	wire _07616_;
	wire _07617_;
	wire _07618_;
	wire _07619_;
	wire _07620_;
	wire _07621_;
	wire _07622_;
	wire _07623_;
	wire _07624_;
	wire _07625_;
	wire _07626_;
	wire _07627_;
	wire _07628_;
	wire _07629_;
	wire _07630_;
	wire _07631_;
	wire _07632_;
	wire _07633_;
	wire _07634_;
	wire _07635_;
	wire _07636_;
	wire _07637_;
	wire _07638_;
	wire _07639_;
	wire _07640_;
	wire _07641_;
	wire _07642_;
	wire _07643_;
	wire _07644_;
	wire _07645_;
	wire _07646_;
	wire _07647_;
	wire _07648_;
	wire _07649_;
	wire _07650_;
	wire _07651_;
	wire _07652_;
	wire _07653_;
	wire _07654_;
	wire _07655_;
	wire _07656_;
	wire _07657_;
	wire _07658_;
	wire _07659_;
	wire _07660_;
	wire _07661_;
	wire _07662_;
	wire _07663_;
	wire _07664_;
	wire _07665_;
	wire _07666_;
	wire _07667_;
	wire _07668_;
	wire _07669_;
	wire _07670_;
	wire _07671_;
	wire _07672_;
	wire _07673_;
	wire _07674_;
	wire _07675_;
	wire _07676_;
	wire _07677_;
	wire _07678_;
	wire _07679_;
	wire _07680_;
	wire _07681_;
	wire _07682_;
	wire _07683_;
	wire _07684_;
	wire _07685_;
	wire _07686_;
	wire _07687_;
	wire _07688_;
	wire _07689_;
	wire _07690_;
	wire _07691_;
	wire _07692_;
	wire _07693_;
	wire _07694_;
	wire _07695_;
	wire _07696_;
	wire _07697_;
	wire _07698_;
	wire _07699_;
	wire _07700_;
	wire _07701_;
	wire _07702_;
	wire _07703_;
	wire _07704_;
	wire _07705_;
	wire _07706_;
	wire _07707_;
	wire _07708_;
	wire _07709_;
	wire _07710_;
	wire _07711_;
	wire _07712_;
	wire _07713_;
	wire _07714_;
	wire _07715_;
	wire _07716_;
	wire _07717_;
	wire _07718_;
	wire _07719_;
	wire _07720_;
	wire _07721_;
	wire _07722_;
	wire _07723_;
	wire _07724_;
	wire _07725_;
	wire _07726_;
	wire _07727_;
	wire _07728_;
	wire _07729_;
	wire _07730_;
	wire _07731_;
	wire _07732_;
	wire _07733_;
	wire _07734_;
	wire _07735_;
	wire _07736_;
	wire _07737_;
	wire _07738_;
	wire _07739_;
	wire _07740_;
	wire _07741_;
	wire _07742_;
	wire _07743_;
	wire _07744_;
	wire _07745_;
	wire _07746_;
	wire _07747_;
	wire _07748_;
	wire _07749_;
	wire _07750_;
	wire _07751_;
	wire _07752_;
	wire _07753_;
	wire _07754_;
	wire _07755_;
	wire _07756_;
	wire _07757_;
	wire _07758_;
	wire _07759_;
	wire _07760_;
	wire _07761_;
	wire _07762_;
	wire _07763_;
	wire _07764_;
	wire _07765_;
	wire _07766_;
	wire _07767_;
	wire _07768_;
	wire _07769_;
	wire _07770_;
	wire _07771_;
	wire _07772_;
	wire _07773_;
	wire _07774_;
	wire _07775_;
	wire _07776_;
	wire _07777_;
	wire _07778_;
	wire _07779_;
	wire _07780_;
	wire _07781_;
	wire _07782_;
	wire _07783_;
	wire _07784_;
	wire _07785_;
	wire _07786_;
	wire _07787_;
	wire _07788_;
	wire _07789_;
	wire _07790_;
	wire _07791_;
	wire _07792_;
	wire _07793_;
	wire _07794_;
	wire _07795_;
	wire _07796_;
	wire _07797_;
	wire _07798_;
	wire _07799_;
	wire _07800_;
	wire _07801_;
	wire _07802_;
	wire _07803_;
	wire _07804_;
	wire _07805_;
	wire _07806_;
	wire _07807_;
	wire _07808_;
	wire _07809_;
	wire _07810_;
	wire _07811_;
	wire _07812_;
	wire _07813_;
	wire _07814_;
	wire _07815_;
	wire _07816_;
	wire _07817_;
	wire _07818_;
	wire _07819_;
	wire _07820_;
	wire _07821_;
	wire _07822_;
	wire _07823_;
	wire _07824_;
	wire _07825_;
	wire _07826_;
	wire _07827_;
	wire _07828_;
	wire _07829_;
	wire _07830_;
	wire _07831_;
	wire _07832_;
	wire _07833_;
	wire _07834_;
	wire _07835_;
	wire _07836_;
	wire _07837_;
	wire _07838_;
	wire _07839_;
	wire _07840_;
	wire _07841_;
	wire _07842_;
	wire _07843_;
	wire _07844_;
	wire _07845_;
	wire _07846_;
	wire _07847_;
	wire _07848_;
	wire _07849_;
	wire _07850_;
	wire _07851_;
	wire _07852_;
	wire _07853_;
	wire _07854_;
	wire _07855_;
	wire _07856_;
	wire _07857_;
	wire _07858_;
	wire _07859_;
	wire _07860_;
	wire _07861_;
	wire _07862_;
	wire _07863_;
	wire _07864_;
	wire _07865_;
	wire _07866_;
	wire _07867_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	reg [11:0] \mchip.index ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire [7:0] \mchip.val ;
	assign _01098_ = ~\mchip.index [4];
	assign _01209_ = ~(\mchip.index [2] & \mchip.index [0]);
	assign _01320_ = _01209_ | \mchip.index [3];
	assign _01431_ = _01320_ | _01098_;
	assign _01542_ = _01431_ | \mchip.index [7];
	assign _01653_ = _01542_ | \mchip.index [9];
	assign _01764_ = \mchip.index [10] & ~_01653_;
	assign _01875_ = ~\mchip.index [11];
	assign _01986_ = ~\mchip.index [10];
	assign _02097_ = ~\mchip.index [7];
	assign _02208_ = ~\mchip.index [2];
	assign _02319_ = \mchip.index [1] | ~\mchip.index [0];
	assign _02430_ = _02319_ | _02208_;
	assign _02540_ = _02430_ | \mchip.index [4];
	assign _02651_ = _02540_ | _02097_;
	assign _02762_ = _02651_ | _01986_;
	assign _02873_ = _01875_ & ~_02762_;
	assign _02984_ = ~\mchip.index [6];
	assign _03095_ = ~(\mchip.index [0] & \mchip.index [5]);
	assign _03206_ = _03095_ | _02984_;
	assign _03317_ = _03206_ | _02097_;
	assign _03428_ = _03317_ | \mchip.index [8];
	assign _03539_ = \mchip.index [10] & ~_03428_;
	assign _03650_ = \mchip.index [0] | ~\mchip.index [2];
	assign _03761_ = _03650_ | \mchip.index [6];
	assign _03871_ = _03761_ | _02097_;
	assign _03982_ = _03871_ | \mchip.index [9];
	assign _04093_ = \mchip.index [10] & ~_03982_;
	assign _04204_ = _02319_ | _01098_;
	assign _04315_ = _04204_ | _02097_;
	assign _04426_ = _04315_ | \mchip.index [8];
	assign _04537_ = \mchip.index [10] & ~_04426_;
	assign _04648_ = ~\mchip.index [8];
	assign _04759_ = \mchip.index [1] | ~\mchip.index [2];
	assign _04870_ = _04759_ | \mchip.index [4];
	assign _04981_ = _04870_ | \mchip.index [5];
	assign _05091_ = _04981_ | \mchip.index [6];
	assign _05202_ = _05091_ | _04648_;
	assign _05313_ = \mchip.index [11] & ~_05202_;
	assign _05424_ = ~\mchip.index [5];
	assign _05535_ = _04870_ | _05424_;
	assign _05646_ = _05535_ | \mchip.index [7];
	assign _05757_ = \mchip.index [11] & ~_05646_;
	assign _05868_ = \mchip.index [0] | ~\mchip.index [1];
	assign _05979_ = _05868_ | \mchip.index [3];
	assign _06090_ = _05979_ | _01098_;
	assign _06201_ = _06090_ | \mchip.index [8];
	assign _06312_ = _06201_ | \mchip.index [9];
	assign _06422_ = _01875_ & ~_06312_;
	assign _06533_ = _04759_ | \mchip.index [6];
	assign _06644_ = _06533_ | _04648_;
	assign _06755_ = _06644_ | \mchip.index [9];
	assign _06866_ = \mchip.index [10] & ~_06755_;
	assign _06977_ = ~(\mchip.index [1] & \mchip.index [0]);
	assign _07088_ = _06977_ | \mchip.index [2];
	assign _07199_ = _07088_ | \mchip.index [3];
	assign _07310_ = _07199_ | \mchip.index [4];
	assign _07421_ = _07310_ | \mchip.index [7];
	assign _07532_ = _04648_ & ~_07421_;
	assign _07637_ = \mchip.index [2] | ~\mchip.index [0];
	assign _07648_ = _07637_ | \mchip.index [3];
	assign _07659_ = _07648_ | _02984_;
	assign _07670_ = _07659_ | \mchip.index [7];
	assign _07681_ = _07670_ | \mchip.index [8];
	assign _07692_ = \mchip.index [9] & ~_07681_;
	assign _07703_ = ~(\mchip.index [2] & \mchip.index [1]);
	assign _07714_ = _07703_ | \mchip.index [3];
	assign _07725_ = _07714_ | _01098_;
	assign _07736_ = _07725_ | \mchip.index [7];
	assign _07747_ = \mchip.index [11] & ~_07736_;
	assign _07758_ = ~\mchip.index [9];
	assign _07769_ = ~(\mchip.index [3] & \mchip.index [2]);
	assign _07780_ = _07769_ | _01098_;
	assign _07791_ = _07780_ | \mchip.index [8];
	assign _07802_ = _07791_ | _07758_;
	assign _07813_ = \mchip.index [10] & ~_07802_;
	assign _07824_ = _07703_ | _01098_;
	assign _07835_ = _07824_ | \mchip.index [6];
	assign _07846_ = _07835_ | \mchip.index [8];
	assign _07857_ = _07758_ & ~_07846_;
	assign _00000_ = _05868_ | \mchip.index [2];
	assign _00011_ = _00000_ | \mchip.index [5];
	assign _00022_ = _00011_ | \mchip.index [6];
	assign _00033_ = _00022_ | _02097_;
	assign _00044_ = \mchip.index [9] & ~_00033_;
	assign _00055_ = _02319_ | \mchip.index [4];
	assign _00066_ = _00055_ | \mchip.index [6];
	assign _00077_ = _00066_ | _04648_;
	assign _00088_ = \mchip.index [11] & ~_00077_;
	assign _00099_ = ~(\mchip.index [3] & \mchip.index [1]);
	assign _00110_ = _00099_ | _01098_;
	assign _00121_ = _00110_ | _04648_;
	assign _00132_ = _00121_ | \mchip.index [10];
	assign _00143_ = \mchip.index [11] & ~_00132_;
	assign _00154_ = _01320_ | \mchip.index [4];
	assign _00165_ = _00154_ | _04648_;
	assign _00176_ = _00165_ | \mchip.index [10];
	assign _00187_ = \mchip.index [11] & ~_00176_;
	assign _00198_ = ~\mchip.index [3];
	assign _00209_ = _06977_ | _00198_;
	assign _00220_ = _00209_ | _02984_;
	assign _00231_ = _00220_ | _02097_;
	assign _00242_ = _00231_ | _04648_;
	assign _00252_ = _01986_ & ~_00242_;
	assign _00263_ = \mchip.index [0] | ~\mchip.index [3];
	assign _00274_ = _00263_ | \mchip.index [7];
	assign _00285_ = _00274_ | \mchip.index [8];
	assign _00296_ = _00285_ | _07758_;
	assign _00307_ = \mchip.index [10] & ~_00296_;
	assign _00318_ = \mchip.index [2] | \mchip.index [0];
	assign _00329_ = _00318_ | \mchip.index [3];
	assign _00340_ = _00329_ | \mchip.index [5];
	assign _00351_ = _00340_ | \mchip.index [6];
	assign _00362_ = _00351_ | _01986_;
	assign _00373_ = _01875_ & ~_00362_;
	assign _00384_ = _07637_ | _00198_;
	assign _00395_ = _00384_ | _01098_;
	assign _00406_ = _00395_ | _02984_;
	assign _00417_ = _00406_ | \mchip.index [7];
	assign _00428_ = _00417_ | _04648_;
	assign _00439_ = \mchip.index [9] & ~_00428_;
	assign _00450_ = _02319_ | \mchip.index [3];
	assign _00461_ = _00450_ | \mchip.index [4];
	assign _00472_ = _00461_ | \mchip.index [5];
	assign _00483_ = _00472_ | _02097_;
	assign _00494_ = \mchip.index [9] & ~_00483_;
	assign _00505_ = _03650_ | _00198_;
	assign _00516_ = _00505_ | _01098_;
	assign _00527_ = _00516_ | \mchip.index [6];
	assign _00538_ = _00527_ | _04648_;
	assign _00549_ = _01875_ & ~_00538_;
	assign _00560_ = \mchip.index [1] | \mchip.index [0];
	assign _00571_ = _00560_ | _00198_;
	assign _00582_ = _00571_ | _01098_;
	assign _00593_ = _00582_ | \mchip.index [6];
	assign _00604_ = _00593_ | \mchip.index [8];
	assign _00615_ = \mchip.index [9] & ~_00604_;
	assign _00626_ = _00384_ | _02984_;
	assign _00637_ = _00626_ | _02097_;
	assign _00648_ = _00637_ | _04648_;
	assign _00659_ = _01986_ & ~_00648_;
	assign _00670_ = _00000_ | \mchip.index [3];
	assign _00681_ = _00670_ | \mchip.index [5];
	assign _00692_ = _00681_ | _02984_;
	assign _00703_ = _00692_ | _02097_;
	assign _00714_ = _01875_ & ~_00703_;
	assign _00725_ = \mchip.index [1] | ~\mchip.index [5];
	assign _00736_ = _00725_ | \mchip.index [7];
	assign _00747_ = _00736_ | _04648_;
	assign _00758_ = _00747_ | _07758_;
	assign _00769_ = _01875_ & ~_00758_;
	assign _00780_ = \mchip.index [3] | \mchip.index [0];
	assign _00791_ = _00780_ | _01098_;
	assign _00802_ = _00791_ | _05424_;
	assign _00813_ = _02097_ & ~_00802_;
	assign _00824_ = _07703_ | _00198_;
	assign _00835_ = _00824_ | \mchip.index [4];
	assign _00846_ = _00835_ | _02097_;
	assign _00857_ = _00846_ | _07758_;
	assign _00868_ = _01986_ & ~_00857_;
	assign _00879_ = _01209_ | _00198_;
	assign _00890_ = _00879_ | _02097_;
	assign _00901_ = _00890_ | \mchip.index [8];
	assign _00912_ = \mchip.index [11] & ~_00901_;
	assign _00923_ = _00560_ | \mchip.index [2];
	assign _00934_ = _00923_ | \mchip.index [4];
	assign _00945_ = _00934_ | \mchip.index [5];
	assign _00956_ = _00945_ | _04648_;
	assign _00967_ = _00956_ | \mchip.index [10];
	assign _00978_ = _01875_ & ~_00967_;
	assign _00989_ = _04759_ | _00198_;
	assign _01000_ = _00989_ | \mchip.index [4];
	assign _01011_ = _01000_ | \mchip.index [7];
	assign _01022_ = _01011_ | _07758_;
	assign _01033_ = _01875_ & ~_01022_;
	assign _01044_ = _07637_ | \mchip.index [4];
	assign _01055_ = _01044_ | \mchip.index [6];
	assign _01066_ = _01055_ | \mchip.index [7];
	assign _01077_ = _01066_ | _04648_;
	assign _01088_ = \mchip.index [10] & ~_01077_;
	assign _01099_ = _00923_ | \mchip.index [3];
	assign _01110_ = _01099_ | _05424_;
	assign _01121_ = _01110_ | _02097_;
	assign _01132_ = _01875_ & ~_01121_;
	assign _01143_ = _00571_ | \mchip.index [5];
	assign _01154_ = _01143_ | _04648_;
	assign _01165_ = _01154_ | \mchip.index [9];
	assign _01176_ = \mchip.index [10] & ~_01165_;
	assign _01187_ = _07824_ | _02984_;
	assign _01198_ = _01187_ | \mchip.index [7];
	assign _01210_ = _01198_ | _07758_;
	assign _01221_ = \mchip.index [11] & ~_01210_;
	assign _01232_ = ~(\mchip.index [4] & \mchip.index [2]);
	assign _01243_ = _01232_ | \mchip.index [6];
	assign _01254_ = _01243_ | _02097_;
	assign _01265_ = _01254_ | _04648_;
	assign _01276_ = _01265_ | \mchip.index [10];
	assign _01287_ = _01875_ & ~_01276_;
	assign _01298_ = _00450_ | _02984_;
	assign _01309_ = _01298_ | _02097_;
	assign _01321_ = _01309_ | \mchip.index [9];
	assign _01332_ = \mchip.index [11] & ~_01321_;
	assign _01343_ = _02430_ | _01098_;
	assign _01354_ = _01343_ | \mchip.index [7];
	assign _01365_ = _01875_ & ~_01354_;
	assign _01376_ = _02430_ | \mchip.index [3];
	assign _01387_ = _01376_ | _01098_;
	assign _01398_ = _01387_ | \mchip.index [5];
	assign _01409_ = _01398_ | \mchip.index [7];
	assign _01420_ = \mchip.index [8] & ~_01409_;
	assign _01432_ = _01209_ | \mchip.index [6];
	assign _01443_ = _01432_ | _02097_;
	assign _01454_ = _01443_ | _01986_;
	assign _01465_ = \mchip.index [11] & ~_01454_;
	assign _01476_ = _00670_ | \mchip.index [4];
	assign _01487_ = _01476_ | \mchip.index [9];
	assign _01498_ = \mchip.index [11] & ~_01487_;
	assign _01509_ = \mchip.index [2] | ~\mchip.index [4];
	assign _01520_ = _01509_ | _02097_;
	assign _01531_ = _01520_ | _04648_;
	assign _01543_ = _01531_ | \mchip.index [9];
	assign _01554_ = \mchip.index [11] & ~_01543_;
	assign _01565_ = _05979_ | \mchip.index [5];
	assign _01576_ = _01565_ | \mchip.index [6];
	assign _01587_ = _01576_ | _02097_;
	assign _01598_ = _01587_ | _07758_;
	assign _01609_ = _01875_ & ~_01598_;
	assign _01620_ = \mchip.index [2] | ~\mchip.index [1];
	assign _01631_ = _01620_ | \mchip.index [4];
	assign _01642_ = _01631_ | \mchip.index [5];
	assign _01654_ = _01642_ | \mchip.index [6];
	assign _01665_ = _01654_ | \mchip.index [7];
	assign _01676_ = \mchip.index [11] & ~_01665_;
	assign _01687_ = _07637_ | _01098_;
	assign _01698_ = _01687_ | \mchip.index [8];
	assign _01709_ = _01698_ | _07758_;
	assign _01720_ = \mchip.index [11] & ~_01709_;
	assign _01731_ = _00000_ | \mchip.index [4];
	assign _01742_ = _01731_ | \mchip.index [5];
	assign _01753_ = _01742_ | \mchip.index [7];
	assign _01765_ = _04648_ & ~_01753_;
	assign _01776_ = _03650_ | \mchip.index [3];
	assign _01787_ = _01776_ | \mchip.index [6];
	assign _01798_ = _01787_ | \mchip.index [8];
	assign _01809_ = _01798_ | \mchip.index [9];
	assign _01820_ = \mchip.index [11] & ~_01809_;
	assign _01831_ = \mchip.index [1] | ~\mchip.index [3];
	assign _01842_ = _01831_ | \mchip.index [4];
	assign _01853_ = _01842_ | \mchip.index [8];
	assign _01864_ = _01853_ | \mchip.index [9];
	assign _01876_ = _01864_ | \mchip.index [10];
	assign _01887_ = _01875_ & ~_01876_;
	assign _01898_ = _07769_ | \mchip.index [5];
	assign _01909_ = _01898_ | \mchip.index [6];
	assign _01920_ = _01909_ | _02097_;
	assign _01931_ = _01920_ | \mchip.index [8];
	assign _01942_ = \mchip.index [10] & ~_01931_;
	assign _01953_ = \mchip.index [2] | \mchip.index [1];
	assign _01964_ = _01953_ | \mchip.index [3];
	assign _01975_ = _01964_ | \mchip.index [5];
	assign _01987_ = _01975_ | \mchip.index [6];
	assign _01998_ = _01987_ | _04648_;
	assign _02009_ = _01998_ | \mchip.index [9];
	assign _02020_ = _01986_ & ~_02009_;
	assign _02031_ = _01776_ | _05424_;
	assign _02042_ = _02031_ | _02984_;
	assign _02053_ = \mchip.index [10] & ~_02042_;
	assign _02064_ = _05979_ | \mchip.index [6];
	assign _02075_ = _02064_ | \mchip.index [7];
	assign _02086_ = _02075_ | _07758_;
	assign _02098_ = \mchip.index [11] & ~_02086_;
	assign _02109_ = _00450_ | \mchip.index [5];
	assign _02120_ = _02109_ | \mchip.index [8];
	assign _02131_ = _02120_ | \mchip.index [9];
	assign _02142_ = \mchip.index [10] & ~_02131_;
	assign _02153_ = _05868_ | _00198_;
	assign _02164_ = _02153_ | \mchip.index [5];
	assign _02175_ = _02164_ | \mchip.index [6];
	assign _02186_ = _02175_ | \mchip.index [8];
	assign _02197_ = \mchip.index [10] & ~_02186_;
	assign _02209_ = _00000_ | _01098_;
	assign _02220_ = _02209_ | _02984_;
	assign _02231_ = _02220_ | _02097_;
	assign _02242_ = _07758_ & ~_02231_;
	assign _02253_ = ~(\mchip.index [3] & \mchip.index [0]);
	assign _02264_ = _02253_ | _01098_;
	assign _02275_ = _02264_ | _02097_;
	assign _02286_ = _02275_ | _07758_;
	assign _02297_ = _02286_ | _01986_;
	assign _02308_ = _01875_ & ~_02297_;
	assign _02320_ = _00923_ | _00198_;
	assign _02331_ = _02320_ | \mchip.index [8];
	assign _02342_ = _02331_ | \mchip.index [9];
	assign _02353_ = _01986_ & ~_02342_;
	assign _02364_ = _00989_ | _01098_;
	assign _02375_ = _02364_ | \mchip.index [6];
	assign _02386_ = _02375_ | _02097_;
	assign _02397_ = \mchip.index [9] & ~_02386_;
	assign _02408_ = _05868_ | _02208_;
	assign _02419_ = _02408_ | _01098_;
	assign _02431_ = _02419_ | _02984_;
	assign _02441_ = _02431_ | \mchip.index [7];
	assign _02452_ = _01875_ & ~_02441_;
	assign _02463_ = ~(\mchip.index [4] & \mchip.index [1]);
	assign _02474_ = _02463_ | _02984_;
	assign _02485_ = _02474_ | \mchip.index [8];
	assign _02496_ = _02485_ | _07758_;
	assign _02507_ = _01986_ & ~_02496_;
	assign _02518_ = _01776_ | \mchip.index [5];
	assign _02529_ = _02518_ | _02984_;
	assign _02541_ = _02529_ | \mchip.index [9];
	assign _02552_ = _02541_ | \mchip.index [10];
	assign _02563_ = _01875_ & ~_02552_;
	assign _02574_ = _04870_ | \mchip.index [6];
	assign _02585_ = _02574_ | _02097_;
	assign _02596_ = _02585_ | \mchip.index [8];
	assign _02607_ = _01875_ & ~_02596_;
	assign _02618_ = \mchip.index [3] | \mchip.index [1];
	assign _02629_ = _02618_ | \mchip.index [4];
	assign _02640_ = _02629_ | _02097_;
	assign _02652_ = _02640_ | \mchip.index [8];
	assign _02663_ = _02652_ | _07758_;
	assign _02674_ = _01986_ & ~_02663_;
	assign _02685_ = _02319_ | \mchip.index [2];
	assign _02696_ = _02685_ | \mchip.index [3];
	assign _02707_ = _02696_ | _01098_;
	assign _02718_ = _02707_ | _02984_;
	assign _02729_ = _04648_ & ~_02718_;
	assign _02740_ = _07637_ | _02984_;
	assign _02751_ = _02740_ | _02097_;
	assign _02763_ = _02751_ | \mchip.index [8];
	assign _02774_ = _02763_ | \mchip.index [9];
	assign _02785_ = \mchip.index [10] & ~_02774_;
	assign _02796_ = _01509_ | _02984_;
	assign _02807_ = _02796_ | _04648_;
	assign _02818_ = _02807_ | _07758_;
	assign _02829_ = _01986_ & ~_02818_;
	assign _02840_ = _00384_ | \mchip.index [4];
	assign _02851_ = _02840_ | \mchip.index [6];
	assign _02862_ = _02851_ | \mchip.index [7];
	assign _02874_ = \mchip.index [10] & ~_02862_;
	assign _02885_ = _00055_ | \mchip.index [5];
	assign _02896_ = _02885_ | _02984_;
	assign _02907_ = _02896_ | \mchip.index [8];
	assign _02918_ = \mchip.index [10] & ~_02907_;
	assign _02929_ = \mchip.index [2] | \mchip.index [5];
	assign _02940_ = _02929_ | _02984_;
	assign _02951_ = _02940_ | _02097_;
	assign _02962_ = _02951_ | _04648_;
	assign _02973_ = _02962_ | _07758_;
	assign _02985_ = _01875_ & ~_02973_;
	assign _02996_ = _00582_ | _02984_;
	assign _03007_ = _02996_ | _01986_;
	assign _03018_ = _01875_ & ~_03007_;
	assign _03029_ = _00450_ | _01098_;
	assign _03040_ = _03029_ | _02984_;
	assign _03051_ = _03040_ | \mchip.index [7];
	assign _03062_ = _03051_ | _01986_;
	assign _03073_ = _01875_ & ~_03062_;
	assign _03084_ = _01209_ | \mchip.index [4];
	assign _03096_ = _03084_ | \mchip.index [5];
	assign _03107_ = _03096_ | \mchip.index [6];
	assign _03118_ = _03107_ | _02097_;
	assign _03129_ = _03118_ | _04648_;
	assign _03140_ = _07758_ & ~_03129_;
	assign _03151_ = _07703_ | _02984_;
	assign _03162_ = _03151_ | _02097_;
	assign _03173_ = _03162_ | \mchip.index [8];
	assign _03184_ = _03173_ | \mchip.index [10];
	assign _03195_ = _01875_ & ~_03184_;
	assign _03207_ = _01432_ | \mchip.index [7];
	assign _03218_ = _03207_ | _07758_;
	assign _03229_ = _01875_ & ~_03218_;
	assign _03240_ = _02320_ | \mchip.index [4];
	assign _03251_ = _03240_ | _02097_;
	assign _03262_ = _01986_ & ~_03251_;
	assign _03273_ = _07725_ | _02097_;
	assign _03284_ = _03273_ | \mchip.index [10];
	assign _03295_ = _01875_ & ~_03284_;
	assign _03306_ = _02319_ | \mchip.index [5];
	assign _03318_ = _03306_ | _02984_;
	assign _03329_ = _03318_ | \mchip.index [8];
	assign _03340_ = _03329_ | \mchip.index [9];
	assign _03351_ = \mchip.index [10] & ~_03340_;
	assign _03362_ = _02209_ | _04648_;
	assign _03373_ = _03362_ | _07758_;
	assign _03384_ = _01875_ & ~_03373_;
	assign _03395_ = _01620_ | _00198_;
	assign _03406_ = _03395_ | _01098_;
	assign _03417_ = _03406_ | _02097_;
	assign _03429_ = _03417_ | \mchip.index [8];
	assign _03440_ = _01986_ & ~_03429_;
	assign _03451_ = _00505_ | _02984_;
	assign _03462_ = _03451_ | \mchip.index [7];
	assign _03473_ = _03462_ | _07758_;
	assign _03484_ = _03473_ | _01986_;
	assign _03495_ = _01875_ & ~_03484_;
	assign _03506_ = _02109_ | _02097_;
	assign _03517_ = _03506_ | _04648_;
	assign _03528_ = _01986_ & ~_03517_;
	assign _03540_ = _06977_ | \mchip.index [4];
	assign _03551_ = _03540_ | \mchip.index [7];
	assign _03562_ = _03551_ | \mchip.index [8];
	assign _03573_ = _03562_ | \mchip.index [9];
	assign _03584_ = _01986_ & ~_03573_;
	assign _03595_ = _06533_ | \mchip.index [7];
	assign _03606_ = _03595_ | _07758_;
	assign _03617_ = _01875_ & ~_03606_;
	assign _03628_ = _00560_ | _05424_;
	assign _03639_ = _03628_ | \mchip.index [6];
	assign _03651_ = _03639_ | _02097_;
	assign _03662_ = _01875_ & ~_03651_;
	assign _03673_ = _02419_ | _04648_;
	assign _03684_ = _03673_ | \mchip.index [9];
	assign _03695_ = _01986_ & ~_03684_;
	assign _03706_ = _02696_ | _02097_;
	assign _03717_ = _03706_ | \mchip.index [8];
	assign _03728_ = \mchip.index [9] & ~_03717_;
	assign _03739_ = _00450_ | \mchip.index [6];
	assign _03750_ = _03739_ | \mchip.index [7];
	assign _03762_ = _03750_ | _04648_;
	assign _03772_ = \mchip.index [11] & ~_03762_;
	assign _03783_ = \mchip.index [4] | \mchip.index [2];
	assign _03794_ = _03783_ | \mchip.index [5];
	assign _03805_ = _03794_ | \mchip.index [6];
	assign _03816_ = _03805_ | _04648_;
	assign _03827_ = _03816_ | _07758_;
	assign _03838_ = _03827_ | _01986_;
	assign _03849_ = \mchip.index [11] & ~_03838_;
	assign _03860_ = _01831_ | _01098_;
	assign _03872_ = _03860_ | \mchip.index [7];
	assign _03883_ = _03872_ | \mchip.index [8];
	assign _03894_ = _03883_ | \mchip.index [9];
	assign _03905_ = \mchip.index [11] & ~_03894_;
	assign _03916_ = _06977_ | _05424_;
	assign _03927_ = _03916_ | _02984_;
	assign _03938_ = _03927_ | _04648_;
	assign _03949_ = \mchip.index [11] & ~_03938_;
	assign _03960_ = _03650_ | \mchip.index [4];
	assign _03971_ = _03960_ | \mchip.index [5];
	assign _03983_ = _03971_ | _02984_;
	assign _03994_ = _03983_ | _02097_;
	assign _04005_ = _03994_ | \mchip.index [8];
	assign _04016_ = _07758_ & ~_04005_;
	assign _04027_ = _02796_ | _02097_;
	assign _04038_ = _04027_ | \mchip.index [9];
	assign _04049_ = \mchip.index [11] & ~_04038_;
	assign _04060_ = _02209_ | \mchip.index [5];
	assign _04071_ = _04060_ | \mchip.index [6];
	assign _04082_ = _04071_ | _07758_;
	assign _04094_ = \mchip.index [10] & ~_04082_;
	assign _04105_ = _01232_ | _02984_;
	assign _04116_ = _04105_ | \mchip.index [7];
	assign _04127_ = _04116_ | \mchip.index [8];
	assign _04138_ = \mchip.index [9] & ~_04127_;
	assign _04149_ = _02153_ | \mchip.index [6];
	assign _04160_ = _04149_ | _02097_;
	assign _04171_ = _04160_ | _04648_;
	assign _04182_ = \mchip.index [9] & ~_04171_;
	assign _04193_ = _00560_ | \mchip.index [3];
	assign _04205_ = _04193_ | \mchip.index [4];
	assign _04216_ = _04205_ | \mchip.index [7];
	assign _04227_ = _04216_ | _01986_;
	assign _04238_ = _01875_ & ~_04227_;
	assign _04249_ = \mchip.index [2] | ~\mchip.index [3];
	assign _04260_ = _04249_ | \mchip.index [4];
	assign _04271_ = _04260_ | _02984_;
	assign _04282_ = _04271_ | _02097_;
	assign _04293_ = \mchip.index [8] & ~_04282_;
	assign _04304_ = _02629_ | _05424_;
	assign _04316_ = _04304_ | \mchip.index [6];
	assign _04327_ = _04316_ | _02097_;
	assign _04338_ = \mchip.index [10] & ~_04327_;
	assign _04349_ = _02320_ | _02097_;
	assign _04360_ = _04349_ | \mchip.index [8];
	assign _04371_ = _01986_ & ~_04360_;
	assign _04382_ = \mchip.index [3] | ~\mchip.index [1];
	assign _04393_ = _04382_ | \mchip.index [5];
	assign _04404_ = _04393_ | \mchip.index [6];
	assign _04415_ = _04404_ | \mchip.index [7];
	assign _04427_ = _04415_ | \mchip.index [10];
	assign _04438_ = \mchip.index [11] & ~_04427_;
	assign _04449_ = _00516_ | _02984_;
	assign _04460_ = _04449_ | \mchip.index [7];
	assign _04471_ = \mchip.index [10] & ~_04460_;
	assign _04482_ = _03650_ | _01098_;
	assign _04493_ = _04482_ | \mchip.index [5];
	assign _04504_ = _04493_ | \mchip.index [6];
	assign _04515_ = _04504_ | _02097_;
	assign _04526_ = _04515_ | _04648_;
	assign _04538_ = \mchip.index [9] & ~_04526_;
	assign _04549_ = _01000_ | _02097_;
	assign _04560_ = _04549_ | \mchip.index [9];
	assign _04571_ = _01875_ & ~_04560_;
	assign _04582_ = _01044_ | _02984_;
	assign _04593_ = _04582_ | \mchip.index [7];
	assign _04604_ = _04593_ | \mchip.index [10];
	assign _04615_ = \mchip.index [11] & ~_04604_;
	assign _04626_ = _00780_ | _05424_;
	assign _04637_ = _04626_ | _02984_;
	assign _04649_ = _04637_ | _04648_;
	assign _04660_ = _04649_ | _07758_;
	assign _04671_ = _01875_ & ~_04660_;
	assign _04682_ = _00099_ | \mchip.index [4];
	assign _04693_ = _04682_ | \mchip.index [7];
	assign _04704_ = _04693_ | \mchip.index [9];
	assign _04715_ = _04704_ | \mchip.index [10];
	assign _04726_ = _01875_ & ~_04715_;
	assign _04737_ = _02109_ | \mchip.index [6];
	assign _04748_ = _04737_ | _02097_;
	assign _04760_ = \mchip.index [11] & ~_04748_;
	assign _04771_ = _00318_ | \mchip.index [4];
	assign _04782_ = _04771_ | \mchip.index [5];
	assign _04793_ = _04782_ | _02097_;
	assign _04804_ = _04793_ | _04648_;
	assign _04815_ = _04804_ | _07758_;
	assign _04826_ = \mchip.index [10] & ~_04815_;
	assign _04837_ = _07780_ | \mchip.index [6];
	assign _04848_ = _04837_ | _02097_;
	assign _04859_ = \mchip.index [10] & ~_04848_;
	assign _04871_ = _07088_ | _00198_;
	assign _04882_ = _04871_ | _01098_;
	assign _04893_ = _04882_ | _02984_;
	assign _04904_ = _04893_ | \mchip.index [8];
	assign _04915_ = _01875_ & ~_04904_;
	assign _04926_ = _00670_ | \mchip.index [6];
	assign _04937_ = _04926_ | \mchip.index [7];
	assign _04948_ = \mchip.index [8] & ~_04937_;
	assign _04959_ = _00472_ | _02984_;
	assign _04970_ = _04959_ | \mchip.index [8];
	assign _04982_ = \mchip.index [9] & ~_04970_;
	assign _04993_ = _00560_ | _02208_;
	assign _05004_ = _04993_ | \mchip.index [3];
	assign _05015_ = _05004_ | _02984_;
	assign _05026_ = _05015_ | \mchip.index [8];
	assign _05037_ = \mchip.index [9] & ~_05026_;
	assign _05048_ = _01953_ | _00198_;
	assign _05059_ = _05048_ | \mchip.index [4];
	assign _05070_ = _05059_ | \mchip.index [6];
	assign _05081_ = _05070_ | _07758_;
	assign _05092_ = _01986_ & ~_05081_;
	assign _05103_ = _00450_ | _04648_;
	assign _05114_ = _05103_ | \mchip.index [10];
	assign _05125_ = \mchip.index [11] & ~_05114_;
	assign _05136_ = _07714_ | _02984_;
	assign _05147_ = _05136_ | \mchip.index [8];
	assign _05158_ = _05147_ | \mchip.index [10];
	assign _05169_ = _01875_ & ~_05158_;
	assign _05180_ = \mchip.index [3] | \mchip.index [2];
	assign _05191_ = _05180_ | \mchip.index [4];
	assign _05203_ = _05191_ | _02984_;
	assign _05214_ = _05203_ | \mchip.index [7];
	assign _05225_ = _05214_ | _07758_;
	assign _05236_ = _05225_ | _01986_;
	assign _05247_ = _01875_ & ~_05236_;
	assign _05258_ = _05048_ | \mchip.index [6];
	assign _05269_ = _05258_ | \mchip.index [7];
	assign _05280_ = _05269_ | \mchip.index [10];
	assign _05291_ = _01875_ & ~_05280_;
	assign _05302_ = _01143_ | _02984_;
	assign _05314_ = _05302_ | \mchip.index [8];
	assign _05325_ = _07758_ & ~_05314_;
	assign _05336_ = _03650_ | _02984_;
	assign _05347_ = _05336_ | \mchip.index [7];
	assign _05358_ = _05347_ | \mchip.index [8];
	assign _05369_ = \mchip.index [9] & ~_05358_;
	assign _05380_ = _01964_ | _05424_;
	assign _05391_ = _05380_ | _02984_;
	assign _05402_ = _05391_ | \mchip.index [7];
	assign _05413_ = \mchip.index [9] & ~_05402_;
	assign _05425_ = _03860_ | _02984_;
	assign _05436_ = _05425_ | _02097_;
	assign _05447_ = _05436_ | _04648_;
	assign _05458_ = _05447_ | _07758_;
	assign _05469_ = _01875_ & ~_05458_;
	assign _05480_ = \mchip.index [3] | ~\mchip.index [2];
	assign _05491_ = _05480_ | \mchip.index [4];
	assign _05502_ = _05491_ | \mchip.index [5];
	assign _05513_ = _05502_ | \mchip.index [6];
	assign _05524_ = _05513_ | \mchip.index [7];
	assign _05536_ = _05524_ | _04648_;
	assign _05547_ = _05536_ | _07758_;
	assign _05558_ = _01875_ & ~_05547_;
	assign _05569_ = _04404_ | _04648_;
	assign _05580_ = _05569_ | _07758_;
	assign _05591_ = _05580_ | _01986_;
	assign _05602_ = _01875_ & ~_05591_;
	assign _05613_ = _01953_ | \mchip.index [5];
	assign _05624_ = _05613_ | \mchip.index [6];
	assign _05635_ = _05624_ | \mchip.index [8];
	assign _05647_ = _05635_ | _07758_;
	assign _05658_ = _05647_ | \mchip.index [10];
	assign _05669_ = \mchip.index [11] & ~_05658_;
	assign _05680_ = _01620_ | \mchip.index [3];
	assign _05691_ = _05680_ | \mchip.index [5];
	assign _05702_ = _05691_ | _02097_;
	assign _05713_ = _05702_ | _04648_;
	assign _05724_ = _05713_ | _01986_;
	assign _05735_ = _01875_ & ~_05724_;
	assign _05746_ = \mchip.index [4] | ~\mchip.index [1];
	assign _05758_ = _05746_ | \mchip.index [5];
	assign _05769_ = _05758_ | _02984_;
	assign _05780_ = _05769_ | \mchip.index [8];
	assign _05791_ = _05780_ | \mchip.index [9];
	assign _05802_ = \mchip.index [11] & ~_05791_;
	assign _05813_ = _00318_ | _02984_;
	assign _05824_ = _05813_ | _02097_;
	assign _05835_ = _05824_ | _04648_;
	assign _05846_ = _05835_ | _01986_;
	assign _05857_ = _01875_ & ~_05846_;
	assign _05869_ = _03084_ | \mchip.index [6];
	assign _05880_ = _05869_ | _02097_;
	assign _05891_ = _05880_ | _07758_;
	assign _05902_ = \mchip.index [11] & ~_05891_;
	assign _05913_ = _00670_ | _04648_;
	assign _05924_ = _05913_ | _01986_;
	assign _05935_ = _01875_ & ~_05924_;
	assign _05946_ = _00263_ | \mchip.index [4];
	assign _05957_ = _05946_ | \mchip.index [5];
	assign _05968_ = _05957_ | _02097_;
	assign _05980_ = _05968_ | _07758_;
	assign _05991_ = _05980_ | \mchip.index [10];
	assign _06002_ = _01875_ & ~_05991_;
	assign _06013_ = _01642_ | \mchip.index [8];
	assign _06024_ = _06013_ | _07758_;
	assign _06035_ = \mchip.index [10] & ~_06024_;
	assign _06046_ = _02518_ | \mchip.index [7];
	assign _06057_ = _06046_ | \mchip.index [10];
	assign _06068_ = \mchip.index [11] & ~_06057_;
	assign _06079_ = _01620_ | _02984_;
	assign _06091_ = _06079_ | _02097_;
	assign _06102_ = _06091_ | _07758_;
	assign _06113_ = _06102_ | \mchip.index [10];
	assign _06124_ = _01875_ & ~_06113_;
	assign _06135_ = _04759_ | \mchip.index [3];
	assign _06146_ = _06135_ | \mchip.index [6];
	assign _06157_ = _06146_ | _07758_;
	assign _06168_ = _06157_ | \mchip.index [10];
	assign _06179_ = _01875_ & ~_06168_;
	assign _06190_ = _05979_ | _02984_;
	assign _06202_ = _06190_ | _02097_;
	assign _06213_ = _06202_ | \mchip.index [8];
	assign _06224_ = _01986_ & ~_06213_;
	assign _06235_ = _01964_ | _01098_;
	assign _06246_ = _06235_ | \mchip.index [6];
	assign _06257_ = _06246_ | _02097_;
	assign _06268_ = _06257_ | \mchip.index [9];
	assign _06279_ = _01875_ & ~_06268_;
	assign _06290_ = _07703_ | \mchip.index [4];
	assign _06301_ = _06290_ | \mchip.index [7];
	assign _06313_ = _06301_ | _04648_;
	assign _06324_ = _06313_ | \mchip.index [9];
	assign _06335_ = \mchip.index [10] & ~_06324_;
	assign _06346_ = _03395_ | _05424_;
	assign _06356_ = _06346_ | _02984_;
	assign _06367_ = \mchip.index [10] & ~_06356_;
	assign _06378_ = _06977_ | \mchip.index [3];
	assign _06389_ = _06378_ | \mchip.index [4];
	assign _06400_ = _06389_ | _02097_;
	assign _06411_ = _06400_ | \mchip.index [8];
	assign _06423_ = _06411_ | \mchip.index [9];
	assign _06434_ = _01875_ & ~_06423_;
	assign _06445_ = _05191_ | \mchip.index [5];
	assign _06456_ = _06445_ | _02097_;
	assign _06467_ = _06456_ | _04648_;
	assign _06478_ = _01875_ & ~_06467_;
	assign _06489_ = _00263_ | \mchip.index [5];
	assign _06500_ = _06489_ | \mchip.index [6];
	assign _06511_ = _06500_ | \mchip.index [8];
	assign _06522_ = _06511_ | _07758_;
	assign _06534_ = \mchip.index [10] & ~_06522_;
	assign _06545_ = _00879_ | \mchip.index [4];
	assign _06556_ = _06545_ | \mchip.index [6];
	assign _06567_ = \mchip.index [11] & ~_06556_;
	assign _06578_ = _04993_ | \mchip.index [4];
	assign _06589_ = _06578_ | _02984_;
	assign _06600_ = _06589_ | _02097_;
	assign _06611_ = \mchip.index [10] & ~_06600_;
	assign _06622_ = _01964_ | \mchip.index [6];
	assign _06633_ = _06622_ | _02097_;
	assign _06645_ = _06633_ | _04648_;
	assign _06656_ = _01875_ & ~_06645_;
	assign _06667_ = _07659_ | \mchip.index [8];
	assign _06678_ = \mchip.index [11] & ~_06667_;
	assign _06689_ = _05979_ | \mchip.index [4];
	assign _06700_ = _06689_ | _02984_;
	assign _06711_ = _06700_ | _02097_;
	assign _06722_ = _06711_ | _07758_;
	assign _06733_ = \mchip.index [11] & ~_06722_;
	assign _06744_ = _06090_ | \mchip.index [5];
	assign _06756_ = _06744_ | \mchip.index [6];
	assign _06767_ = \mchip.index [11] & ~_06756_;
	assign _06778_ = _01209_ | _02984_;
	assign _06789_ = _06778_ | \mchip.index [7];
	assign _06800_ = _06789_ | \mchip.index [8];
	assign _06811_ = _06800_ | \mchip.index [9];
	assign _06822_ = \mchip.index [10] & ~_06811_;
	assign _06833_ = \mchip.index [4] | \mchip.index [1];
	assign _06844_ = _06833_ | \mchip.index [6];
	assign _06855_ = _06844_ | \mchip.index [7];
	assign _06867_ = _06855_ | _07758_;
	assign _06878_ = _06867_ | _01986_;
	assign _06889_ = _01875_ & ~_06878_;
	assign _06900_ = _01209_ | _01098_;
	assign _06911_ = _06900_ | \mchip.index [6];
	assign _06922_ = _06911_ | _04648_;
	assign _06933_ = _06922_ | \mchip.index [10];
	assign _06944_ = _01875_ & ~_06933_;
	assign _06955_ = _00923_ | \mchip.index [5];
	assign _06966_ = _06955_ | _02984_;
	assign _06978_ = _06966_ | \mchip.index [9];
	assign _06989_ = _06978_ | \mchip.index [10];
	assign _07000_ = \mchip.index [11] & ~_06989_;
	assign _07011_ = _05480_ | _05424_;
	assign _07022_ = _07011_ | \mchip.index [6];
	assign _07033_ = _07022_ | \mchip.index [8];
	assign _07044_ = \mchip.index [10] & ~_07033_;
	assign _07055_ = _03783_ | \mchip.index [6];
	assign _07066_ = _07055_ | _02097_;
	assign _07077_ = _07066_ | \mchip.index [8];
	assign _07089_ = _07077_ | \mchip.index [9];
	assign _07100_ = _07089_ | \mchip.index [10];
	assign _07111_ = \mchip.index [11] & ~_07100_;
	assign _07122_ = _00736_ | \mchip.index [9];
	assign _07133_ = \mchip.index [11] & ~_07122_;
	assign _07144_ = _03794_ | _02984_;
	assign _07155_ = _07144_ | _04648_;
	assign _07166_ = _07155_ | \mchip.index [9];
	assign _07177_ = _01875_ & ~_07166_;
	assign _07188_ = _06778_ | _02097_;
	assign _07200_ = _07188_ | \mchip.index [8];
	assign _07211_ = _07200_ | _07758_;
	assign _07222_ = \mchip.index [10] & ~_07211_;
	assign _07233_ = _05180_ | \mchip.index [5];
	assign _07244_ = _07233_ | \mchip.index [6];
	assign _07255_ = _07244_ | _02097_;
	assign _07266_ = _07255_ | _07758_;
	assign _07277_ = _07266_ | _01986_;
	assign _07288_ = _01875_ & ~_07277_;
	assign _07299_ = _07088_ | _01098_;
	assign _07311_ = _07299_ | \mchip.index [6];
	assign _07322_ = _07311_ | _04648_;
	assign _07333_ = _07322_ | _01986_;
	assign _07344_ = _01875_ & ~_07333_;
	assign _07355_ = _02629_ | _02984_;
	assign _07366_ = _07355_ | _04648_;
	assign _07377_ = _07366_ | \mchip.index [9];
	assign _07388_ = _01986_ & ~_07377_;
	assign _07399_ = _03395_ | \mchip.index [4];
	assign _07410_ = _07399_ | \mchip.index [6];
	assign _07422_ = _07410_ | _02097_;
	assign _07433_ = _07422_ | \mchip.index [8];
	assign _07444_ = _07758_ & ~_07433_;
	assign _07455_ = _02264_ | _02984_;
	assign _07466_ = _07455_ | _07758_;
	assign _07477_ = _01986_ & ~_07466_;
	assign _07488_ = _05491_ | _02097_;
	assign _07499_ = _07488_ | \mchip.index [8];
	assign _07510_ = \mchip.index [10] & ~_07499_;
	assign _07521_ = _00209_ | \mchip.index [5];
	assign _07533_ = _07521_ | \mchip.index [6];
	assign _07544_ = _07533_ | _02097_;
	assign _07555_ = \mchip.index [11] & ~_07544_;
	assign _07566_ = _03628_ | \mchip.index [8];
	assign _07577_ = \mchip.index [9] & ~_07566_;
	assign _07588_ = _02430_ | _00198_;
	assign _07599_ = _07588_ | \mchip.index [7];
	assign _07610_ = _07599_ | \mchip.index [9];
	assign _07621_ = _01986_ & ~_07610_;
	assign _07632_ = _07188_ | _04648_;
	assign _07638_ = _07632_ | \mchip.index [9];
	assign _07639_ = \mchip.index [10] & ~_07638_;
	assign _07640_ = _02253_ | _05424_;
	assign _07641_ = _07640_ | _07758_;
	assign _07642_ = _01875_ & ~_07641_;
	assign _07643_ = _00055_ | _04648_;
	assign _07644_ = _07643_ | \mchip.index [9];
	assign _07645_ = \mchip.index [11] & ~_07644_;
	assign _07646_ = _03960_ | \mchip.index [6];
	assign _07647_ = _07646_ | \mchip.index [9];
	assign _07649_ = \mchip.index [10] & ~_07647_;
	assign _07650_ = _04993_ | _04648_;
	assign _07651_ = _07650_ | \mchip.index [9];
	assign _07652_ = \mchip.index [10] & ~_07651_;
	assign _07653_ = _02319_ | _00198_;
	assign _07654_ = _07653_ | _01098_;
	assign _07655_ = _07654_ | _04648_;
	assign _07656_ = _07655_ | _07758_;
	assign _07657_ = _01875_ & ~_07656_;
	assign _07658_ = _00154_ | \mchip.index [5];
	assign _07660_ = _07658_ | _02097_;
	assign _07661_ = \mchip.index [10] & ~_07660_;
	assign _07662_ = _03306_ | \mchip.index [6];
	assign _07663_ = _07662_ | _02097_;
	assign _07664_ = _07663_ | \mchip.index [9];
	assign _07665_ = \mchip.index [10] & ~_07664_;
	assign _07666_ = _06545_ | \mchip.index [7];
	assign _07667_ = _07666_ | _04648_;
	assign _07668_ = _07667_ | _01986_;
	assign _07669_ = _01875_ & ~_07668_;
	assign _07671_ = _00923_ | _01098_;
	assign _07672_ = _07671_ | \mchip.index [6];
	assign _07673_ = _07672_ | \mchip.index [7];
	assign _07674_ = _01986_ & ~_07673_;
	assign _07675_ = _00318_ | _00198_;
	assign _07676_ = _07675_ | _01098_;
	assign _07677_ = _07676_ | _02984_;
	assign _07678_ = _07677_ | \mchip.index [9];
	assign _07679_ = \mchip.index [11] & ~_07678_;
	assign _07680_ = _02463_ | \mchip.index [7];
	assign _07682_ = _07680_ | \mchip.index [8];
	assign _07683_ = _07682_ | \mchip.index [9];
	assign _07684_ = \mchip.index [10] & ~_07683_;
	assign _07685_ = _00560_ | _01098_;
	assign _07686_ = _07685_ | \mchip.index [7];
	assign _07687_ = _07686_ | \mchip.index [8];
	assign _07688_ = _07687_ | \mchip.index [9];
	assign _07689_ = _01986_ & ~_07688_;
	assign _07690_ = _07658_ | _02984_;
	assign _07691_ = _07690_ | _07758_;
	assign _07693_ = _07691_ | \mchip.index [10];
	assign _07694_ = _01875_ & ~_07693_;
	assign _07695_ = _06445_ | _01986_;
	assign _07696_ = _01875_ & ~_07695_;
	assign _07697_ = _00923_ | \mchip.index [7];
	assign _07698_ = _07697_ | \mchip.index [8];
	assign _07699_ = _07698_ | _01986_;
	assign _07700_ = _01875_ & ~_07699_;
	assign _07701_ = _01099_ | \mchip.index [5];
	assign _07702_ = _07701_ | _04648_;
	assign _07704_ = _07702_ | \mchip.index [9];
	assign _07705_ = _01986_ & ~_07704_;
	assign _07706_ = _07199_ | _05424_;
	assign _07707_ = _07706_ | _02097_;
	assign _07708_ = \mchip.index [11] & ~_07707_;
	assign _07709_ = _00824_ | \mchip.index [6];
	assign _07710_ = _07709_ | \mchip.index [7];
	assign _07711_ = _04648_ & ~_07710_;
	assign _07712_ = _00263_ | _01098_;
	assign _07713_ = _07712_ | _02984_;
	assign _07715_ = _07713_ | _02097_;
	assign _07716_ = _07715_ | \mchip.index [10];
	assign _07717_ = \mchip.index [11] & ~_07716_;
	assign _07718_ = _01476_ | \mchip.index [7];
	assign _07719_ = _07758_ & ~_07718_;
	assign _07720_ = _06977_ | _02208_;
	assign _07721_ = _07720_ | _00198_;
	assign _07722_ = _07721_ | \mchip.index [8];
	assign _07723_ = \mchip.index [11] & ~_07722_;
	assign _07724_ = _07399_ | _04648_;
	assign _07726_ = _07724_ | \mchip.index [10];
	assign _07727_ = _01875_ & ~_07726_;
	assign _07728_ = _07088_ | _02984_;
	assign _07729_ = _07728_ | \mchip.index [7];
	assign _07730_ = _07729_ | _04648_;
	assign _07731_ = _07730_ | \mchip.index [9];
	assign _07732_ = _01986_ & ~_07731_;
	assign _07733_ = _06689_ | \mchip.index [6];
	assign _07734_ = _07733_ | _02097_;
	assign _07735_ = _07734_ | _04648_;
	assign _07737_ = _07758_ & ~_07735_;
	assign _07738_ = _02740_ | \mchip.index [8];
	assign _07739_ = _07738_ | _07758_;
	assign _07740_ = \mchip.index [11] & ~_07739_;
	assign _07741_ = _02408_ | _02984_;
	assign _07742_ = _07741_ | \mchip.index [7];
	assign _07743_ = _07742_ | _04648_;
	assign _07744_ = _01986_ & ~_07743_;
	assign _07745_ = _04993_ | _02984_;
	assign _07746_ = _07745_ | _02097_;
	assign _07748_ = _07746_ | _01986_;
	assign _07749_ = _01875_ & ~_07748_;
	assign _07750_ = _03406_ | \mchip.index [7];
	assign _07751_ = _07750_ | \mchip.index [9];
	assign _07752_ = \mchip.index [10] & ~_07751_;
	assign _07753_ = \mchip.index [4] | \mchip.index [0];
	assign _07754_ = _07753_ | \mchip.index [5];
	assign _07755_ = _07754_ | _02097_;
	assign _07756_ = _07755_ | \mchip.index [8];
	assign _07757_ = _07756_ | \mchip.index [9];
	assign _07759_ = _07757_ | \mchip.index [10];
	assign _07760_ = \mchip.index [11] & ~_07759_;
	assign _07761_ = \mchip.index [0] | ~\mchip.index [4];
	assign _07762_ = _07761_ | _02984_;
	assign _07763_ = _07762_ | _02097_;
	assign _07764_ = _07763_ | \mchip.index [8];
	assign _07765_ = _07764_ | \mchip.index [9];
	assign _07766_ = _07765_ | \mchip.index [10];
	assign _07767_ = _01875_ & ~_07766_;
	assign _07768_ = _06378_ | _01098_;
	assign _07770_ = _07768_ | \mchip.index [5];
	assign _07771_ = _07770_ | \mchip.index [6];
	assign _07772_ = _02097_ & ~_07771_;
	assign _07773_ = _00670_ | _01098_;
	assign _07774_ = _07773_ | \mchip.index [6];
	assign _07775_ = \mchip.index [9] & ~_07774_;
	assign _07776_ = _00780_ | \mchip.index [4];
	assign _07777_ = _07776_ | \mchip.index [6];
	assign _07778_ = _07777_ | _02097_;
	assign _07779_ = _07778_ | \mchip.index [8];
	assign _07781_ = _07779_ | _07758_;
	assign _07782_ = _01875_ & ~_07781_;
	assign _07783_ = _02320_ | \mchip.index [6];
	assign _07784_ = _07783_ | _07758_;
	assign _07785_ = \mchip.index [11] & ~_07784_;
	assign _07786_ = \mchip.index [5] & ~_07685_;
	assign _07787_ = _07088_ | \mchip.index [6];
	assign _07788_ = _07787_ | \mchip.index [8];
	assign _07789_ = _07788_ | \mchip.index [9];
	assign _07790_ = _01986_ & ~_07789_;
	assign _07792_ = _01431_ | \mchip.index [6];
	assign _07793_ = _07792_ | \mchip.index [7];
	assign _07794_ = _07758_ & ~_07793_;
	assign _07795_ = _02696_ | _02984_;
	assign _07796_ = _07795_ | _02097_;
	assign _07797_ = _04648_ & ~_07796_;
	assign _07798_ = _07088_ | \mchip.index [4];
	assign _07799_ = _07798_ | _02097_;
	assign _07800_ = _07799_ | _04648_;
	assign _07801_ = _07800_ | _07758_;
	assign _07803_ = _01875_ & ~_07801_;
	assign _07804_ = _04382_ | _01098_;
	assign _07805_ = _07804_ | _02097_;
	assign _07806_ = _07805_ | _04648_;
	assign _07807_ = _07806_ | _07758_;
	assign _07808_ = _01875_ & ~_07807_;
	assign _07809_ = _00824_ | _02097_;
	assign _07810_ = _07809_ | \mchip.index [9];
	assign _07811_ = \mchip.index [11] & ~_07810_;
	assign _07812_ = ~(\mchip.index [1] & \mchip.index [5]);
	assign _07814_ = _07812_ | \mchip.index [6];
	assign _07815_ = _07814_ | _02097_;
	assign _07816_ = _07815_ | \mchip.index [9];
	assign _07817_ = \mchip.index [11] & ~_07816_;
	assign _07818_ = _05336_ | \mchip.index [8];
	assign _07819_ = _07818_ | _07758_;
	assign _07820_ = \mchip.index [11] & ~_07819_;
	assign _07821_ = _04759_ | _01098_;
	assign _07822_ = _07821_ | _02984_;
	assign _07823_ = _07822_ | _02097_;
	assign _07825_ = _07823_ | \mchip.index [8];
	assign _07826_ = _07825_ | \mchip.index [9];
	assign _07827_ = _01875_ & ~_07826_;
	assign _07828_ = _05004_ | \mchip.index [4];
	assign _07829_ = _07828_ | \mchip.index [10];
	assign _07830_ = \mchip.index [11] & ~_07829_;
	assign _07831_ = _00527_ | _02097_;
	assign _07832_ = \mchip.index [8] & ~_07831_;
	assign _07833_ = _07653_ | _02984_;
	assign _07834_ = _07833_ | _02097_;
	assign _07836_ = _07834_ | _01986_;
	assign _07837_ = _01875_ & ~_07836_;
	assign _07838_ = _01875_ & ~_04804_;
	assign _07839_ = _06135_ | \mchip.index [4];
	assign _07840_ = _07839_ | _02097_;
	assign _07841_ = _07840_ | _07758_;
	assign _07842_ = _01986_ & ~_07841_;
	assign _07843_ = _05048_ | _01098_;
	assign _07844_ = _07843_ | \mchip.index [7];
	assign _07845_ = _07844_ | _01986_;
	assign _07847_ = \mchip.index [11] & ~_07845_;
	assign _07848_ = _02153_ | \mchip.index [4];
	assign _07849_ = _07848_ | _02097_;
	assign _07850_ = _07849_ | _04648_;
	assign _07851_ = _07850_ | _07758_;
	assign _07852_ = _01875_ & ~_07851_;
	assign _07853_ = _07088_ | _04648_;
	assign _07854_ = _07853_ | _07758_;
	assign _07855_ = _07854_ | _01986_;
	assign _07856_ = _01875_ & ~_07855_;
	assign _07858_ = _02618_ | \mchip.index [5];
	assign _07859_ = _07858_ | _02984_;
	assign _07860_ = _07859_ | \mchip.index [8];
	assign _07861_ = _07860_ | _07758_;
	assign _07862_ = _07861_ | _01986_;
	assign _07863_ = _01875_ & ~_07862_;
	assign _07864_ = _00835_ | \mchip.index [6];
	assign _07865_ = _07864_ | _07758_;
	assign _07866_ = \mchip.index [11] & ~_07865_;
	assign _07867_ = _04870_ | \mchip.index [7];
	assign _00001_ = _07867_ | _04648_;
	assign _00002_ = _00001_ | \mchip.index [10];
	assign _00003_ = \mchip.index [11] & ~_00002_;
	assign _00004_ = _03628_ | _02984_;
	assign _00005_ = _00004_ | \mchip.index [7];
	assign _00006_ = \mchip.index [9] & ~_00005_;
	assign _00007_ = _00006_ | _00003_;
	assign _00008_ = _00007_ | _07866_;
	assign _00009_ = _00008_ | _07863_;
	assign _00010_ = _00009_ | _07856_;
	assign _00012_ = _00010_ | _07852_;
	assign _00013_ = _00012_ | _07847_;
	assign _00014_ = _00013_ | _07842_;
	assign _00015_ = _00014_ | _07838_;
	assign _00016_ = _00015_ | _07837_;
	assign _00017_ = _00016_ | _07832_;
	assign _00018_ = _00017_ | _07830_;
	assign _00019_ = _00018_ | _07827_;
	assign _00020_ = _00019_ | _07820_;
	assign _00021_ = _00020_ | _07817_;
	assign _00023_ = _00021_ | _07811_;
	assign _00024_ = _00023_ | _07808_;
	assign _00025_ = _00024_ | _07803_;
	assign _00026_ = _00025_ | _07797_;
	assign _00027_ = _00026_ | _07794_;
	assign _00028_ = _00027_ | _07790_;
	assign _00029_ = _00028_ | _07786_;
	assign _00030_ = _00029_ | _07785_;
	assign _00031_ = _00030_ | _07782_;
	assign _00032_ = _00031_ | _07775_;
	assign _00034_ = _00032_ | _07772_;
	assign _00035_ = _00034_ | _07767_;
	assign _00036_ = _00035_ | _07760_;
	assign _00037_ = _00036_ | _07752_;
	assign _00038_ = _00037_ | _07749_;
	assign _00039_ = _00038_ | _07744_;
	assign _00040_ = _00039_ | _07740_;
	assign _00041_ = _00040_ | _07737_;
	assign _00042_ = _00041_ | _07732_;
	assign _00043_ = _00042_ | _07727_;
	assign _00045_ = _00043_ | _07723_;
	assign _00046_ = _00045_ | _07719_;
	assign _00047_ = _00046_ | _07717_;
	assign _00048_ = _00047_ | _07711_;
	assign _00049_ = _00048_ | _07708_;
	assign _00050_ = _00049_ | _07705_;
	assign _00051_ = _00050_ | _07700_;
	assign _00052_ = _00051_ | _07696_;
	assign _00053_ = _00052_ | _07694_;
	assign _00054_ = _00053_ | _07689_;
	assign _00056_ = _00054_ | _07684_;
	assign _00057_ = _00056_ | _07679_;
	assign _00058_ = _00057_ | _07674_;
	assign _00059_ = _00058_ | _07669_;
	assign _00060_ = _00059_ | _07665_;
	assign _00061_ = _00060_ | _07661_;
	assign _00062_ = _00061_ | _07657_;
	assign _00063_ = _00062_ | _07652_;
	assign _00064_ = _00063_ | _07649_;
	assign _00065_ = _00064_ | _07645_;
	assign _00067_ = _00065_ | _07642_;
	assign _00068_ = _00067_ | _07639_;
	assign _00069_ = _00068_ | _07621_;
	assign _00070_ = _00069_ | _07577_;
	assign _00071_ = _00070_ | _07555_;
	assign _00072_ = _00071_ | _07510_;
	assign _00073_ = _00072_ | _07477_;
	assign _00074_ = _00073_ | _07444_;
	assign _00075_ = _00074_ | _07388_;
	assign _00076_ = _00075_ | _07344_;
	assign _00078_ = _00076_ | _07288_;
	assign _00079_ = _00078_ | _07222_;
	assign _00080_ = _00079_ | _07177_;
	assign _00081_ = _00080_ | _07133_;
	assign _00082_ = _00081_ | _07111_;
	assign _00083_ = _00082_ | _07044_;
	assign _00084_ = _00083_ | _07000_;
	assign _00085_ = _00084_ | _06944_;
	assign _00086_ = _00085_ | _06889_;
	assign _00087_ = _00086_ | _06822_;
	assign _00089_ = _00087_ | _06767_;
	assign _00090_ = _00089_ | _06733_;
	assign _00091_ = _00090_ | _06678_;
	assign _00092_ = _00091_ | _06656_;
	assign _00093_ = _00092_ | _06611_;
	assign _00094_ = _00093_ | _06567_;
	assign _00095_ = _00094_ | _06534_;
	assign _00096_ = _00095_ | _06478_;
	assign _00097_ = _00096_ | _06434_;
	assign _00098_ = _00097_ | _06367_;
	assign _00100_ = _00098_ | _06335_;
	assign _00101_ = _00100_ | _06279_;
	assign _00102_ = _00101_ | _06224_;
	assign _00103_ = _00102_ | _06179_;
	assign _00104_ = _00103_ | _06124_;
	assign _00105_ = _00104_ | _06068_;
	assign _00106_ = _00105_ | _06035_;
	assign _00107_ = _00106_ | _06002_;
	assign _00108_ = _00107_ | _05935_;
	assign _00109_ = _00108_ | _05902_;
	assign _00111_ = _00109_ | _05857_;
	assign _00112_ = _00111_ | _05802_;
	assign _00113_ = _00112_ | _05735_;
	assign _00114_ = _00113_ | _05669_;
	assign _00115_ = _00114_ | _05602_;
	assign _00116_ = _00115_ | _05558_;
	assign _00117_ = _00116_ | _05469_;
	assign _00118_ = _00117_ | _05413_;
	assign _00119_ = _00118_ | _05369_;
	assign _00120_ = _00119_ | _05325_;
	assign _00122_ = _00120_ | _05291_;
	assign _00123_ = _00122_ | _05247_;
	assign _00124_ = _00123_ | _05169_;
	assign _00125_ = _00124_ | _05125_;
	assign _00126_ = _00125_ | _05092_;
	assign _00127_ = _00126_ | _05037_;
	assign _00128_ = _00127_ | _04982_;
	assign _00129_ = _00128_ | _04948_;
	assign _00130_ = _00129_ | _04915_;
	assign _00131_ = _00130_ | _04859_;
	assign _00133_ = _00131_ | _04826_;
	assign _00134_ = _00133_ | _04760_;
	assign _00135_ = _00134_ | _04726_;
	assign _00136_ = _00135_ | _04671_;
	assign _00137_ = _00136_ | _04615_;
	assign _00138_ = _00137_ | _04571_;
	assign _00139_ = _00138_ | _04538_;
	assign _00140_ = _00139_ | _04471_;
	assign _00141_ = _00140_ | _04438_;
	assign _00142_ = _00141_ | _04371_;
	assign _00144_ = _00142_ | _04338_;
	assign _00145_ = _00144_ | _04293_;
	assign _00146_ = _00145_ | _04238_;
	assign _00147_ = _00146_ | _04182_;
	assign _00148_ = _00147_ | _04138_;
	assign _00149_ = _00148_ | _04094_;
	assign _00150_ = _00149_ | _04049_;
	assign _00151_ = _00150_ | _04016_;
	assign _00152_ = _00151_ | _03949_;
	assign _00153_ = _00152_ | _03905_;
	assign _00155_ = _00153_ | _03849_;
	assign _00156_ = _00155_ | _03772_;
	assign _00157_ = _00156_ | _03728_;
	assign _00158_ = _00157_ | _03695_;
	assign _00159_ = _00158_ | _03662_;
	assign _00160_ = _00159_ | _03617_;
	assign _00161_ = _00160_ | _03584_;
	assign _00162_ = _00161_ | _03528_;
	assign _00163_ = _00162_ | _03495_;
	assign _00164_ = _00163_ | _03440_;
	assign _00166_ = _00164_ | _03384_;
	assign _00167_ = _00166_ | _03351_;
	assign _00168_ = _00167_ | _03295_;
	assign _00169_ = _00168_ | _03262_;
	assign _00170_ = _00169_ | _03229_;
	assign _00171_ = _00170_ | _03195_;
	assign _00172_ = _00171_ | _03140_;
	assign _00173_ = _00172_ | _03073_;
	assign _00174_ = _00173_ | _03018_;
	assign _00175_ = _00174_ | _02985_;
	assign _00177_ = _00175_ | _02918_;
	assign _00178_ = _00177_ | _02874_;
	assign _00179_ = _00178_ | _02829_;
	assign _00180_ = _00179_ | _02785_;
	assign _00181_ = _00180_ | _02729_;
	assign _00182_ = _00181_ | _02674_;
	assign _00183_ = _00182_ | _02607_;
	assign _00184_ = _00183_ | _02563_;
	assign _00185_ = _00184_ | _02507_;
	assign _00186_ = _00185_ | _02452_;
	assign _00188_ = _00186_ | _02397_;
	assign _00189_ = _00188_ | _02353_;
	assign _00190_ = _00189_ | _02308_;
	assign _00191_ = _00190_ | _02242_;
	assign _00192_ = _00191_ | _02197_;
	assign _00193_ = _00192_ | _02142_;
	assign _00194_ = _00193_ | _02098_;
	assign _00195_ = _00194_ | _02053_;
	assign _00196_ = _00195_ | _02020_;
	assign _00197_ = _00196_ | _01942_;
	assign _00199_ = _00197_ | _01887_;
	assign _00200_ = _00199_ | _01820_;
	assign _00201_ = _00200_ | _01765_;
	assign _00202_ = _00201_ | _01720_;
	assign _00203_ = _00202_ | _01676_;
	assign _00204_ = _00203_ | _01609_;
	assign _00205_ = _00204_ | _01554_;
	assign _00206_ = _00205_ | _01498_;
	assign _00207_ = _00206_ | _01465_;
	assign _00208_ = _00207_ | _01420_;
	assign _00210_ = _00208_ | _01365_;
	assign _00211_ = _00210_ | _01332_;
	assign _00212_ = _00211_ | _01287_;
	assign _00213_ = _00212_ | _01221_;
	assign _00214_ = _00213_ | _01176_;
	assign _00215_ = _00214_ | _01132_;
	assign _00216_ = _00215_ | _01088_;
	assign _00217_ = _00216_ | _01033_;
	assign _00218_ = _00217_ | _00978_;
	assign _00219_ = _00218_ | _00912_;
	assign _00221_ = _00219_ | _00868_;
	assign _00222_ = _00221_ | _00813_;
	assign _00223_ = _00222_ | _00769_;
	assign _00224_ = _00223_ | _00714_;
	assign _00225_ = _00224_ | _00659_;
	assign _00226_ = _00225_ | _00615_;
	assign _00227_ = _00226_ | _00549_;
	assign _00228_ = _00227_ | _00494_;
	assign _00229_ = _00228_ | _00439_;
	assign _00230_ = _00229_ | _00373_;
	assign _00232_ = _00230_ | _00307_;
	assign _00233_ = _00232_ | _00252_;
	assign _00234_ = _00233_ | _00187_;
	assign _00235_ = _00234_ | _00143_;
	assign _00236_ = _00235_ | _00088_;
	assign _00237_ = _00236_ | _00044_;
	assign _00238_ = _00237_ | _07857_;
	assign _00239_ = _00238_ | _07813_;
	assign _00240_ = _00239_ | _07747_;
	assign _00241_ = _00240_ | _07692_;
	assign _00243_ = _00241_ | _07532_;
	assign _00244_ = _00243_ | _06866_;
	assign _00245_ = _00244_ | _06422_;
	assign _00246_ = _00245_ | _05757_;
	assign _00247_ = _00246_ | _05313_;
	assign _00248_ = _00247_ | _04537_;
	assign _00249_ = _00248_ | _04093_;
	assign _00250_ = _00249_ | _03539_;
	assign _00251_ = _00250_ | _02873_;
	assign \mchip.val [6] = _00251_ | _01764_;
	assign _00253_ = _07839_ | \mchip.index [8];
	assign _00254_ = \mchip.index [11] & ~_00253_;
	assign _00255_ = _00329_ | _01098_;
	assign _00256_ = _00255_ | _02984_;
	assign _00257_ = _04648_ & ~_00256_;
	assign _00258_ = _07821_ | _02097_;
	assign _00259_ = _00258_ | _04648_;
	assign _00260_ = _07758_ & ~_00259_;
	assign _00261_ = _00879_ | _01098_;
	assign _00262_ = _00261_ | _02097_;
	assign _00264_ = _01875_ & ~_00262_;
	assign _00265_ = _01298_ | _04648_;
	assign _00266_ = _07758_ & ~_00265_;
	assign _00267_ = _01953_ | _01098_;
	assign _00268_ = _00267_ | \mchip.index [6];
	assign _00269_ = _00268_ | _07758_;
	assign _00270_ = _00269_ | \mchip.index [10];
	assign _00271_ = _01875_ & ~_00270_;
	assign _00272_ = _07804_ | \mchip.index [9];
	assign _00273_ = _00272_ | \mchip.index [10];
	assign _00275_ = _01875_ & ~_00273_;
	assign _00276_ = _07685_ | \mchip.index [5];
	assign _00277_ = _00276_ | \mchip.index [6];
	assign _00278_ = _00277_ | \mchip.index [7];
	assign _00279_ = \mchip.index [8] & ~_00278_;
	assign _00280_ = _02408_ | \mchip.index [6];
	assign _00281_ = _00280_ | _02097_;
	assign _00282_ = _00281_ | \mchip.index [9];
	assign _00283_ = _01875_ & ~_00282_;
	assign _00284_ = _05957_ | _04648_;
	assign _00286_ = \mchip.index [11] & ~_00284_;
	assign _00287_ = ~(\mchip.index [4] & \mchip.index [0]);
	assign _00288_ = _00287_ | _02097_;
	assign _00289_ = _00288_ | _04648_;
	assign _00290_ = \mchip.index [11] & ~_00289_;
	assign _00291_ = _04981_ | \mchip.index [7];
	assign _00292_ = _00291_ | _04648_;
	assign _00293_ = \mchip.index [11] & ~_00292_;
	assign _00294_ = _05491_ | \mchip.index [6];
	assign _00295_ = _00294_ | \mchip.index [7];
	assign _00297_ = _00295_ | \mchip.index [9];
	assign _00298_ = _01875_ & ~_00297_;
	assign _00299_ = _01953_ | _05424_;
	assign _00300_ = _00299_ | \mchip.index [7];
	assign _00301_ = \mchip.index [11] & ~_00300_;
	assign _00302_ = _01620_ | \mchip.index [5];
	assign _00303_ = _00302_ | \mchip.index [7];
	assign _00304_ = _00303_ | _07758_;
	assign _00305_ = \mchip.index [11] & ~_00304_;
	assign _00306_ = _05680_ | _02984_;
	assign _00308_ = _00306_ | _02097_;
	assign _00309_ = _00308_ | \mchip.index [8];
	assign _00310_ = _01986_ & ~_00309_;
	assign _00311_ = _03540_ | \mchip.index [5];
	assign _00312_ = _00311_ | \mchip.index [7];
	assign _00313_ = _00312_ | _07758_;
	assign _00314_ = \mchip.index [11] & ~_00313_;
	assign _00315_ = _01964_ | \mchip.index [4];
	assign _00316_ = _00315_ | _05424_;
	assign _00317_ = _00316_ | _02097_;
	assign _00319_ = _01875_ & ~_00317_;
	assign _00320_ = _01620_ | _01098_;
	assign _00321_ = _00320_ | _02097_;
	assign _00322_ = _00321_ | \mchip.index [10];
	assign _00323_ = \mchip.index [11] & ~_00322_;
	assign _00324_ = _07720_ | _01098_;
	assign _00325_ = _00324_ | _04648_;
	assign _00326_ = \mchip.index [11] & ~_00325_;
	assign _00327_ = \mchip.index [5] | ~\mchip.index [0];
	assign _00328_ = _00327_ | _02984_;
	assign _00330_ = _00328_ | _02097_;
	assign _00331_ = _00330_ | \mchip.index [8];
	assign _00332_ = _00331_ | \mchip.index [9];
	assign _00333_ = \mchip.index [11] & ~_00332_;
	assign _00334_ = _04870_ | \mchip.index [8];
	assign _00335_ = _00334_ | \mchip.index [9];
	assign _00336_ = \mchip.index [10] & ~_00335_;
	assign _00337_ = _07199_ | \mchip.index [6];
	assign _00338_ = _02097_ & ~_00337_;
	assign _00339_ = _00299_ | \mchip.index [6];
	assign _00341_ = \mchip.index [9] & ~_00339_;
	assign _00342_ = _07399_ | _02097_;
	assign _00343_ = _00342_ | _04648_;
	assign _00344_ = _01875_ & ~_00343_;
	assign _00345_ = _07721_ | \mchip.index [5];
	assign _00346_ = _00345_ | \mchip.index [7];
	assign _00347_ = \mchip.index [9] & ~_00346_;
	assign _00348_ = _00670_ | _05424_;
	assign _00349_ = _00348_ | \mchip.index [7];
	assign _00350_ = \mchip.index [8] & ~_00349_;
	assign _00352_ = _06977_ | _01098_;
	assign _00353_ = _00352_ | \mchip.index [6];
	assign _00354_ = _00353_ | _07758_;
	assign _00355_ = \mchip.index [10] & ~_00354_;
	assign _00356_ = _04637_ | _02097_;
	assign _00357_ = _04648_ & ~_00356_;
	assign _00358_ = _00835_ | \mchip.index [8];
	assign _00359_ = _01986_ & ~_00358_;
	assign _00360_ = _07761_ | \mchip.index [6];
	assign _00361_ = _00360_ | _02097_;
	assign _00363_ = _00361_ | \mchip.index [8];
	assign _00364_ = _00363_ | \mchip.index [9];
	assign _00365_ = _01986_ & ~_00364_;
	assign _00366_ = _05868_ | _01098_;
	assign _00367_ = _00366_ | _02097_;
	assign _00368_ = _00367_ | \mchip.index [8];
	assign _00369_ = \mchip.index [10] & ~_00368_;
	assign _00370_ = _03650_ | \mchip.index [5];
	assign _00371_ = _00370_ | _02097_;
	assign _00372_ = _00371_ | \mchip.index [8];
	assign _00374_ = \mchip.index [11] & ~_00372_;
	assign _00375_ = _07780_ | \mchip.index [9];
	assign _00376_ = _00375_ | \mchip.index [10];
	assign _00377_ = _01875_ & ~_00376_;
	assign _00378_ = _04926_ | _02097_;
	assign _00379_ = _01875_ & ~_00378_;
	assign _00380_ = _07648_ | \mchip.index [4];
	assign _00381_ = _00380_ | \mchip.index [5];
	assign _00382_ = _00381_ | _01986_;
	assign _00383_ = _01875_ & ~_00382_;
	assign _00385_ = \mchip.index [0] | \mchip.index [5];
	assign _00386_ = _00385_ | _02984_;
	assign _00387_ = _00386_ | \mchip.index [7];
	assign _00388_ = _00387_ | \mchip.index [8];
	assign _00389_ = _00388_ | _07758_;
	assign _00390_ = _00389_ | \mchip.index [10];
	assign _00391_ = \mchip.index [11] & ~_00390_;
	assign _00392_ = _07839_ | \mchip.index [7];
	assign _00393_ = _00392_ | _04648_;
	assign _00394_ = \mchip.index [10] & ~_00393_;
	assign _00396_ = _02685_ | \mchip.index [5];
	assign _00397_ = _00396_ | _02984_;
	assign _00398_ = _00397_ | \mchip.index [7];
	assign _00399_ = _07758_ & ~_00398_;
	assign _00400_ = _01654_ | \mchip.index [8];
	assign _00401_ = \mchip.index [11] & ~_00400_;
	assign _00402_ = _00461_ | _02097_;
	assign _00403_ = _00402_ | \mchip.index [8];
	assign _00404_ = \mchip.index [9] & ~_00403_;
	assign _00405_ = \mchip.index [6] | ~\mchip.index [0];
	assign _00407_ = _00405_ | _02097_;
	assign _00408_ = _00407_ | \mchip.index [8];
	assign _00409_ = _00408_ | _07758_;
	assign _00410_ = _01875_ & ~_00409_;
	assign _00411_ = _04871_ | \mchip.index [6];
	assign _00412_ = _04648_ & ~_00411_;
	assign _00413_ = _02796_ | _01986_;
	assign _00414_ = \mchip.index [11] & ~_00413_;
	assign _00415_ = _02618_ | _05424_;
	assign _00416_ = _00415_ | \mchip.index [6];
	assign _00418_ = _00416_ | _02097_;
	assign _00419_ = _00418_ | _04648_;
	assign _00420_ = \mchip.index [9] & ~_00419_;
	assign _00421_ = _07685_ | \mchip.index [6];
	assign _00422_ = _00421_ | \mchip.index [7];
	assign _00423_ = _07758_ & ~_00422_;
	assign _00424_ = \mchip.index [10] & ~_01753_;
	assign _00425_ = _00320_ | _02984_;
	assign _00426_ = _00425_ | _07758_;
	assign _00427_ = _01986_ & ~_00426_;
	assign _00429_ = _04193_ | _05424_;
	assign _00430_ = _00429_ | _02984_;
	assign _00431_ = _00430_ | _02097_;
	assign _00432_ = _01875_ & ~_00431_;
	assign _00433_ = _03650_ | _05424_;
	assign _00434_ = _00433_ | _02984_;
	assign _00435_ = _02097_ & ~_00434_;
	assign _00436_ = _07709_ | _07758_;
	assign _00437_ = \mchip.index [10] & ~_00436_;
	assign _00438_ = _01631_ | _02984_;
	assign _00440_ = _00438_ | \mchip.index [7];
	assign _00441_ = _00440_ | _01986_;
	assign _00442_ = _01875_ & ~_00441_;
	assign _00443_ = _04648_ & ~_00339_;
	assign _00444_ = \mchip.index [11] & ~_00846_;
	assign _00445_ = _00261_ | _07758_;
	assign _00446_ = \mchip.index [10] & ~_00445_;
	assign _00447_ = _07703_ | \mchip.index [5];
	assign _00448_ = _00447_ | \mchip.index [6];
	assign _00449_ = _00448_ | \mchip.index [7];
	assign _00451_ = _00449_ | _04648_;
	assign _00452_ = \mchip.index [10] & ~_00451_;
	assign _00453_ = _07648_ | \mchip.index [6];
	assign _00454_ = _00453_ | _07758_;
	assign _00455_ = \mchip.index [10] & ~_00454_;
	assign _00456_ = \mchip.index [0] | \mchip.index [6];
	assign _00457_ = _00456_ | _02097_;
	assign _00458_ = _00457_ | \mchip.index [8];
	assign _00459_ = _00458_ | \mchip.index [9];
	assign _00460_ = _00459_ | \mchip.index [10];
	assign _00462_ = _01875_ & ~_00460_;
	assign _00463_ = _00505_ | \mchip.index [4];
	assign _00464_ = _00463_ | \mchip.index [7];
	assign _00465_ = _01986_ & ~_00464_;
	assign _00466_ = _04682_ | _02097_;
	assign _00467_ = _00466_ | _04648_;
	assign _00468_ = \mchip.index [10] & ~_00467_;
	assign _00469_ = _02408_ | \mchip.index [5];
	assign _00470_ = _00469_ | \mchip.index [6];
	assign _00471_ = _00470_ | \mchip.index [7];
	assign _00473_ = \mchip.index [8] & ~_00471_;
	assign _00474_ = _05070_ | \mchip.index [7];
	assign _00475_ = \mchip.index [9] & ~_00474_;
	assign _00476_ = _07828_ | \mchip.index [5];
	assign _00477_ = \mchip.index [10] & ~_00476_;
	assign _00478_ = _07011_ | _02984_;
	assign _00479_ = _00478_ | _02097_;
	assign _00480_ = _01875_ & ~_00479_;
	assign _00481_ = _07839_ | _02984_;
	assign _00482_ = _07758_ & ~_00481_;
	assign _00484_ = _07648_ | \mchip.index [5];
	assign _00485_ = _00484_ | \mchip.index [9];
	assign _00486_ = \mchip.index [10] & ~_00485_;
	assign _00487_ = _07654_ | _02097_;
	assign _00488_ = \mchip.index [9] & ~_00487_;
	assign _00489_ = _00267_ | _01986_;
	assign _00490_ = \mchip.index [11] & ~_00489_;
	assign _00491_ = _00433_ | \mchip.index [7];
	assign _00492_ = _04648_ & ~_00491_;
	assign _00493_ = _07533_ | \mchip.index [8];
	assign _00495_ = _01875_ & ~_00493_;
	assign _00496_ = _01831_ | \mchip.index [5];
	assign _00497_ = _00496_ | _02984_;
	assign _00498_ = _00497_ | _02097_;
	assign _00499_ = _00498_ | _04648_;
	assign _00500_ = \mchip.index [9] & ~_00499_;
	assign _00501_ = _05048_ | \mchip.index [5];
	assign _00502_ = _00501_ | _04648_;
	assign _00503_ = _00502_ | \mchip.index [9];
	assign _00504_ = \mchip.index [10] & ~_00503_;
	assign _00506_ = _02253_ | \mchip.index [4];
	assign _00507_ = _00506_ | \mchip.index [5];
	assign _00508_ = _00507_ | _02984_;
	assign _00509_ = _00508_ | _04648_;
	assign _00510_ = \mchip.index [9] & ~_00509_;
	assign _00511_ = _00429_ | _04648_;
	assign _00512_ = _00511_ | \mchip.index [10];
	assign _00513_ = _01875_ & ~_00512_;
	assign _00514_ = _06578_ | \mchip.index [5];
	assign _00515_ = _00514_ | _02097_;
	assign _00517_ = _00515_ | _04648_;
	assign _00518_ = \mchip.index [9] & ~_00517_;
	assign _00519_ = _02463_ | \mchip.index [8];
	assign _00520_ = _00519_ | \mchip.index [9];
	assign _00521_ = \mchip.index [10] & ~_00520_;
	assign _00522_ = _02840_ | _04648_;
	assign _00523_ = _00522_ | \mchip.index [10];
	assign _00524_ = _01875_ & ~_00523_;
	assign _00525_ = _07804_ | _02984_;
	assign _00526_ = _00525_ | \mchip.index [7];
	assign _00528_ = _00526_ | \mchip.index [9];
	assign _00529_ = _01875_ & ~_00528_;
	assign _00530_ = _05004_ | \mchip.index [5];
	assign _00531_ = _00530_ | _02984_;
	assign _00532_ = \mchip.index [9] & ~_00531_;
	assign _00533_ = _05769_ | \mchip.index [7];
	assign _00534_ = _00533_ | _07758_;
	assign _00535_ = \mchip.index [10] & ~_00534_;
	assign _00536_ = _02463_ | _02097_;
	assign _00537_ = _00536_ | _04648_;
	assign _00539_ = _00537_ | _07758_;
	assign _00540_ = _01986_ & ~_00539_;
	assign _00541_ = _06977_ | \mchip.index [5];
	assign _00542_ = _00541_ | _01986_;
	assign _00543_ = \mchip.index [11] & ~_00542_;
	assign _00544_ = \mchip.index [6] | ~\mchip.index [2];
	assign _00545_ = _00544_ | \mchip.index [7];
	assign _00546_ = _00545_ | _04648_;
	assign _00547_ = _00546_ | \mchip.index [9];
	assign _00548_ = \mchip.index [10] & ~_00547_;
	assign _00550_ = _07637_ | \mchip.index [5];
	assign _00551_ = _00550_ | \mchip.index [7];
	assign _00552_ = _00551_ | \mchip.index [8];
	assign _00553_ = _07758_ & ~_00552_;
	assign _00554_ = _00267_ | \mchip.index [7];
	assign _00555_ = _00554_ | \mchip.index [8];
	assign _00556_ = _01875_ & ~_00555_;
	assign _00557_ = _06356_ | _02097_;
	assign _00558_ = \mchip.index [10] & ~_00557_;
	assign _00559_ = _01099_ | _01098_;
	assign _00561_ = _00559_ | \mchip.index [7];
	assign _00562_ = \mchip.index [10] & ~_00561_;
	assign _00563_ = _07646_ | _01986_;
	assign _00564_ = \mchip.index [11] & ~_00563_;
	assign _00565_ = \mchip.index [10] & ~_07736_;
	assign _00566_ = _02153_ | _01098_;
	assign _00567_ = _00566_ | _04648_;
	assign _00568_ = _00567_ | _07758_;
	assign _00569_ = _01875_ & ~_00568_;
	assign _00570_ = _06489_ | _02984_;
	assign _00572_ = _00570_ | \mchip.index [7];
	assign _00573_ = _00572_ | \mchip.index [8];
	assign _00574_ = _01986_ & ~_00573_;
	assign _00575_ = _02386_ | \mchip.index [8];
	assign _00576_ = \mchip.index [9] & ~_00575_;
	assign _00577_ = _07725_ | \mchip.index [6];
	assign _00578_ = _07758_ & ~_00577_;
	assign _00579_ = _04981_ | \mchip.index [8];
	assign _00580_ = \mchip.index [10] & ~_00579_;
	assign _00581_ = _01698_ | \mchip.index [9];
	assign _00583_ = _01875_ & ~_00581_;
	assign _00584_ = _00352_ | _02097_;
	assign _00585_ = _00584_ | \mchip.index [8];
	assign _00586_ = _07758_ & ~_00585_;
	assign _00587_ = _01320_ | _02984_;
	assign _00588_ = _00587_ | \mchip.index [9];
	assign _00589_ = _00588_ | \mchip.index [10];
	assign _00590_ = _01875_ & ~_00589_;
	assign _00591_ = _01376_ | \mchip.index [9];
	assign _00592_ = \mchip.index [11] & ~_00591_;
	assign _00594_ = \mchip.index [4] | ~\mchip.index [2];
	assign _00595_ = _00594_ | \mchip.index [5];
	assign _00596_ = _00595_ | _02984_;
	assign _00597_ = _00596_ | \mchip.index [7];
	assign _00598_ = _00597_ | _04648_;
	assign _00599_ = \mchip.index [11] & ~_00598_;
	assign _00600_ = _01044_ | \mchip.index [5];
	assign _00601_ = _00600_ | _02097_;
	assign _00602_ = _00601_ | _04648_;
	assign _00603_ = _01875_ & ~_00602_;
	assign _00605_ = _03739_ | \mchip.index [8];
	assign _00606_ = \mchip.index [9] & ~_00605_;
	assign _00607_ = _06135_ | _01098_;
	assign _00608_ = _00607_ | _07758_;
	assign _00609_ = _00608_ | _01986_;
	assign _00610_ = _01875_ & ~_00609_;
	assign _00611_ = _00370_ | _02984_;
	assign _00612_ = _00611_ | \mchip.index [8];
	assign _00613_ = \mchip.index [10] & ~_00612_;
	assign _00614_ = _00791_ | _02984_;
	assign _00616_ = _00614_ | _04648_;
	assign _00617_ = \mchip.index [11] & ~_00616_;
	assign _00618_ = _00384_ | \mchip.index [5];
	assign _00619_ = _00618_ | \mchip.index [8];
	assign _00620_ = _00619_ | \mchip.index [9];
	assign _00621_ = _01986_ & ~_00620_;
	assign _00622_ = _00596_ | _07758_;
	assign _00623_ = \mchip.index [11] & ~_00622_;
	assign _00624_ = _01209_ | \mchip.index [5];
	assign _00625_ = _00624_ | \mchip.index [6];
	assign _00627_ = _00625_ | _02097_;
	assign _00628_ = _00627_ | _04648_;
	assign _00629_ = \mchip.index [11] & ~_00628_;
	assign _00630_ = _05680_ | \mchip.index [4];
	assign _00631_ = _00630_ | \mchip.index [5];
	assign _00632_ = _00631_ | _02984_;
	assign _00633_ = _00632_ | _04648_;
	assign _00634_ = _01875_ & ~_00633_;
	assign _00635_ = _02319_ | _04648_;
	assign _00636_ = _00635_ | \mchip.index [9];
	assign _00638_ = \mchip.index [10] & ~_00636_;
	assign _00639_ = \mchip.index [4] | ~\mchip.index [0];
	assign _00640_ = _00639_ | \mchip.index [5];
	assign _00641_ = _00640_ | _02984_;
	assign _00642_ = _00641_ | \mchip.index [7];
	assign _00643_ = _00642_ | _04648_;
	assign _00644_ = \mchip.index [10] & ~_00643_;
	assign _00645_ = \mchip.index [10] & ~_03994_;
	assign _00646_ = _00302_ | \mchip.index [6];
	assign _00647_ = _00646_ | \mchip.index [7];
	assign _00649_ = _00647_ | _04648_;
	assign _00650_ = \mchip.index [11] & ~_00649_;
	assign _00651_ = _01831_ | _02984_;
	assign _00652_ = _00651_ | \mchip.index [7];
	assign _00653_ = _00652_ | \mchip.index [8];
	assign _00654_ = _07758_ & ~_00653_;
	assign _00655_ = _01687_ | \mchip.index [7];
	assign _00656_ = _00655_ | \mchip.index [9];
	assign _00657_ = _01875_ & ~_00656_;
	assign _00658_ = _06778_ | \mchip.index [8];
	assign _00660_ = _00658_ | \mchip.index [10];
	assign _00661_ = _01875_ & ~_00660_;
	assign _00662_ = _00571_ | \mchip.index [4];
	assign _00663_ = _00662_ | _02097_;
	assign _00664_ = _00663_ | \mchip.index [8];
	assign _00665_ = \mchip.index [10] & ~_00664_;
	assign _00666_ = _02685_ | _04648_;
	assign _00667_ = _00666_ | _07758_;
	assign _00668_ = _01986_ & ~_00667_;
	assign _00669_ = _00287_ | \mchip.index [5];
	assign _00671_ = _00669_ | _02097_;
	assign _00672_ = _00671_ | _04648_;
	assign _00673_ = _00672_ | _07758_;
	assign _00674_ = \mchip.index [10] & ~_00673_;
	assign _00675_ = _02529_ | _04648_;
	assign _00676_ = \mchip.index [11] & ~_00675_;
	assign _00677_ = _02618_ | \mchip.index [6];
	assign _00678_ = _00677_ | \mchip.index [7];
	assign _00679_ = _00678_ | \mchip.index [8];
	assign _00680_ = _00679_ | \mchip.index [9];
	assign _00682_ = _00680_ | \mchip.index [10];
	assign _00683_ = \mchip.index [11] & ~_00682_;
	assign _00684_ = _00923_ | _05424_;
	assign _00685_ = _00684_ | \mchip.index [8];
	assign _00686_ = \mchip.index [10] & ~_00685_;
	assign _00687_ = _02840_ | _02984_;
	assign _00688_ = _00687_ | _02097_;
	assign _00689_ = \mchip.index [8] & ~_00688_;
	assign _00690_ = _00099_ | \mchip.index [7];
	assign _00691_ = _00690_ | \mchip.index [9];
	assign _00693_ = _00691_ | \mchip.index [10];
	assign _00694_ = _01875_ & ~_00693_;
	assign _00695_ = _05957_ | _07758_;
	assign _00696_ = \mchip.index [11] & ~_00695_;
	assign _00697_ = _00626_ | _04648_;
	assign _00698_ = \mchip.index [9] & ~_00697_;
	assign _00699_ = _00639_ | \mchip.index [6];
	assign _00700_ = _00699_ | _02097_;
	assign _00701_ = _00700_ | \mchip.index [8];
	assign _00702_ = _00701_ | \mchip.index [9];
	assign _00704_ = \mchip.index [11] & ~_00702_;
	assign _00705_ = _04193_ | _01098_;
	assign _00706_ = _00705_ | \mchip.index [10];
	assign _00707_ = \mchip.index [11] & ~_00706_;
	assign _00708_ = _00395_ | \mchip.index [7];
	assign _00709_ = _07758_ & ~_00708_;
	assign _00710_ = _02408_ | \mchip.index [3];
	assign _00711_ = _00710_ | \mchip.index [8];
	assign _00712_ = \mchip.index [10] & ~_00711_;
	assign _00713_ = _07685_ | _02984_;
	assign _00715_ = _00713_ | _02097_;
	assign _00716_ = _00715_ | _04648_;
	assign _00717_ = _00716_ | \mchip.index [10];
	assign _00718_ = _01875_ & ~_00717_;
	assign _00719_ = _03650_ | _04648_;
	assign _00720_ = _00719_ | \mchip.index [9];
	assign _00721_ = _00720_ | \mchip.index [10];
	assign _00722_ = _01875_ & ~_00721_;
	assign _00723_ = _07804_ | \mchip.index [5];
	assign _00724_ = _00723_ | _02097_;
	assign _00726_ = \mchip.index [11] & ~_00724_;
	assign _00727_ = _00640_ | \mchip.index [6];
	assign _00728_ = _00727_ | _07758_;
	assign _00729_ = _00728_ | \mchip.index [10];
	assign _00730_ = _01875_ & ~_00729_;
	assign _00731_ = _00267_ | \mchip.index [9];
	assign _00732_ = \mchip.index [10] & ~_00731_;
	assign _00733_ = _00497_ | \mchip.index [9];
	assign _00734_ = \mchip.index [10] & ~_00733_;
	assign _00735_ = _00624_ | _02097_;
	assign _00737_ = _00735_ | \mchip.index [8];
	assign _00738_ = _00737_ | \mchip.index [9];
	assign _00739_ = \mchip.index [10] & ~_00738_;
	assign _00740_ = _00989_ | _02984_;
	assign _00741_ = \mchip.index [10] & ~_00740_;
	assign _00742_ = _00299_ | _07758_;
	assign _00743_ = \mchip.index [11] & ~_00742_;
	assign _00744_ = _06378_ | \mchip.index [5];
	assign _00745_ = _00744_ | _02984_;
	assign _00746_ = _00745_ | \mchip.index [8];
	assign _00748_ = _01986_ & ~_00746_;
	assign _00749_ = \mchip.index [5] | ~\mchip.index [2];
	assign _00750_ = _00749_ | _02984_;
	assign _00751_ = _00750_ | \mchip.index [7];
	assign _00752_ = _00751_ | \mchip.index [8];
	assign _00753_ = \mchip.index [9] & ~_00752_;
	assign _00754_ = _05048_ | _02984_;
	assign _00755_ = _00754_ | \mchip.index [8];
	assign _00756_ = _00755_ | \mchip.index [10];
	assign _00757_ = _01875_ & ~_00756_;
	assign _00759_ = _01642_ | _02984_;
	assign _00760_ = _00759_ | _07758_;
	assign _00761_ = _00760_ | _01986_;
	assign _00762_ = _01875_ & ~_00761_;
	assign _00763_ = _00055_ | _02984_;
	assign _00764_ = _00763_ | _02097_;
	assign _00765_ = _00764_ | _04648_;
	assign _00766_ = _01875_ & ~_00765_;
	assign _00767_ = _00570_ | _02097_;
	assign _00768_ = \mchip.index [10] & ~_00767_;
	assign _00770_ = _00670_ | _02097_;
	assign _00771_ = _00770_ | \mchip.index [8];
	assign _00772_ = _07758_ & ~_00771_;
	assign _00773_ = _05491_ | \mchip.index [7];
	assign _00774_ = _00773_ | _01986_;
	assign _00775_ = \mchip.index [11] & ~_00774_;
	assign _00776_ = _07653_ | \mchip.index [4];
	assign _00777_ = _00776_ | _02097_;
	assign _00778_ = _00777_ | \mchip.index [10];
	assign _00779_ = _01875_ & ~_00778_;
	assign _00781_ = _00318_ | _05424_;
	assign _00782_ = _00781_ | _02984_;
	assign _00783_ = _00782_ | _02097_;
	assign _00784_ = _07758_ & ~_00783_;
	assign _00785_ = _00662_ | _02984_;
	assign _00786_ = \mchip.index [11] & ~_00785_;
	assign _00787_ = \mchip.index [4] | ~\mchip.index [3];
	assign _00788_ = _00787_ | \mchip.index [5];
	assign _00789_ = _00788_ | _02984_;
	assign _00790_ = _00789_ | _04648_;
	assign _00792_ = \mchip.index [10] & ~_00790_;
	assign _00793_ = _01831_ | \mchip.index [7];
	assign _00794_ = _00793_ | _01986_;
	assign _00795_ = \mchip.index [11] & ~_00794_;
	assign _00796_ = _07675_ | \mchip.index [5];
	assign _00797_ = _00796_ | \mchip.index [6];
	assign _00798_ = _00797_ | _02097_;
	assign _00799_ = _00798_ | \mchip.index [9];
	assign _00800_ = _01875_ & ~_00799_;
	assign _00801_ = _07011_ | \mchip.index [8];
	assign _00803_ = _00801_ | \mchip.index [9];
	assign _00804_ = _01875_ & ~_00803_;
	assign _00805_ = _00453_ | \mchip.index [7];
	assign _00806_ = \mchip.index [11] & ~_00805_;
	assign _00807_ = _06966_ | \mchip.index [8];
	assign _00808_ = _00807_ | \mchip.index [9];
	assign _00809_ = _00808_ | \mchip.index [10];
	assign _00810_ = _01875_ & ~_00809_;
	assign _00811_ = _02618_ | _01098_;
	assign _00812_ = _00811_ | \mchip.index [8];
	assign _00814_ = _00812_ | _07758_;
	assign _00815_ = \mchip.index [10] & ~_00814_;
	assign _00816_ = _02685_ | _00198_;
	assign _00817_ = _00816_ | _02097_;
	assign _00818_ = \mchip.index [11] & ~_00817_;
	assign _00819_ = _04682_ | \mchip.index [6];
	assign _00820_ = _00819_ | \mchip.index [8];
	assign _00821_ = _01986_ & ~_00820_;
	assign _00822_ = _01776_ | _01098_;
	assign _00823_ = _00822_ | _04648_;
	assign _00825_ = _01986_ & ~_00823_;
	assign _00826_ = _05480_ | _01098_;
	assign _00827_ = _00826_ | _02984_;
	assign _00828_ = _00827_ | \mchip.index [7];
	assign _00829_ = _00828_ | _04648_;
	assign _00830_ = _01986_ & ~_00829_;
	assign _00831_ = _07745_ | \mchip.index [7];
	assign _00832_ = \mchip.index [9] & ~_00831_;
	assign _00833_ = _02364_ | _07758_;
	assign _00834_ = \mchip.index [11] & ~_00833_;
	assign _00836_ = _00000_ | _00198_;
	assign _00837_ = _00836_ | \mchip.index [4];
	assign _00838_ = _00837_ | \mchip.index [6];
	assign _00839_ = \mchip.index [8] & ~_00838_;
	assign _00840_ = _00554_ | _04648_;
	assign _00841_ = \mchip.index [11] & ~_00840_;
	assign _00842_ = _05702_ | _07758_;
	assign _00843_ = _01875_ & ~_00842_;
	assign _00844_ = _07714_ | \mchip.index [5];
	assign _00845_ = _00844_ | \mchip.index [6];
	assign _00847_ = _00845_ | _04648_;
	assign _00848_ = _07758_ & ~_00847_;
	assign _00849_ = _00630_ | _02984_;
	assign _00850_ = _00849_ | \mchip.index [9];
	assign _00851_ = \mchip.index [11] & ~_00850_;
	assign _00852_ = _02319_ | \mchip.index [6];
	assign _00853_ = _00852_ | _07758_;
	assign _00854_ = _00853_ | \mchip.index [10];
	assign _00855_ = _01875_ & ~_00854_;
	assign _00856_ = _02685_ | \mchip.index [4];
	assign _00858_ = _00856_ | _05424_;
	assign _00859_ = \mchip.index [9] & ~_00858_;
	assign _00860_ = _00461_ | \mchip.index [6];
	assign _00861_ = _04648_ & ~_00860_;
	assign _00862_ = _02419_ | \mchip.index [9];
	assign _00863_ = _01875_ & ~_00862_;
	assign _00864_ = _01565_ | _02097_;
	assign _00865_ = _00864_ | _04648_;
	assign _00866_ = _00865_ | \mchip.index [10];
	assign _00867_ = _01875_ & ~_00866_;
	assign _00869_ = _05502_ | _02984_;
	assign _00870_ = _00869_ | \mchip.index [8];
	assign _00871_ = \mchip.index [9] & ~_00870_;
	assign _00872_ = _06235_ | _02984_;
	assign _00873_ = _07758_ & ~_00872_;
	assign _00874_ = _07848_ | \mchip.index [9];
	assign _00875_ = _00874_ | \mchip.index [10];
	assign _00876_ = _01875_ & ~_00875_;
	assign _00877_ = _06833_ | _02984_;
	assign _00878_ = _00877_ | \mchip.index [7];
	assign _00880_ = _00878_ | _04648_;
	assign _00881_ = _00880_ | _07758_;
	assign _00882_ = _00881_ | _01986_;
	assign _00883_ = \mchip.index [11] & ~_00882_;
	assign _00884_ = _00450_ | _05424_;
	assign _00885_ = _00884_ | \mchip.index [6];
	assign _00886_ = \mchip.index [10] & ~_00885_;
	assign _00887_ = _00630_ | \mchip.index [6];
	assign _00888_ = _00887_ | _04648_;
	assign _00889_ = \mchip.index [10] & ~_00888_;
	assign _00891_ = _00626_ | \mchip.index [7];
	assign _00892_ = _01875_ & ~_00891_;
	assign _00893_ = \mchip.index [11] & ~_00337_;
	assign _00894_ = _04648_ & ~_01587_;
	assign _00895_ = _04582_ | _02097_;
	assign _00896_ = _00895_ | _04648_;
	assign _00897_ = _00896_ | _07758_;
	assign _00898_ = _01875_ & ~_00897_;
	assign _00899_ = _00898_ | _00894_;
	assign _00900_ = _00899_ | _00893_;
	assign _00902_ = _00900_ | _00892_;
	assign _00903_ = _00902_ | _00889_;
	assign _00904_ = _00903_ | _00886_;
	assign _00905_ = _00904_ | _00883_;
	assign _00906_ = _00905_ | _00876_;
	assign _00907_ = _00906_ | _00873_;
	assign _00908_ = _00907_ | _00871_;
	assign _00909_ = _00908_ | _00867_;
	assign _00910_ = _00909_ | _00863_;
	assign _00911_ = _00910_ | _00861_;
	assign _00913_ = _00911_ | _00859_;
	assign _00914_ = _00913_ | _00855_;
	assign _00915_ = _00914_ | _00851_;
	assign _00916_ = _00915_ | _00848_;
	assign _00917_ = _00916_ | _00843_;
	assign _00918_ = _00917_ | _00841_;
	assign _00919_ = _00918_ | _00839_;
	assign _00920_ = _00919_ | _00834_;
	assign _00921_ = _00920_ | _00832_;
	assign _00922_ = _00921_ | _00830_;
	assign _00924_ = _00922_ | _00825_;
	assign _00925_ = _00924_ | _00821_;
	assign _00926_ = _00925_ | _00818_;
	assign _00927_ = _00926_ | _00815_;
	assign _00928_ = _00927_ | _00810_;
	assign _00929_ = _00928_ | _00806_;
	assign _00930_ = _00929_ | _00804_;
	assign _00931_ = _00930_ | _00800_;
	assign _00932_ = _00931_ | _00795_;
	assign _00933_ = _00932_ | _00792_;
	assign _00935_ = _00933_ | _00786_;
	assign _00936_ = _00935_ | _00784_;
	assign _00937_ = _00936_ | _00779_;
	assign _00938_ = _00937_ | _00775_;
	assign _00939_ = _00938_ | _00772_;
	assign _00940_ = _00939_ | _00768_;
	assign _00941_ = _00940_ | _00766_;
	assign _00942_ = _00941_ | _00762_;
	assign _00943_ = _00942_ | _00757_;
	assign _00944_ = _00943_ | _00753_;
	assign _00946_ = _00944_ | _00748_;
	assign _00947_ = _00946_ | _00743_;
	assign _00948_ = _00947_ | _00741_;
	assign _00949_ = _00948_ | _00739_;
	assign _00950_ = _00949_ | _00734_;
	assign _00951_ = _00950_ | _00732_;
	assign _00952_ = _00951_ | _00730_;
	assign _00953_ = _00952_ | _00726_;
	assign _00954_ = _00953_ | _00722_;
	assign _00955_ = _00954_ | _00718_;
	assign _00957_ = _00955_ | _00712_;
	assign _00958_ = _00957_ | _00709_;
	assign _00959_ = _00958_ | _00707_;
	assign _00960_ = _00959_ | _00704_;
	assign _00961_ = _00960_ | _00698_;
	assign _00962_ = _00961_ | _00696_;
	assign _00963_ = _00962_ | _00694_;
	assign _00964_ = _00963_ | _00689_;
	assign _00965_ = _00964_ | _00686_;
	assign _00966_ = _00965_ | _00683_;
	assign _00968_ = _00966_ | _00676_;
	assign _00969_ = _00968_ | _00674_;
	assign _00970_ = _00969_ | _00668_;
	assign _00971_ = _00970_ | _00665_;
	assign _00972_ = _00971_ | _00661_;
	assign _00973_ = _00972_ | _00657_;
	assign _00974_ = _00973_ | _00654_;
	assign _00975_ = _00974_ | _00650_;
	assign _00976_ = _00975_ | _00645_;
	assign _00977_ = _00976_ | _00644_;
	assign _00979_ = _00977_ | _00638_;
	assign _00980_ = _00979_ | _00634_;
	assign _00981_ = _00980_ | _00629_;
	assign _00982_ = _00981_ | _00623_;
	assign _00983_ = _00982_ | _00621_;
	assign _00984_ = _00983_ | _00617_;
	assign _00985_ = _00984_ | _00613_;
	assign _00986_ = _00985_ | _00610_;
	assign _00987_ = _00986_ | _00606_;
	assign _00988_ = _00987_ | _00603_;
	assign _00990_ = _00988_ | _00599_;
	assign _00991_ = _00990_ | _00592_;
	assign _00992_ = _00991_ | _00590_;
	assign _00993_ = _00992_ | _00586_;
	assign _00994_ = _00993_ | _00583_;
	assign _00995_ = _00994_ | _00580_;
	assign _00996_ = _00995_ | _00578_;
	assign _00997_ = _00996_ | _00576_;
	assign _00998_ = _00997_ | _00574_;
	assign _00999_ = _00998_ | _00569_;
	assign _01001_ = _00999_ | _00565_;
	assign _01002_ = _01001_ | _00564_;
	assign _01003_ = _01002_ | _00562_;
	assign _01004_ = _01003_ | _00558_;
	assign _01005_ = _01004_ | _00556_;
	assign _01006_ = _01005_ | _00553_;
	assign _01007_ = _01006_ | _00548_;
	assign _01008_ = _01007_ | _00543_;
	assign _01009_ = _01008_ | _00540_;
	assign _01010_ = _01009_ | _00535_;
	assign _01012_ = _01010_ | _00532_;
	assign _01013_ = _01012_ | _00529_;
	assign _01014_ = _01013_ | _00524_;
	assign _01015_ = _01014_ | _00521_;
	assign _01016_ = _01015_ | _00518_;
	assign _01017_ = _01016_ | _00513_;
	assign _01018_ = _01017_ | _00510_;
	assign _01019_ = _01018_ | _00504_;
	assign _01020_ = _01019_ | _00500_;
	assign _01021_ = _01020_ | _00495_;
	assign _01023_ = _01021_ | _00492_;
	assign _01024_ = _01023_ | _00490_;
	assign _01025_ = _01024_ | _00488_;
	assign _01026_ = _01025_ | _00486_;
	assign _01027_ = _01026_ | _00482_;
	assign _01028_ = _01027_ | _00480_;
	assign _01029_ = _01028_ | _00477_;
	assign _01030_ = _01029_ | _00475_;
	assign _01031_ = _01030_ | _00473_;
	assign _01032_ = _01031_ | _00468_;
	assign _01034_ = _01032_ | _00465_;
	assign _01035_ = _01034_ | _00462_;
	assign _01036_ = _01035_ | _00455_;
	assign _01037_ = _01036_ | _00452_;
	assign _01038_ = _01037_ | _00446_;
	assign _01039_ = _01038_ | _00444_;
	assign _01040_ = _01039_ | _00443_;
	assign _01041_ = _01040_ | _00442_;
	assign _01042_ = _01041_ | _00437_;
	assign _01043_ = _01042_ | _00435_;
	assign _01045_ = _01043_ | _00432_;
	assign _01046_ = _01045_ | _00427_;
	assign _01047_ = _01046_ | _00424_;
	assign _01048_ = _01047_ | _00423_;
	assign _01049_ = _01048_ | _00420_;
	assign _01050_ = _01049_ | _00414_;
	assign _01051_ = _01050_ | _00412_;
	assign _01052_ = _01051_ | _00410_;
	assign _01053_ = _01052_ | _00404_;
	assign _01054_ = _01053_ | _00401_;
	assign _01056_ = _01054_ | _00399_;
	assign _01057_ = _01056_ | _00394_;
	assign _01058_ = _01057_ | _00391_;
	assign _01059_ = _01058_ | _00383_;
	assign _01060_ = _01059_ | _00379_;
	assign _01061_ = _01060_ | _00377_;
	assign _01062_ = _01061_ | _00374_;
	assign _01063_ = _01062_ | _00369_;
	assign _01064_ = _01063_ | _00365_;
	assign _01065_ = _01064_ | _00359_;
	assign _01067_ = _01065_ | _00357_;
	assign _01068_ = _01067_ | _00355_;
	assign _01069_ = _01068_ | _00350_;
	assign _01070_ = _01069_ | _00347_;
	assign _01071_ = _01070_ | _00344_;
	assign _01072_ = _01071_ | _00341_;
	assign _01073_ = _01072_ | _00338_;
	assign _01074_ = _01073_ | _00336_;
	assign _01075_ = _01074_ | _00333_;
	assign _01076_ = _01075_ | _00326_;
	assign _01078_ = _01076_ | _00323_;
	assign _01079_ = _01078_ | _00319_;
	assign _01080_ = _01079_ | _00314_;
	assign _01081_ = _01080_ | _00310_;
	assign _01082_ = _01081_ | _00305_;
	assign _01083_ = _01082_ | _00301_;
	assign _01084_ = _01083_ | _00298_;
	assign _01085_ = _01084_ | _00293_;
	assign _01086_ = _01085_ | _00290_;
	assign _01087_ = _01086_ | _00286_;
	assign _01089_ = _01087_ | _00283_;
	assign _01090_ = _01089_ | _00279_;
	assign _01091_ = _01090_ | _00275_;
	assign _01092_ = _01091_ | _00271_;
	assign _01093_ = _01092_ | _00266_;
	assign _01094_ = _01093_ | _00264_;
	assign _01095_ = _01094_ | _00260_;
	assign _01096_ = _01095_ | _00257_;
	assign \mchip.val [5] = _01096_ | _00254_;
	assign _01097_ = _03406_ | _02984_;
	assign _01100_ = _01097_ | _02097_;
	assign _01101_ = _01100_ | _04648_;
	assign _01102_ = _01101_ | _07758_;
	assign _01103_ = \mchip.index [10] & ~_01102_;
	assign _01104_ = _01476_ | \mchip.index [5];
	assign _01105_ = _01104_ | _02984_;
	assign _01106_ = _01105_ | _02097_;
	assign _01107_ = _01106_ | _04648_;
	assign _01108_ = _01107_ | \mchip.index [10];
	assign _01109_ = \mchip.index [11] & ~_01108_;
	assign _01111_ = _01099_ | \mchip.index [4];
	assign _01112_ = _01111_ | \mchip.index [5];
	assign _01113_ = _01112_ | \mchip.index [6];
	assign _01114_ = _01113_ | _02097_;
	assign _01115_ = _01114_ | _07758_;
	assign _01116_ = _01875_ & ~_01115_;
	assign _01117_ = _04071_ | _02097_;
	assign _01118_ = _01117_ | _01986_;
	assign _01119_ = \mchip.index [11] & ~_01118_;
	assign _01120_ = _07310_ | \mchip.index [5];
	assign _01122_ = _01120_ | \mchip.index [6];
	assign _01123_ = _01122_ | _04648_;
	assign _01124_ = _01123_ | _01986_;
	assign _01125_ = _01875_ & ~_01124_;
	assign _01126_ = _00710_ | \mchip.index [6];
	assign _01127_ = _01126_ | _02097_;
	assign _01128_ = _01127_ | _04648_;
	assign _01129_ = _01128_ | _01986_;
	assign _01130_ = _01875_ & ~_01129_;
	assign _01131_ = _07199_ | _01098_;
	assign _01133_ = _01131_ | \mchip.index [6];
	assign _01134_ = _01133_ | \mchip.index [7];
	assign _01135_ = _01134_ | _04648_;
	assign _01136_ = _01135_ | _07758_;
	assign _01137_ = _01986_ & ~_01136_;
	assign _01138_ = _03628_ | _02097_;
	assign _01139_ = _01138_ | _07758_;
	assign _01140_ = _01139_ | \mchip.index [10];
	assign _01141_ = \mchip.index [11] & ~_01140_;
	assign _01142_ = _07812_ | _02984_;
	assign _01144_ = _01142_ | _02097_;
	assign _01145_ = _01144_ | _07758_;
	assign _01146_ = \mchip.index [11] & ~_01145_;
	assign _01147_ = _05004_ | _01098_;
	assign _01148_ = _01147_ | \mchip.index [8];
	assign _01149_ = _01148_ | _07758_;
	assign _01150_ = _01149_ | \mchip.index [10];
	assign _01151_ = _01875_ & ~_01150_;
	assign _01152_ = _01376_ | \mchip.index [4];
	assign _01153_ = _01152_ | \mchip.index [5];
	assign _01155_ = _01153_ | _02984_;
	assign _01156_ = _01155_ | \mchip.index [8];
	assign _01157_ = _01156_ | \mchip.index [9];
	assign _01158_ = \mchip.index [10] & ~_01157_;
	assign _01159_ = _00710_ | _02984_;
	assign _01160_ = _01159_ | _02097_;
	assign _01161_ = _01160_ | _04648_;
	assign _01162_ = _01161_ | \mchip.index [9];
	assign _01163_ = _01162_ | \mchip.index [10];
	assign _01164_ = _01875_ & ~_01163_;
	assign _01166_ = _06689_ | \mchip.index [5];
	assign _01167_ = _01166_ | _02984_;
	assign _01168_ = _01167_ | \mchip.index [7];
	assign _01169_ = _01168_ | _04648_;
	assign _01170_ = _01169_ | _07758_;
	assign _01171_ = _01875_ & ~_01170_;
	assign _01172_ = _00559_ | _02984_;
	assign _01173_ = _01172_ | \mchip.index [7];
	assign _01174_ = _01173_ | \mchip.index [8];
	assign _01175_ = _01174_ | \mchip.index [9];
	assign _01177_ = \mchip.index [11] & ~_01175_;
	assign _01178_ = _07721_ | \mchip.index [4];
	assign _01179_ = _01178_ | _02984_;
	assign _01180_ = _01179_ | \mchip.index [7];
	assign _01181_ = _01180_ | _04648_;
	assign _01182_ = _01181_ | \mchip.index [9];
	assign _01183_ = \mchip.index [10] & ~_01182_;
	assign _01184_ = _07774_ | _02097_;
	assign _01185_ = _01184_ | _07758_;
	assign _01186_ = _01185_ | \mchip.index [10];
	assign _01188_ = _01875_ & ~_01186_;
	assign _01189_ = _02408_ | _00198_;
	assign _01190_ = _01189_ | _01098_;
	assign _01191_ = _01190_ | _02984_;
	assign _01192_ = _01191_ | _02097_;
	assign _01193_ = _01192_ | \mchip.index [8];
	assign _01194_ = _01193_ | \mchip.index [10];
	assign _01195_ = _01875_ & ~_01194_;
	assign _01196_ = _02685_ | _01098_;
	assign _01197_ = _01196_ | _02984_;
	assign _01199_ = _01197_ | _02097_;
	assign _01200_ = _01199_ | _07758_;
	assign _01201_ = \mchip.index [11] & ~_01200_;
	assign _01202_ = _06389_ | \mchip.index [6];
	assign _01203_ = _01202_ | \mchip.index [7];
	assign _01204_ = _01203_ | \mchip.index [8];
	assign _01205_ = _01204_ | _07758_;
	assign _01206_ = \mchip.index [10] & ~_01205_;
	assign _01207_ = _07798_ | \mchip.index [6];
	assign _01208_ = _01207_ | \mchip.index [7];
	assign _01211_ = _01208_ | _04648_;
	assign _01212_ = _01211_ | \mchip.index [9];
	assign _01213_ = \mchip.index [10] & ~_01212_;
	assign _01214_ = _00281_ | _04648_;
	assign _01215_ = _01214_ | _07758_;
	assign _01216_ = _01215_ | _01986_;
	assign _01217_ = _01875_ & ~_01216_;
	assign _01218_ = _00836_ | \mchip.index [6];
	assign _01219_ = _01218_ | _02097_;
	assign _01220_ = _01219_ | _04648_;
	assign _01222_ = _01220_ | \mchip.index [9];
	assign _01223_ = _01222_ | \mchip.index [10];
	assign _01224_ = _01875_ & ~_01223_;
	assign _01225_ = _00945_ | _02984_;
	assign _01226_ = _01225_ | _04648_;
	assign _01227_ = _01226_ | _07758_;
	assign _01228_ = _01227_ | _01986_;
	assign _01229_ = \mchip.index [11] & ~_01228_;
	assign _01230_ = _04993_ | _01098_;
	assign _01231_ = _01230_ | \mchip.index [6];
	assign _01233_ = _01231_ | _02097_;
	assign _01234_ = _01233_ | _04648_;
	assign _01235_ = _01234_ | \mchip.index [9];
	assign _01236_ = \mchip.index [10] & ~_01235_;
	assign _01237_ = _06689_ | \mchip.index [7];
	assign _01238_ = _01237_ | _04648_;
	assign _01239_ = _01238_ | \mchip.index [9];
	assign _01240_ = _01239_ | \mchip.index [10];
	assign _01241_ = _01875_ & ~_01240_;
	assign _01242_ = _07720_ | \mchip.index [3];
	assign _01244_ = _01242_ | _01098_;
	assign _01245_ = _01244_ | \mchip.index [6];
	assign _01246_ = _01245_ | _02097_;
	assign _01247_ = _01246_ | _04648_;
	assign _01248_ = \mchip.index [9] & ~_01247_;
	assign _01249_ = _07773_ | _02984_;
	assign _01250_ = _01249_ | _02097_;
	assign _01251_ = _01250_ | \mchip.index [8];
	assign _01252_ = \mchip.index [10] & ~_01251_;
	assign _01253_ = _07588_ | _01098_;
	assign _01255_ = _01253_ | _02984_;
	assign _01256_ = _01255_ | _02097_;
	assign _01257_ = _01256_ | \mchip.index [9];
	assign _01258_ = \mchip.index [10] & ~_01257_;
	assign _01259_ = _02441_ | _04648_;
	assign _01260_ = _01259_ | \mchip.index [9];
	assign _01261_ = \mchip.index [10] & ~_01260_;
	assign _01262_ = _07798_ | _02984_;
	assign _01263_ = _01262_ | _02097_;
	assign _01264_ = _01263_ | \mchip.index [8];
	assign _01266_ = _01264_ | \mchip.index [9];
	assign _01267_ = \mchip.index [10] & ~_01266_;
	assign _01268_ = _02153_ | _02984_;
	assign _01269_ = _01268_ | _02097_;
	assign _01270_ = _01269_ | _01986_;
	assign _01271_ = \mchip.index [11] & ~_01270_;
	assign _01272_ = _00816_ | _05424_;
	assign _01273_ = _01272_ | _02984_;
	assign _01274_ = _01273_ | \mchip.index [8];
	assign _01275_ = \mchip.index [9] & ~_01274_;
	assign _01277_ = _07676_ | \mchip.index [6];
	assign _01278_ = _01277_ | \mchip.index [7];
	assign _01279_ = _01278_ | _04648_;
	assign _01280_ = _01279_ | \mchip.index [9];
	assign _01281_ = \mchip.index [10] & ~_01280_;
	assign _01282_ = _00066_ | \mchip.index [8];
	assign _01283_ = _01282_ | \mchip.index [9];
	assign _01284_ = _01283_ | \mchip.index [10];
	assign _01285_ = _01875_ & ~_01284_;
	assign _01286_ = _07673_ | _04648_;
	assign _01288_ = _01286_ | \mchip.index [10];
	assign _01289_ = \mchip.index [11] & ~_01288_;
	assign _01290_ = _05680_ | _01098_;
	assign _01291_ = _01290_ | \mchip.index [5];
	assign _01292_ = _01291_ | _02984_;
	assign _01293_ = _01292_ | \mchip.index [7];
	assign _01294_ = _01293_ | _04648_;
	assign _01295_ = _01294_ | _07758_;
	assign _01296_ = \mchip.index [10] & ~_01295_;
	assign _01297_ = _02696_ | \mchip.index [5];
	assign _01299_ = _01297_ | _02984_;
	assign _01300_ = _01299_ | \mchip.index [7];
	assign _01301_ = _01300_ | \mchip.index [8];
	assign _01302_ = _01301_ | _07758_;
	assign _01303_ = \mchip.index [10] & ~_01302_;
	assign _01304_ = _07399_ | \mchip.index [5];
	assign _01305_ = _01304_ | \mchip.index [6];
	assign _01306_ = _01305_ | _02097_;
	assign _01307_ = _01306_ | \mchip.index [8];
	assign _01308_ = _01307_ | \mchip.index [9];
	assign _01310_ = \mchip.index [11] & ~_01308_;
	assign _01311_ = _07199_ | _02984_;
	assign _01312_ = _01311_ | _02097_;
	assign _01313_ = _01312_ | \mchip.index [8];
	assign _01314_ = _01313_ | \mchip.index [9];
	assign _01315_ = \mchip.index [10] & ~_01314_;
	assign _01316_ = _00209_ | \mchip.index [4];
	assign _01317_ = _01316_ | _02984_;
	assign _01318_ = _01317_ | \mchip.index [7];
	assign _01319_ = _01318_ | \mchip.index [8];
	assign _01322_ = _01319_ | \mchip.index [9];
	assign _01323_ = \mchip.index [11] & ~_01322_;
	assign _01324_ = _00329_ | \mchip.index [4];
	assign _01325_ = _01324_ | \mchip.index [5];
	assign _01326_ = _01325_ | _02984_;
	assign _01327_ = _01326_ | \mchip.index [7];
	assign _01328_ = _01327_ | \mchip.index [8];
	assign _01329_ = _01328_ | \mchip.index [9];
	assign _01330_ = _01329_ | _01986_;
	assign _01331_ = _01875_ & ~_01330_;
	assign _01333_ = _01172_ | _02097_;
	assign _01334_ = _01333_ | _04648_;
	assign _01335_ = \mchip.index [10] & ~_01334_;
	assign _01336_ = _00154_ | \mchip.index [6];
	assign _01337_ = _01336_ | \mchip.index [7];
	assign _01338_ = _01337_ | \mchip.index [8];
	assign _01339_ = _01338_ | _07758_;
	assign _01340_ = \mchip.index [10] & ~_01339_;
	assign _01341_ = _00710_ | _01098_;
	assign _01342_ = _01341_ | _02984_;
	assign _01344_ = _01342_ | \mchip.index [7];
	assign _01345_ = _01344_ | _07758_;
	assign _01346_ = _01875_ & ~_01345_;
	assign _01347_ = _01242_ | \mchip.index [5];
	assign _01348_ = _01347_ | \mchip.index [6];
	assign _01349_ = _01348_ | _02097_;
	assign _01350_ = _01349_ | \mchip.index [8];
	assign _01351_ = _01350_ | \mchip.index [9];
	assign _01352_ = \mchip.index [10] & ~_01351_;
	assign _01353_ = _05004_ | \mchip.index [6];
	assign _01355_ = _01353_ | \mchip.index [8];
	assign _01356_ = _01355_ | _07758_;
	assign _01357_ = _01356_ | \mchip.index [10];
	assign _01358_ = _01875_ & ~_01357_;
	assign _01359_ = _00261_ | \mchip.index [6];
	assign _01360_ = _01359_ | _02097_;
	assign _01361_ = _01360_ | \mchip.index [8];
	assign _01362_ = _01361_ | _07758_;
	assign _01363_ = \mchip.index [10] & ~_01362_;
	assign _01364_ = _00684_ | _02984_;
	assign _01366_ = _01364_ | _02097_;
	assign _01367_ = _01366_ | _04648_;
	assign _01368_ = \mchip.index [11] & ~_01367_;
	assign _01369_ = _01147_ | _02097_;
	assign _01370_ = _01369_ | \mchip.index [8];
	assign _01371_ = _01370_ | \mchip.index [9];
	assign _01372_ = \mchip.index [10] & ~_01371_;
	assign _01373_ = _02320_ | \mchip.index [5];
	assign _01374_ = _01373_ | \mchip.index [6];
	assign _01375_ = _01374_ | \mchip.index [7];
	assign _01377_ = _01375_ | \mchip.index [8];
	assign _01378_ = \mchip.index [10] & ~_01377_;
	assign _01379_ = _07721_ | _01098_;
	assign _01380_ = _01379_ | \mchip.index [6];
	assign _01381_ = _01380_ | _02097_;
	assign _01382_ = _01986_ & ~_01381_;
	assign _01383_ = _07588_ | \mchip.index [4];
	assign _01384_ = _01383_ | _02984_;
	assign _01385_ = _01384_ | _02097_;
	assign _01386_ = _01385_ | \mchip.index [9];
	assign _01388_ = _01986_ & ~_01386_;
	assign _01389_ = _00824_ | _01098_;
	assign _01390_ = _01389_ | \mchip.index [7];
	assign _01391_ = _01390_ | _04648_;
	assign _01392_ = _01391_ | _07758_;
	assign _01393_ = _01986_ & ~_01392_;
	assign _01394_ = _07706_ | _02984_;
	assign _01395_ = _01394_ | _02097_;
	assign _01396_ = _04648_ & ~_01395_;
	assign _01397_ = _00836_ | _01098_;
	assign _01399_ = _01397_ | _02097_;
	assign _01400_ = _01399_ | \mchip.index [8];
	assign _01401_ = _01400_ | \mchip.index [9];
	assign _01402_ = \mchip.index [10] & ~_01401_;
	assign _01403_ = _04893_ | _07758_;
	assign _01404_ = \mchip.index [11] & ~_01403_;
	assign _01405_ = _00934_ | \mchip.index [6];
	assign _01406_ = _01405_ | \mchip.index [7];
	assign _01407_ = _01406_ | \mchip.index [8];
	assign _01408_ = _01407_ | \mchip.index [9];
	assign _01410_ = _01408_ | \mchip.index [10];
	assign _01411_ = \mchip.index [11] & ~_01410_;
	assign _01412_ = _01341_ | \mchip.index [8];
	assign _01413_ = _01412_ | \mchip.index [9];
	assign _01414_ = \mchip.index [11] & ~_01413_;
	assign _01415_ = _00346_ | _01986_;
	assign _01416_ = \mchip.index [11] & ~_01415_;
	assign _01417_ = _00710_ | _05424_;
	assign _01418_ = _01417_ | _02984_;
	assign _01419_ = _01418_ | _07758_;
	assign _01421_ = \mchip.index [11] & ~_01419_;
	assign _01422_ = _00705_ | \mchip.index [6];
	assign _01423_ = _01422_ | \mchip.index [7];
	assign _01424_ = _01423_ | _04648_;
	assign _01425_ = _01424_ | \mchip.index [9];
	assign _01426_ = \mchip.index [11] & ~_01425_;
	assign _01427_ = _01242_ | \mchip.index [4];
	assign _01428_ = _01427_ | \mchip.index [5];
	assign _01429_ = _01428_ | \mchip.index [7];
	assign _01430_ = _01429_ | \mchip.index [8];
	assign _01433_ = _01430_ | \mchip.index [9];
	assign _01434_ = \mchip.index [11] & ~_01433_;
	assign _01435_ = _06257_ | \mchip.index [8];
	assign _01436_ = _01435_ | _07758_;
	assign _01437_ = \mchip.index [10] & ~_01436_;
	assign _01438_ = _01297_ | \mchip.index [6];
	assign _01439_ = _01438_ | _02097_;
	assign _01440_ = _01439_ | \mchip.index [8];
	assign _01441_ = \mchip.index [10] & ~_01440_;
	assign _01442_ = _00670_ | _02984_;
	assign _01444_ = _01442_ | _04648_;
	assign _01445_ = _01444_ | \mchip.index [9];
	assign _01446_ = \mchip.index [10] & ~_01445_;
	assign _01447_ = _05957_ | _02984_;
	assign _01448_ = _01447_ | \mchip.index [7];
	assign _01449_ = _01448_ | _01986_;
	assign _01450_ = \mchip.index [11] & ~_01449_;
	assign _01451_ = _01397_ | _02984_;
	assign _01452_ = _01451_ | \mchip.index [7];
	assign _01453_ = _01452_ | \mchip.index [8];
	assign _01455_ = \mchip.index [9] & ~_01453_;
	assign _01456_ = _01731_ | _02984_;
	assign _01457_ = _01456_ | \mchip.index [7];
	assign _01458_ = _01457_ | _04648_;
	assign _01459_ = _01458_ | \mchip.index [9];
	assign _01460_ = _01875_ & ~_01459_;
	assign _01461_ = _00816_ | \mchip.index [4];
	assign _01462_ = _01461_ | _02984_;
	assign _01463_ = _01462_ | \mchip.index [7];
	assign _01464_ = _01463_ | _04648_;
	assign _01466_ = _01464_ | _01986_;
	assign _01467_ = _01875_ & ~_01466_;
	assign _01468_ = _07310_ | _02984_;
	assign _01469_ = _01468_ | \mchip.index [8];
	assign _01470_ = _01469_ | \mchip.index [9];
	assign _01471_ = \mchip.index [10] & ~_01470_;
	assign _01472_ = _01197_ | \mchip.index [7];
	assign _01473_ = _01472_ | \mchip.index [8];
	assign _01474_ = _01473_ | \mchip.index [9];
	assign _01475_ = \mchip.index [10] & ~_01474_;
	assign _01477_ = _01190_ | \mchip.index [6];
	assign _01478_ = _01477_ | \mchip.index [7];
	assign _01479_ = _01478_ | _07758_;
	assign _01480_ = \mchip.index [10] & ~_01479_;
	assign _01481_ = _01397_ | \mchip.index [6];
	assign _01482_ = _01481_ | _02097_;
	assign _01483_ = _01482_ | _04648_;
	assign _01484_ = \mchip.index [11] & ~_01483_;
	assign _01485_ = _01244_ | _02984_;
	assign _01486_ = _01485_ | \mchip.index [7];
	assign _01488_ = _07758_ & ~_01486_;
	assign _01489_ = _01488_ & ~_01986_;
	assign _01490_ = \mchip.index [3] | ~\mchip.index [0];
	assign _01491_ = _01490_ | \mchip.index [4];
	assign _01492_ = _01491_ | \mchip.index [5];
	assign _01493_ = _01492_ | _02984_;
	assign _01494_ = _01493_ | \mchip.index [7];
	assign _01495_ = _01494_ | _01986_;
	assign _01496_ = \mchip.index [11] & ~_01495_;
	assign _01497_ = _01468_ | \mchip.index [7];
	assign _01499_ = _01497_ | _07758_;
	assign _01500_ = \mchip.index [11] & ~_01499_;
	assign _01501_ = _04993_ | _00198_;
	assign _01502_ = _01501_ | \mchip.index [4];
	assign _01503_ = _01502_ | _02984_;
	assign _01504_ = _01503_ | _02097_;
	assign _01505_ = _01504_ | \mchip.index [8];
	assign _01506_ = _01505_ | \mchip.index [10];
	assign _01507_ = _01875_ & ~_01506_;
	assign _01508_ = _00822_ | _02984_;
	assign _01510_ = _01508_ | _02097_;
	assign _01511_ = _01510_ | _04648_;
	assign _01512_ = _01511_ | \mchip.index [9];
	assign _01513_ = _01512_ | \mchip.index [10];
	assign _01514_ = _01875_ & ~_01513_;
	assign _01515_ = _07824_ | \mchip.index [5];
	assign _01516_ = _01515_ | \mchip.index [6];
	assign _01517_ = _01516_ | \mchip.index [7];
	assign _01518_ = _01517_ | _01986_;
	assign _01519_ = \mchip.index [11] & ~_01518_;
	assign _01521_ = _01256_ | _04648_;
	assign _01522_ = \mchip.index [9] & ~_01521_;
	assign _01523_ = _07654_ | _02984_;
	assign _01524_ = _01523_ | \mchip.index [7];
	assign _01525_ = _01524_ | \mchip.index [8];
	assign _01526_ = \mchip.index [11] & ~_01525_;
	assign _01527_ = _00315_ | \mchip.index [5];
	assign _01528_ = _01527_ | _02984_;
	assign _01529_ = _01528_ | _04648_;
	assign _01530_ = _01529_ | _07758_;
	assign _01532_ = _01530_ | \mchip.index [10];
	assign _01533_ = _01875_ & ~_01532_;
	assign _01534_ = _01189_ | \mchip.index [4];
	assign _01535_ = _01534_ | \mchip.index [6];
	assign _01536_ = _01535_ | \mchip.index [7];
	assign _01537_ = _01536_ | _04648_;
	assign _01538_ = _01537_ | \mchip.index [9];
	assign _01539_ = \mchip.index [10] & ~_01538_;
	assign _01540_ = _01534_ | \mchip.index [5];
	assign _01541_ = _01540_ | _02097_;
	assign _01544_ = _01541_ | \mchip.index [8];
	assign _01545_ = _01544_ | \mchip.index [9];
	assign _01546_ = \mchip.index [10] & ~_01545_;
	assign _01547_ = _01209_ | _05424_;
	assign _01548_ = _01547_ | _02984_;
	assign _01549_ = _01548_ | _04648_;
	assign _01550_ = _07758_ & ~_01549_;
	assign _01551_ = _00816_ | _01098_;
	assign _01552_ = _01551_ | _02984_;
	assign _01553_ = _01552_ | _02097_;
	assign _01555_ = _01553_ | _04648_;
	assign _01556_ = _01555_ | \mchip.index [10];
	assign _01557_ = _01875_ & ~_01556_;
	assign _01558_ = _00989_ | _05424_;
	assign _01559_ = _01558_ | _02984_;
	assign _01560_ = _07758_ & ~_01559_;
	assign _01561_ = _02408_ | \mchip.index [4];
	assign _01562_ = _01561_ | \mchip.index [5];
	assign _01563_ = _01562_ | _02984_;
	assign _01564_ = _01563_ | _02097_;
	assign _01566_ = _01564_ | \mchip.index [8];
	assign _01567_ = _01566_ | \mchip.index [9];
	assign _01568_ = \mchip.index [10] & ~_01567_;
	assign _01569_ = _00381_ | _02984_;
	assign _01570_ = _01569_ | _04648_;
	assign _01571_ = _01570_ | _07758_;
	assign _01572_ = _01986_ & ~_01571_;
	assign _01573_ = _01427_ | \mchip.index [6];
	assign _01574_ = _01573_ | _02097_;
	assign _01575_ = _01574_ | _07758_;
	assign _01577_ = _01575_ | \mchip.index [10];
	assign _01578_ = \mchip.index [11] & ~_01577_;
	assign _01579_ = _01180_ | \mchip.index [8];
	assign _01580_ = \mchip.index [11] & ~_01579_;
	assign _01581_ = _04759_ | _05424_;
	assign _01582_ = _01581_ | \mchip.index [6];
	assign _01583_ = _01582_ | _02097_;
	assign _01584_ = _01583_ | \mchip.index [8];
	assign _01585_ = \mchip.index [9] & ~_01584_;
	assign _01586_ = _06135_ | _05424_;
	assign _01588_ = _01586_ | _02984_;
	assign _01589_ = _01588_ | _07758_;
	assign _01590_ = _01986_ & ~_01589_;
	assign _01591_ = _01114_ | \mchip.index [10];
	assign _01592_ = _01875_ & ~_01591_;
	assign _01593_ = _07839_ | _05424_;
	assign _01594_ = _01593_ | \mchip.index [6];
	assign _01595_ = _01594_ | \mchip.index [7];
	assign _01596_ = _01595_ | _01986_;
	assign _01597_ = \mchip.index [11] & ~_01596_;
	assign _01599_ = _00824_ | _02984_;
	assign _01600_ = _01599_ | _02097_;
	assign _01601_ = _01600_ | _01986_;
	assign _01602_ = \mchip.index [11] & ~_01601_;
	assign _01603_ = _07780_ | _02984_;
	assign _01604_ = _01603_ | _02097_;
	assign _01605_ = _01604_ | _07758_;
	assign _01606_ = \mchip.index [11] & ~_01605_;
	assign _01607_ = _01551_ | \mchip.index [7];
	assign _01608_ = _01607_ | _04648_;
	assign _01610_ = _01608_ | _07758_;
	assign _01611_ = _01610_ | _01986_;
	assign _01612_ = _01875_ & ~_01611_;
	assign _01613_ = _01428_ | _02984_;
	assign _01614_ = _01613_ | \mchip.index [7];
	assign _01615_ = _01614_ | _04648_;
	assign _01616_ = _01615_ | _07758_;
	assign _01617_ = \mchip.index [10] & ~_01616_;
	assign _01618_ = _02540_ | \mchip.index [5];
	assign _01619_ = _01618_ | _02984_;
	assign _01621_ = _01619_ | _02097_;
	assign _01622_ = _01621_ | \mchip.index [8];
	assign _01623_ = _01622_ | \mchip.index [9];
	assign _01624_ = \mchip.index [11] & ~_01623_;
	assign _01625_ = _00476_ | _02984_;
	assign _01626_ = _01625_ | \mchip.index [7];
	assign _01627_ = _01626_ | \mchip.index [8];
	assign _01628_ = _01986_ & ~_01627_;
	assign _01629_ = _01383_ | \mchip.index [6];
	assign _01630_ = _01629_ | _04648_;
	assign _01632_ = _01630_ | _07758_;
	assign _01633_ = _01632_ | _01986_;
	assign _01634_ = _01875_ & ~_01633_;
	assign _01635_ = _01534_ | _02984_;
	assign _01636_ = _01635_ | \mchip.index [7];
	assign _01637_ = _01636_ | \mchip.index [8];
	assign _01638_ = _01637_ | _07758_;
	assign _01639_ = \mchip.index [10] & ~_01638_;
	assign _01640_ = _00776_ | \mchip.index [5];
	assign _01641_ = _01640_ | _02984_;
	assign _01643_ = _01641_ | _02097_;
	assign _01644_ = _01643_ | \mchip.index [9];
	assign _01645_ = _01644_ | \mchip.index [10];
	assign _01646_ = _01875_ & ~_01645_;
	assign _01647_ = _01625_ | _02097_;
	assign _01648_ = _01647_ | \mchip.index [8];
	assign _01649_ = \mchip.index [10] & ~_01648_;
	assign _01650_ = _01131_ | _02097_;
	assign _01651_ = _01650_ | _04648_;
	assign _01652_ = _01651_ | \mchip.index [10];
	assign _01655_ = \mchip.index [11] & ~_01652_;
	assign _01656_ = _06090_ | \mchip.index [6];
	assign _01657_ = _01656_ | _02097_;
	assign _01658_ = _01657_ | _04648_;
	assign _01659_ = _01658_ | \mchip.index [9];
	assign _01660_ = \mchip.index [10] & ~_01659_;
	assign _01661_ = _01462_ | _04648_;
	assign _01662_ = _01661_ | \mchip.index [10];
	assign _01663_ = \mchip.index [11] & ~_01662_;
	assign _01664_ = _01341_ | \mchip.index [6];
	assign _01666_ = _01664_ | _02097_;
	assign _01667_ = _01666_ | _07758_;
	assign _01668_ = _01667_ | _01986_;
	assign _01669_ = _01875_ & ~_01668_;
	assign _01670_ = _00476_ | \mchip.index [6];
	assign _01671_ = _01670_ | _02097_;
	assign _01672_ = _01671_ | _04648_;
	assign _01673_ = \mchip.index [11] & ~_01672_;
	assign _01674_ = _02540_ | _02984_;
	assign _01675_ = _01674_ | \mchip.index [7];
	assign _01677_ = _01675_ | \mchip.index [8];
	assign _01678_ = _01677_ | \mchip.index [9];
	assign _01679_ = \mchip.index [10] & ~_01678_;
	assign _01680_ = _04993_ | _05424_;
	assign _01681_ = _01680_ | _02984_;
	assign _01682_ = _01681_ | _02097_;
	assign _01683_ = _01682_ | \mchip.index [8];
	assign _01684_ = \mchip.index [11] & ~_01683_;
	assign _01685_ = _00476_ | _04648_;
	assign _01686_ = _01685_ | \mchip.index [10];
	assign _01688_ = \mchip.index [11] & ~_01686_;
	assign _01689_ = _01187_ | _02097_;
	assign _01690_ = _01689_ | _01986_;
	assign _01691_ = \mchip.index [11] & ~_01690_;
	assign _01692_ = _01394_ | \mchip.index [8];
	assign _01693_ = _01875_ & ~_01692_;
	assign _01694_ = _07770_ | \mchip.index [7];
	assign _01695_ = _01694_ | _01986_;
	assign _01696_ = \mchip.index [11] & ~_01695_;
	assign _01697_ = _02540_ | _05424_;
	assign _01699_ = _01697_ | \mchip.index [7];
	assign _01700_ = _01699_ | _07758_;
	assign _01701_ = \mchip.index [11] & ~_01700_;
	assign _01702_ = _01379_ | \mchip.index [7];
	assign _01703_ = _01702_ | \mchip.index [8];
	assign _01704_ = _01703_ | _07758_;
	assign _01705_ = \mchip.index [10] & ~_01704_;
	assign _01706_ = _03251_ | _01986_;
	assign _01707_ = \mchip.index [11] & ~_01706_;
	assign _01708_ = _04205_ | \mchip.index [5];
	assign _01710_ = _01708_ | \mchip.index [6];
	assign _01711_ = _01710_ | _02097_;
	assign _01712_ = _01711_ | _04648_;
	assign _01713_ = _01712_ | \mchip.index [9];
	assign _01714_ = _01713_ | \mchip.index [10];
	assign _01715_ = \mchip.index [11] & ~_01714_;
	assign _01716_ = _07721_ | \mchip.index [6];
	assign _01717_ = _01716_ | _02097_;
	assign _01718_ = _01717_ | _04648_;
	assign _01719_ = _01718_ | \mchip.index [9];
	assign _01721_ = _01986_ & ~_01719_;
	assign _01722_ = _07588_ | _02097_;
	assign _01723_ = _01722_ | \mchip.index [8];
	assign _01724_ = _01723_ | \mchip.index [9];
	assign _01725_ = _01724_ | \mchip.index [10];
	assign _01726_ = _01875_ & ~_01725_;
	assign _01727_ = _06900_ | \mchip.index [5];
	assign _01728_ = _01727_ | \mchip.index [6];
	assign _01729_ = _01728_ | \mchip.index [7];
	assign _01730_ = _01729_ | _01986_;
	assign _01732_ = \mchip.index [11] & ~_01730_;
	assign _01733_ = _05015_ | \mchip.index [7];
	assign _01734_ = _01733_ | _04648_;
	assign _01735_ = _01734_ | \mchip.index [9];
	assign _01736_ = \mchip.index [10] & ~_01735_;
	assign _01737_ = _00836_ | \mchip.index [5];
	assign _01738_ = _01737_ | \mchip.index [6];
	assign _01739_ = _01738_ | _02097_;
	assign _01740_ = _01739_ | \mchip.index [8];
	assign _01741_ = _01740_ | _07758_;
	assign _01743_ = \mchip.index [10] & ~_01741_;
	assign _01744_ = _07310_ | _05424_;
	assign _01745_ = _01744_ | \mchip.index [7];
	assign _01746_ = _01745_ | _01986_;
	assign _01747_ = \mchip.index [11] & ~_01746_;
	assign _01748_ = _01501_ | _01098_;
	assign _01749_ = _01748_ | \mchip.index [6];
	assign _01750_ = _01749_ | \mchip.index [7];
	assign _01751_ = _01750_ | _07758_;
	assign _01752_ = \mchip.index [11] & ~_01751_;
	assign _01754_ = _00315_ | _02984_;
	assign _01755_ = _01754_ | _02097_;
	assign _01756_ = _01755_ | _04648_;
	assign _01757_ = _01756_ | \mchip.index [9];
	assign _01758_ = _01757_ | _01986_;
	assign _01759_ = _01875_ & ~_01758_;
	assign _01760_ = _01629_ | \mchip.index [7];
	assign _01761_ = _01760_ | _04648_;
	assign _01762_ = _01761_ | _01986_;
	assign _01763_ = _01875_ & ~_01762_;
	assign _01766_ = _01155_ | _02097_;
	assign _01767_ = _01766_ | _04648_;
	assign _01768_ = _01767_ | _07758_;
	assign _01769_ = _01768_ | _01986_;
	assign _01770_ = _01875_ & ~_01769_;
	assign _01771_ = _00777_ | _07758_;
	assign _01772_ = _01771_ | \mchip.index [10];
	assign _01773_ = \mchip.index [11] & ~_01772_;
	assign _01774_ = _00000_ | _05424_;
	assign _01775_ = _01774_ | \mchip.index [6];
	assign _01777_ = _01775_ | \mchip.index [7];
	assign _01778_ = _01777_ | \mchip.index [8];
	assign _01779_ = \mchip.index [11] & ~_01778_;
	assign _01780_ = _01179_ | \mchip.index [8];
	assign _01781_ = _01780_ | \mchip.index [9];
	assign _01782_ = \mchip.index [11] & ~_01781_;
	assign _01783_ = _01178_ | _02097_;
	assign _01784_ = _01783_ | \mchip.index [8];
	assign _01785_ = _01784_ | _07758_;
	assign _01786_ = \mchip.index [10] & ~_01785_;
	assign _01788_ = _01670_ | \mchip.index [7];
	assign _01789_ = _01788_ | \mchip.index [8];
	assign _01790_ = _07758_ & ~_01789_;
	assign _01791_ = _02419_ | \mchip.index [6];
	assign _01792_ = _01791_ | _04648_;
	assign _01793_ = _01792_ | _07758_;
	assign _01794_ = _01793_ | _01986_;
	assign _01795_ = _01875_ & ~_01794_;
	assign _01796_ = _02320_ | _01098_;
	assign _01797_ = _01796_ | \mchip.index [6];
	assign _01799_ = _01797_ | _02097_;
	assign _01800_ = _01799_ | \mchip.index [8];
	assign _01801_ = \mchip.index [11] & ~_01800_;
	assign _01802_ = _00411_ | \mchip.index [7];
	assign _01803_ = _01802_ | \mchip.index [8];
	assign _01804_ = _07758_ & ~_01803_;
	assign _01805_ = _01431_ | _02984_;
	assign _01806_ = _01805_ | _02097_;
	assign _01807_ = _01806_ | \mchip.index [8];
	assign _01808_ = _01807_ | _07758_;
	assign _01810_ = \mchip.index [10] & ~_01808_;
	assign _01811_ = _01439_ | _04648_;
	assign _01812_ = _01811_ | _07758_;
	assign _01813_ = _01986_ & ~_01812_;
	assign _01814_ = _07828_ | _02097_;
	assign _01815_ = _01814_ | _07758_;
	assign _01816_ = _01815_ | \mchip.index [10];
	assign _01817_ = \mchip.index [11] & ~_01816_;
	assign _01818_ = _06246_ | \mchip.index [7];
	assign _01819_ = _01818_ | \mchip.index [8];
	assign _01821_ = _01819_ | _07758_;
	assign _01822_ = \mchip.index [11] & ~_01821_;
	assign _01823_ = _01776_ | \mchip.index [4];
	assign _01824_ = _01823_ | \mchip.index [6];
	assign _01825_ = _01824_ | \mchip.index [7];
	assign _01826_ = _01825_ | \mchip.index [10];
	assign _01827_ = _01875_ & ~_01826_;
	assign _01828_ = _01374_ | _02097_;
	assign _01829_ = _01828_ | \mchip.index [8];
	assign _01830_ = _01829_ | \mchip.index [9];
	assign _01832_ = \mchip.index [11] & ~_01830_;
	assign _01833_ = _05059_ | _02984_;
	assign _01834_ = _01833_ | _02097_;
	assign _01835_ = _01834_ | _04648_;
	assign _01836_ = _01835_ | \mchip.index [9];
	assign _01837_ = _01836_ | \mchip.index [10];
	assign _01838_ = _01875_ & ~_01837_;
	assign _01839_ = _00559_ | \mchip.index [6];
	assign _01840_ = _01839_ | \mchip.index [7];
	assign _01841_ = _01840_ | _04648_;
	assign _01843_ = _01841_ | _07758_;
	assign _01844_ = _01875_ & ~_01843_;
	assign _01845_ = \mchip.index [9] & ~_01193_;
	assign _01846_ = _02718_ | _01986_;
	assign _01847_ = \mchip.index [11] & ~_01846_;
	assign _01848_ = _07720_ | \mchip.index [4];
	assign _01849_ = _01848_ | \mchip.index [5];
	assign _01850_ = _01849_ | _02984_;
	assign _01851_ = _01850_ | _02097_;
	assign _01852_ = _01851_ | _04648_;
	assign _01854_ = _01852_ | _07758_;
	assign _01855_ = _01986_ & ~_01854_;
	assign _01856_ = ~(_02397_ & \mchip.index [10]);
	assign _01857_ = _01875_ & ~_01856_;
	assign _01858_ = _02264_ | \mchip.index [6];
	assign _01859_ = _01858_ | _02097_;
	assign _01860_ = _01859_ | _04648_;
	assign _01861_ = _01860_ | _01986_;
	assign _01862_ = _01875_ & ~_01861_;
	assign _01863_ = _00329_ | _05424_;
	assign _01865_ = _01863_ | \mchip.index [6];
	assign _01866_ = _01865_ | \mchip.index [8];
	assign _01867_ = _01866_ | \mchip.index [9];
	assign _01868_ = \mchip.index [11] & ~_01867_;
	assign _01869_ = _01383_ | \mchip.index [5];
	assign _01870_ = _01869_ | \mchip.index [6];
	assign _01871_ = _01870_ | _02097_;
	assign _01872_ = _01871_ | _07758_;
	assign _01873_ = \mchip.index [11] & ~_01872_;
	assign _01874_ = _07299_ | _02984_;
	assign _01877_ = _01874_ | _02097_;
	assign _01878_ = _01877_ | _07758_;
	assign _01879_ = _01878_ | \mchip.index [10];
	assign _01880_ = _01875_ & ~_01879_;
	assign _01881_ = _07311_ | _02097_;
	assign _01882_ = _01881_ | _07758_;
	assign _01883_ = _01882_ | \mchip.index [10];
	assign _01884_ = \mchip.index [11] & ~_01883_;
	assign _01885_ = _01643_ | \mchip.index [8];
	assign _01886_ = _01885_ | _07758_;
	assign _01888_ = \mchip.index [10] & ~_01886_;
	assign _01889_ = _01341_ | _02097_;
	assign _01890_ = _01889_ | \mchip.index [10];
	assign _01891_ = \mchip.index [11] & ~_01890_;
	assign _01892_ = _02685_ | _05424_;
	assign _01893_ = _01892_ | \mchip.index [6];
	assign _01894_ = _01893_ | _04648_;
	assign _01895_ = _01894_ | \mchip.index [9];
	assign _01896_ = \mchip.index [11] & ~_01895_;
	assign _01897_ = \mchip.index [11] & ~_01626_;
	assign _01899_ = _06389_ | \mchip.index [5];
	assign _01900_ = _01899_ | \mchip.index [6];
	assign _01901_ = _01900_ | _02097_;
	assign _01902_ = _01901_ | \mchip.index [9];
	assign _01903_ = \mchip.index [10] & ~_01902_;
	assign _01904_ = _02430_ | _05424_;
	assign _01905_ = _01904_ | \mchip.index [7];
	assign _01906_ = _01905_ | \mchip.index [9];
	assign _01907_ = \mchip.index [10] & ~_01906_;
	assign _01908_ = _00710_ | \mchip.index [5];
	assign _01910_ = _01908_ | _02097_;
	assign _01911_ = _01910_ | \mchip.index [8];
	assign _01912_ = _01911_ | \mchip.index [9];
	assign _01913_ = \mchip.index [11] & ~_01912_;
	assign _01914_ = _01387_ | \mchip.index [6];
	assign _01915_ = _01914_ | \mchip.index [8];
	assign _01916_ = _01915_ | \mchip.index [9];
	assign _01917_ = \mchip.index [11] & ~_01916_;
	assign _01918_ = _01796_ | _02984_;
	assign _01919_ = _01918_ | _02097_;
	assign _01921_ = _01919_ | \mchip.index [8];
	assign _01922_ = _01921_ | _07758_;
	assign _01923_ = \mchip.index [10] & ~_01922_;
	assign _01924_ = _01000_ | \mchip.index [6];
	assign _01925_ = _01924_ | \mchip.index [7];
	assign _01926_ = _01925_ | _07758_;
	assign _01927_ = _01926_ | _01986_;
	assign _01928_ = _01875_ & ~_01927_;
	assign _01929_ = _04893_ | \mchip.index [7];
	assign _01930_ = _01929_ | \mchip.index [9];
	assign _01932_ = \mchip.index [10] & ~_01930_;
	assign _01933_ = _01131_ | \mchip.index [5];
	assign _01934_ = _01933_ | _02984_;
	assign _01935_ = _01934_ | _04648_;
	assign _01936_ = \mchip.index [11] & ~_01935_;
	assign _01937_ = _07839_ | \mchip.index [6];
	assign _01938_ = _01937_ | \mchip.index [7];
	assign _01939_ = _01938_ | \mchip.index [9];
	assign _01940_ = _01939_ | \mchip.index [10];
	assign _01941_ = _01875_ & ~_01940_;
	assign _01943_ = _04871_ | \mchip.index [4];
	assign _01944_ = _01943_ | \mchip.index [6];
	assign _01945_ = _01944_ | \mchip.index [7];
	assign _01946_ = _01945_ | _04648_;
	assign _01947_ = _01946_ | _07758_;
	assign _01948_ = _01986_ & ~_01947_;
	assign _01949_ = _00710_ | \mchip.index [4];
	assign _01950_ = _01949_ | _02984_;
	assign _01951_ = _01950_ | _02097_;
	assign _01952_ = _01951_ | \mchip.index [8];
	assign _01954_ = _01952_ | _07758_;
	assign _01955_ = _01986_ & ~_01954_;
	assign _01956_ = _01953_ | \mchip.index [4];
	assign _01957_ = _01956_ | \mchip.index [5];
	assign _01958_ = _01957_ | \mchip.index [6];
	assign _01959_ = _01958_ | \mchip.index [7];
	assign _01960_ = _01959_ | _04648_;
	assign _01961_ = _01960_ | _07758_;
	assign _01962_ = _01961_ | _01986_;
	assign _01963_ = \mchip.index [11] & ~_01962_;
	assign _01965_ = _04871_ | \mchip.index [5];
	assign _01966_ = _01965_ | \mchip.index [6];
	assign _01967_ = _01966_ | \mchip.index [8];
	assign _01968_ = _01967_ | \mchip.index [9];
	assign _01969_ = _01986_ & ~_01968_;
	assign _01970_ = _07648_ | _05424_;
	assign _01971_ = _01970_ | _02984_;
	assign _01972_ = _01971_ | _02097_;
	assign _01973_ = _01972_ | \mchip.index [9];
	assign _01974_ = \mchip.index [10] & ~_01973_;
	assign _01976_ = _01511_ | _07758_;
	assign _01977_ = \mchip.index [10] & ~_01976_;
	assign _01978_ = _01833_ | \mchip.index [7];
	assign _01979_ = _01978_ | _04648_;
	assign _01980_ = _01979_ | _07758_;
	assign _01981_ = _01980_ | _01986_;
	assign _01982_ = _01875_ & ~_01981_;
	assign _01983_ = _01207_ | _02097_;
	assign _01984_ = _01983_ | _04648_;
	assign _01985_ = _01984_ | _07758_;
	assign _01988_ = _01985_ | _01986_;
	assign _01989_ = _01875_ & ~_01988_;
	assign _01990_ = _01152_ | _02984_;
	assign _01991_ = _01990_ | _04648_;
	assign _01992_ = _01991_ | \mchip.index [9];
	assign _01993_ = _01992_ | \mchip.index [10];
	assign _01994_ = _01875_ & ~_01993_;
	assign _01995_ = _01387_ | \mchip.index [7];
	assign _01996_ = _01995_ | \mchip.index [8];
	assign _01997_ = _01996_ | _07758_;
	assign _01999_ = \mchip.index [10] & ~_01997_;
	assign _02000_ = _01418_ | _02097_;
	assign _02001_ = \mchip.index [9] & ~_02000_;
	assign _02002_ = _01110_ | _02984_;
	assign _02003_ = _02002_ | _02097_;
	assign _02004_ = _02003_ | _04648_;
	assign _02005_ = \mchip.index [9] & ~_02004_;
	assign _02006_ = _01373_ | _02984_;
	assign _02007_ = _02006_ | \mchip.index [7];
	assign _02008_ = _02007_ | _01986_;
	assign _02010_ = \mchip.index [11] & ~_02008_;
	assign _02011_ = _01242_ | _05424_;
	assign _02012_ = _02011_ | \mchip.index [6];
	assign _02013_ = _02012_ | _02097_;
	assign _02014_ = \mchip.index [11] & ~_02013_;
	assign _02015_ = _00776_ | \mchip.index [6];
	assign _02016_ = _02015_ | \mchip.index [7];
	assign _02017_ = _02016_ | _04648_;
	assign _02018_ = _02017_ | \mchip.index [10];
	assign _02019_ = \mchip.index [11] & ~_02018_;
	assign _02021_ = _03240_ | \mchip.index [6];
	assign _02022_ = _02021_ | \mchip.index [7];
	assign _02023_ = _02022_ | \mchip.index [10];
	assign _02024_ = _01875_ & ~_02023_;
	assign _02025_ = _01796_ | \mchip.index [8];
	assign _02026_ = _02025_ | \mchip.index [9];
	assign _02027_ = _02026_ | \mchip.index [10];
	assign _02028_ = _01875_ & ~_02027_;
	assign _02029_ = _01427_ | _02984_;
	assign _02030_ = _02029_ | _04648_;
	assign _02032_ = _02030_ | \mchip.index [10];
	assign _02033_ = \mchip.index [11] & ~_02032_;
	assign _02034_ = _00571_ | _05424_;
	assign _02035_ = _02034_ | \mchip.index [6];
	assign _02036_ = _02035_ | _02097_;
	assign _02037_ = _02036_ | \mchip.index [9];
	assign _02038_ = \mchip.index [10] & ~_02037_;
	assign _02039_ = _00631_ | \mchip.index [6];
	assign _02040_ = _02039_ | _02097_;
	assign _02041_ = _02040_ | _01986_;
	assign _02043_ = \mchip.index [11] & ~_02041_;
	assign _02044_ = _00945_ | \mchip.index [6];
	assign _02045_ = _02044_ | \mchip.index [7];
	assign _02046_ = _02045_ | \mchip.index [8];
	assign _02047_ = _02046_ | _07758_;
	assign _02048_ = _02047_ | _01986_;
	assign _02049_ = _01875_ & ~_02048_;
	assign _02050_ = _00514_ | _02984_;
	assign _02051_ = _02050_ | _02097_;
	assign _02052_ = _02051_ | \mchip.index [8];
	assign _02054_ = _02052_ | \mchip.index [9];
	assign _02055_ = _02054_ | \mchip.index [10];
	assign _02056_ = _01875_ & ~_02055_;
	assign _02057_ = _01112_ | _02984_;
	assign _02058_ = _02057_ | \mchip.index [7];
	assign _02059_ = _02058_ | \mchip.index [9];
	assign _02060_ = _02059_ | \mchip.index [10];
	assign _02061_ = _01875_ & ~_02060_;
	assign _02062_ = _01636_ | \mchip.index [9];
	assign _02063_ = \mchip.index [11] & ~_02062_;
	assign _02065_ = _00541_ | _02984_;
	assign _02066_ = _02065_ | \mchip.index [7];
	assign _02067_ = _02066_ | _01986_;
	assign _02068_ = \mchip.index [11] & ~_02067_;
	assign _02069_ = _03051_ | _04648_;
	assign _02070_ = _02069_ | \mchip.index [9];
	assign _02071_ = \mchip.index [11] & ~_02070_;
	assign _02072_ = _00776_ | _05424_;
	assign _02073_ = _02072_ | \mchip.index [6];
	assign _02074_ = _02097_ & ~_02073_;
	assign _02076_ = _01451_ | _02097_;
	assign _02077_ = _02076_ | \mchip.index [8];
	assign _02078_ = \mchip.index [11] & ~_02077_;
	assign _02079_ = _02002_ | _04648_;
	assign _02080_ = _02079_ | _01986_;
	assign _02081_ = _01875_ & ~_02080_;
	assign _02082_ = _07654_ | \mchip.index [7];
	assign _02083_ = _02082_ | \mchip.index [8];
	assign _02084_ = _02083_ | \mchip.index [9];
	assign _02085_ = \mchip.index [11] & ~_02084_;
	assign _02087_ = _02696_ | \mchip.index [4];
	assign _02088_ = _02087_ | \mchip.index [5];
	assign _02089_ = _02088_ | _04648_;
	assign _02090_ = _02089_ | _07758_;
	assign _02091_ = _01986_ & ~_02090_;
	assign _02092_ = _07701_ | \mchip.index [6];
	assign _02093_ = _02092_ | \mchip.index [7];
	assign _02094_ = _02093_ | _04648_;
	assign _02095_ = _02094_ | \mchip.index [9];
	assign _02096_ = _02095_ | _01986_;
	assign _02099_ = _01875_ & ~_02096_;
	assign _02100_ = _01502_ | \mchip.index [6];
	assign _02101_ = _02100_ | _02097_;
	assign _02102_ = _02101_ | _04648_;
	assign _02103_ = _02102_ | \mchip.index [10];
	assign _02104_ = _01875_ & ~_02103_;
	assign _02105_ = _00348_ | \mchip.index [6];
	assign _02106_ = _02105_ | _02097_;
	assign _02107_ = _02106_ | \mchip.index [8];
	assign _02108_ = _02107_ | _07758_;
	assign _02110_ = \mchip.index [10] & ~_02108_;
	assign _02111_ = _00220_ | \mchip.index [8];
	assign _02112_ = _02111_ | _07758_;
	assign _02113_ = _02112_ | \mchip.index [10];
	assign _02114_ = _01875_ & ~_02113_;
	assign _02115_ = _01405_ | _02097_;
	assign _02116_ = _02115_ | \mchip.index [8];
	assign _02117_ = _02116_ | _07758_;
	assign _02118_ = _02117_ | \mchip.index [10];
	assign _02119_ = _01875_ & ~_02118_;
	assign _02121_ = _07648_ | _01098_;
	assign _02122_ = _02121_ | _02984_;
	assign _02123_ = _02122_ | _02097_;
	assign _02124_ = _02123_ | \mchip.index [8];
	assign _02125_ = _02124_ | \mchip.index [9];
	assign _02126_ = \mchip.index [11] & ~_02125_;
	assign _02127_ = _01383_ | \mchip.index [7];
	assign _02128_ = _02127_ | _04648_;
	assign _02129_ = _02128_ | _07758_;
	assign _02130_ = _02129_ | _01986_;
	assign _02132_ = _01875_ & ~_02130_;
	assign _02133_ = _00607_ | \mchip.index [6];
	assign _02134_ = _02133_ | _02097_;
	assign _02135_ = _02134_ | \mchip.index [8];
	assign _02136_ = _02135_ | \mchip.index [9];
	assign _02137_ = \mchip.index [11] & ~_02136_;
	assign _02138_ = _07774_ | \mchip.index [7];
	assign _02139_ = _02138_ | \mchip.index [8];
	assign _02140_ = _02139_ | _07758_;
	assign _02141_ = \mchip.index [10] & ~_02140_;
	assign _02143_ = _01540_ | \mchip.index [6];
	assign _02144_ = _02143_ | \mchip.index [7];
	assign _02145_ = _02144_ | _07758_;
	assign _02146_ = \mchip.index [11] & ~_02145_;
	assign _02147_ = _02101_ | \mchip.index [8];
	assign _02148_ = \mchip.index [10] & ~_02147_;
	assign _02149_ = _01166_ | \mchip.index [6];
	assign _02150_ = _02149_ | \mchip.index [7];
	assign _02151_ = _02150_ | _01986_;
	assign _02152_ = \mchip.index [11] & ~_02151_;
	assign _02154_ = _01749_ | _04648_;
	assign _02155_ = _02154_ | \mchip.index [9];
	assign _02156_ = \mchip.index [10] & ~_02155_;
	assign _02157_ = _01153_ | \mchip.index [6];
	assign _02158_ = _02157_ | _02097_;
	assign _02159_ = _02158_ | \mchip.index [8];
	assign _02160_ = _07758_ & ~_02159_;
	assign _02161_ = _00255_ | \mchip.index [6];
	assign _02162_ = _02161_ | \mchip.index [7];
	assign _02163_ = _02162_ | _04648_;
	assign _02165_ = _02163_ | \mchip.index [9];
	assign _02166_ = \mchip.index [11] & ~_02165_;
	assign _02167_ = _02088_ | _02984_;
	assign _02168_ = _02167_ | _07758_;
	assign _02169_ = _02168_ | \mchip.index [10];
	assign _02170_ = _01875_ & ~_02169_;
	assign _02171_ = _01383_ | \mchip.index [8];
	assign _02172_ = _02171_ | \mchip.index [9];
	assign _02173_ = _02172_ | \mchip.index [10];
	assign _02174_ = _01875_ & ~_02173_;
	assign _02176_ = _00566_ | \mchip.index [6];
	assign _02177_ = _02176_ | _02097_;
	assign _02178_ = _02177_ | _04648_;
	assign _02179_ = _02178_ | _07758_;
	assign _02180_ = _01986_ & ~_02179_;
	assign _02181_ = _02696_ | \mchip.index [6];
	assign _02182_ = _02181_ | _02097_;
	assign _02183_ = _02182_ | _04648_;
	assign _02184_ = _02183_ | \mchip.index [10];
	assign _02185_ = \mchip.index [11] & ~_02184_;
	assign _02187_ = _01104_ | _02097_;
	assign _02188_ = _02187_ | \mchip.index [8];
	assign _02189_ = _02188_ | _07758_;
	assign _02190_ = \mchip.index [11] & ~_02189_;
	assign _02191_ = _00209_ | _01098_;
	assign _02192_ = _02191_ | \mchip.index [6];
	assign _02193_ = _02192_ | \mchip.index [7];
	assign _02194_ = _02193_ | \mchip.index [9];
	assign _02195_ = \mchip.index [11] & ~_02194_;
	assign _02196_ = _02195_ | _02190_;
	assign _02198_ = _02196_ | _02185_;
	assign _02199_ = _02198_ | _02180_;
	assign _02200_ = _02199_ | _02174_;
	assign _02201_ = _02200_ | _02170_;
	assign _02202_ = _02201_ | _02166_;
	assign _02203_ = _02202_ | _02160_;
	assign _02204_ = _02203_ | _02156_;
	assign _02205_ = _02204_ | _02152_;
	assign _02206_ = _02205_ | _02148_;
	assign _02207_ = _02206_ | _02146_;
	assign _02210_ = _02207_ | _02141_;
	assign _02211_ = _02210_ | _02137_;
	assign _02212_ = _02211_ | _02132_;
	assign _02213_ = _02212_ | _02126_;
	assign _02214_ = _02213_ | _02119_;
	assign _02215_ = _02214_ | _02114_;
	assign _02216_ = _02215_ | _02110_;
	assign _02217_ = _02216_ | _02104_;
	assign _02218_ = _02217_ | _02099_;
	assign _02219_ = _02218_ | _02091_;
	assign _02221_ = _02219_ | _02085_;
	assign _02222_ = _02221_ | _02081_;
	assign _02223_ = _02222_ | _02078_;
	assign _02224_ = _02223_ | _02074_;
	assign _02225_ = _02224_ | _02071_;
	assign _02226_ = _02225_ | _02068_;
	assign _02227_ = _02226_ | _02063_;
	assign _02228_ = _02227_ | _02061_;
	assign _02229_ = _02228_ | _02056_;
	assign _02230_ = _02229_ | _02049_;
	assign _02232_ = _02230_ | _02043_;
	assign _02233_ = _02232_ | _02038_;
	assign _02234_ = _02233_ | _02033_;
	assign _02235_ = _02234_ | _02028_;
	assign _02236_ = _02235_ | _02024_;
	assign _02237_ = _02236_ | _02019_;
	assign _02238_ = _02237_ | _02014_;
	assign _02239_ = _02238_ | _02010_;
	assign _02240_ = _02239_ | _02005_;
	assign _02241_ = _02240_ | _02001_;
	assign _02243_ = _02241_ | _01999_;
	assign _02244_ = _02243_ | _01994_;
	assign _02245_ = _02244_ | _01989_;
	assign _02246_ = _02245_ | _01982_;
	assign _02247_ = _02246_ | _01977_;
	assign _02248_ = _02247_ | _01974_;
	assign _02249_ = _02248_ | _01969_;
	assign _02250_ = _02249_ | _01963_;
	assign _02251_ = _02250_ | _01955_;
	assign _02252_ = _02251_ | _01948_;
	assign _02254_ = _02252_ | _01941_;
	assign _02255_ = _02254_ | _01936_;
	assign _02256_ = _02255_ | _01932_;
	assign _02257_ = _02256_ | _01928_;
	assign _02258_ = _02257_ | _01923_;
	assign _02259_ = _02258_ | _01917_;
	assign _02260_ = _02259_ | _01913_;
	assign _02261_ = _02260_ | _01907_;
	assign _02262_ = _02261_ | _01903_;
	assign _02263_ = _02262_ | _01897_;
	assign _02265_ = _02263_ | _01896_;
	assign _02266_ = _02265_ | _01891_;
	assign _02267_ = _02266_ | _01888_;
	assign _02268_ = _02267_ | _01884_;
	assign _02269_ = _02268_ | _01880_;
	assign _02270_ = _02269_ | _01873_;
	assign _02271_ = _02270_ | _01868_;
	assign _02272_ = _02271_ | _01862_;
	assign _02273_ = _02272_ | _01857_;
	assign _02274_ = _02273_ | _01855_;
	assign _02276_ = _02274_ | _01847_;
	assign _02277_ = _02276_ | _01845_;
	assign _02278_ = _02277_ | _01844_;
	assign _02279_ = _02278_ | _01838_;
	assign _02280_ = _02279_ | _01832_;
	assign _02281_ = _02280_ | _01827_;
	assign _02282_ = _02281_ | _01822_;
	assign _02283_ = _02282_ | _01817_;
	assign _02284_ = _02283_ | _01813_;
	assign _02285_ = _02284_ | _01810_;
	assign _02287_ = _02285_ | _01804_;
	assign _02288_ = _02287_ | _01801_;
	assign _02289_ = _02288_ | _01795_;
	assign _02290_ = _02289_ | _01790_;
	assign _02291_ = _02290_ | _01786_;
	assign _02292_ = _02291_ | _01782_;
	assign _02293_ = _02292_ | _01779_;
	assign _02294_ = _02293_ | _01773_;
	assign _02295_ = _02294_ | _01770_;
	assign _02296_ = _02295_ | _01763_;
	assign _02298_ = _02296_ | _01759_;
	assign _02299_ = _02298_ | _01752_;
	assign _02300_ = _02299_ | _01747_;
	assign _02301_ = _02300_ | _01743_;
	assign _02302_ = _02301_ | _01736_;
	assign _02303_ = _02302_ | _01732_;
	assign _02304_ = _02303_ | _01726_;
	assign _02305_ = _02304_ | _01721_;
	assign _02306_ = _02305_ | _01715_;
	assign _02307_ = _02306_ | _01707_;
	assign _02309_ = _02307_ | _01705_;
	assign _02310_ = _02309_ | _01701_;
	assign _02311_ = _02310_ | _01696_;
	assign _02312_ = _02311_ | _01693_;
	assign _02313_ = _02312_ | _01691_;
	assign _02314_ = _02313_ | _01688_;
	assign _02315_ = _02314_ | _01684_;
	assign _02316_ = _02315_ | _01679_;
	assign _02317_ = _02316_ | _01673_;
	assign _02318_ = _02317_ | _01669_;
	assign _02321_ = _02318_ | _01663_;
	assign _02322_ = _02321_ | _01660_;
	assign _02323_ = _02322_ | _01655_;
	assign _02324_ = _02323_ | _01649_;
	assign _02325_ = _02324_ | _01646_;
	assign _02326_ = _02325_ | _01639_;
	assign _02327_ = _02326_ | _01634_;
	assign _02328_ = _02327_ | _01628_;
	assign _02329_ = _02328_ | _01624_;
	assign _02330_ = _02329_ | _01617_;
	assign _02332_ = _02330_ | _01612_;
	assign _02333_ = _02332_ | _01606_;
	assign _02334_ = _02333_ | _01602_;
	assign _02335_ = _02334_ | _01597_;
	assign _02336_ = _02335_ | _01592_;
	assign _02337_ = _02336_ | _01590_;
	assign _02338_ = _02337_ | _01585_;
	assign _02339_ = _02338_ | _01580_;
	assign _02340_ = _02339_ | _01578_;
	assign _02341_ = _02340_ | _01572_;
	assign _02343_ = _02341_ | _01568_;
	assign _02344_ = _02343_ | _01560_;
	assign _02345_ = _02344_ | _01557_;
	assign _02346_ = _02345_ | _01550_;
	assign _02347_ = _02346_ | _01546_;
	assign _02348_ = _02347_ | _01539_;
	assign _02349_ = _02348_ | _01533_;
	assign _02350_ = _02349_ | _01526_;
	assign _02351_ = _02350_ | _01522_;
	assign _02352_ = _02351_ | _01519_;
	assign _02354_ = _02352_ | _01514_;
	assign _02355_ = _02354_ | _01507_;
	assign _02356_ = _02355_ | _01500_;
	assign _02357_ = _02356_ | _01496_;
	assign _02358_ = _02357_ | _01489_;
	assign _02359_ = _02358_ | _01484_;
	assign _02360_ = _02359_ | _01480_;
	assign _02361_ = _02360_ | _01475_;
	assign _02362_ = _02361_ | _01471_;
	assign _02363_ = _02362_ | _01467_;
	assign _02365_ = _02363_ | _01460_;
	assign _02366_ = _02365_ | _01455_;
	assign _02367_ = _02366_ | _01450_;
	assign _02368_ = _02367_ | _01446_;
	assign _02369_ = _02368_ | _01441_;
	assign _02370_ = _02369_ | _01437_;
	assign _02371_ = _02370_ | _01434_;
	assign _02372_ = _02371_ | _01426_;
	assign _02373_ = _02372_ | _01421_;
	assign _02374_ = _02373_ | _01416_;
	assign _02376_ = _02374_ | _01414_;
	assign _02377_ = _02376_ | _01411_;
	assign _02378_ = _02377_ | _01404_;
	assign _02379_ = _02378_ | _01402_;
	assign _02380_ = _02379_ | _01396_;
	assign _02381_ = _02380_ | _01393_;
	assign _02382_ = _02381_ | _01388_;
	assign _02383_ = _02382_ | _01382_;
	assign _02384_ = _02383_ | _01378_;
	assign _02385_ = _02384_ | _01372_;
	assign _02387_ = _02385_ | _01368_;
	assign _02388_ = _02387_ | _01363_;
	assign _02389_ = _02388_ | _01358_;
	assign _02390_ = _02389_ | _01352_;
	assign _02391_ = _02390_ | _01346_;
	assign _02392_ = _02391_ | _01340_;
	assign _02393_ = _02392_ | _01335_;
	assign _02394_ = _02393_ | _01331_;
	assign _02395_ = _02394_ | _01323_;
	assign _02396_ = _02395_ | _01315_;
	assign _02398_ = _02396_ | _01310_;
	assign _02399_ = _02398_ | _01303_;
	assign _02400_ = _02399_ | _01296_;
	assign _02401_ = _02400_ | _01289_;
	assign _02402_ = _02401_ | _01285_;
	assign _02403_ = _02402_ | _01281_;
	assign _02404_ = _02403_ | _01275_;
	assign _02405_ = _02404_ | _01271_;
	assign _02406_ = _02405_ | _01267_;
	assign _02407_ = _02406_ | _01261_;
	assign _02409_ = _02407_ | _01258_;
	assign _02410_ = _02409_ | _01252_;
	assign _02411_ = _02410_ | _01248_;
	assign _02412_ = _02411_ | _01241_;
	assign _02413_ = _02412_ | _01236_;
	assign _02414_ = _02413_ | _01229_;
	assign _02415_ = _02414_ | _01224_;
	assign _02416_ = _02415_ | _01217_;
	assign _02417_ = _02416_ | _01213_;
	assign _02418_ = _02417_ | _01206_;
	assign _02420_ = _02418_ | _01201_;
	assign _02421_ = _02420_ | _01195_;
	assign _02422_ = _02421_ | _01188_;
	assign _02423_ = _02422_ | _01183_;
	assign _02424_ = _02423_ | _01177_;
	assign _02425_ = _02424_ | _01171_;
	assign _02426_ = _02425_ | _01164_;
	assign _02427_ = _02426_ | _01158_;
	assign _02428_ = _02427_ | _01151_;
	assign _02429_ = _02428_ | _01146_;
	assign _02432_ = _02429_ | _01141_;
	assign _02433_ = _02432_ | _01137_;
	assign _02434_ = _02433_ | _01130_;
	assign _02435_ = _02434_ | _01125_;
	assign _02436_ = _02435_ | _01119_;
	assign _02437_ = _02436_ | _01116_;
	assign _02438_ = _02437_ | _01109_;
	assign \mchip.val [4] = _02438_ | _01103_;
	assign _02439_ = _00381_ | \mchip.index [6];
	assign _02440_ = _02439_ | \mchip.index [7];
	assign _02442_ = _02440_ | \mchip.index [8];
	assign _02443_ = _07758_ & ~_02442_;
	assign _02444_ = _00856_ | \mchip.index [6];
	assign _02445_ = _02444_ | _02097_;
	assign _02446_ = _02445_ | _04648_;
	assign _02447_ = _02446_ | \mchip.index [9];
	assign _02448_ = \mchip.index [10] & ~_02447_;
	assign _02449_ = _01461_ | \mchip.index [7];
	assign _02450_ = _02449_ | \mchip.index [8];
	assign _02451_ = \mchip.index [10] & ~_02450_;
	assign _02453_ = _01657_ | \mchip.index [8];
	assign _02454_ = \mchip.index [9] & ~_02453_;
	assign _02455_ = _00324_ | \mchip.index [7];
	assign _02456_ = _02455_ | \mchip.index [8];
	assign _02457_ = \mchip.index [11] & ~_02456_;
	assign _02458_ = _01190_ | _02097_;
	assign _02459_ = _02458_ | _04648_;
	assign _02460_ = \mchip.index [11] & ~_02459_;
	assign _02461_ = _06090_ | _02984_;
	assign _02462_ = _02461_ | \mchip.index [7];
	assign _02464_ = _02462_ | _04648_;
	assign _02465_ = _02464_ | \mchip.index [10];
	assign _02466_ = _01875_ & ~_02465_;
	assign _02467_ = _00366_ | _05424_;
	assign _02468_ = \mchip.index [6] & ~_02467_;
	assign _02469_ = _07864_ | \mchip.index [7];
	assign _02470_ = _02469_ | \mchip.index [8];
	assign _02471_ = \mchip.index [10] & ~_02470_;
	assign _02472_ = _07677_ | \mchip.index [7];
	assign _02473_ = _02472_ | \mchip.index [8];
	assign _02475_ = _02473_ | \mchip.index [9];
	assign _02476_ = \mchip.index [11] & ~_02475_;
	assign _02477_ = _01000_ | _02984_;
	assign _02478_ = _02477_ | \mchip.index [7];
	assign _02479_ = _02478_ | _04648_;
	assign _02480_ = _07758_ & ~_02479_;
	assign _02481_ = _01635_ | _02097_;
	assign _02482_ = _02481_ | _04648_;
	assign _02483_ = \mchip.index [9] & ~_02482_;
	assign _02484_ = _02483_ & ~\mchip.index [11];
	assign _02486_ = _07843_ | _02984_;
	assign _02487_ = _02486_ | _02097_;
	assign _02488_ = _02487_ | \mchip.index [8];
	assign _02489_ = _02488_ | _07758_;
	assign _02490_ = _01986_ & ~_02489_;
	assign _02491_ = \mchip.index [9] & ~_01789_;
	assign _02492_ = _01574_ | _04648_;
	assign _02493_ = _02492_ | \mchip.index [9];
	assign _02494_ = _01986_ & ~_02493_;
	assign _02495_ = _03240_ | _02984_;
	assign _02497_ = _02495_ | \mchip.index [8];
	assign _02498_ = _02497_ | \mchip.index [10];
	assign _02499_ = _01875_ & ~_02498_;
	assign _02500_ = _01316_ | \mchip.index [6];
	assign _02501_ = _02500_ | _02097_;
	assign _02502_ = _02501_ | _04648_;
	assign _02503_ = _02502_ | _07758_;
	assign _02504_ = _01875_ & ~_02503_;
	assign _02505_ = _07588_ | \mchip.index [6];
	assign _02506_ = _02505_ | \mchip.index [8];
	assign _02508_ = _02506_ | \mchip.index [9];
	assign _02509_ = \mchip.index [11] & ~_02508_;
	assign _02510_ = _01842_ | \mchip.index [5];
	assign _02511_ = _02510_ | _02984_;
	assign _02512_ = _02511_ | _02097_;
	assign _02513_ = _02512_ | \mchip.index [8];
	assign _02514_ = _02513_ | \mchip.index [9];
	assign _02515_ = \mchip.index [10] & ~_02514_;
	assign _02516_ = _01189_ | _05424_;
	assign _02517_ = _02984_ & ~_02516_;
	assign _02519_ = _02220_ | \mchip.index [7];
	assign _02520_ = _02519_ | _04648_;
	assign _02521_ = _02520_ | \mchip.index [9];
	assign _02522_ = _01875_ & ~_02521_;
	assign _02523_ = _01477_ | _02097_;
	assign _02524_ = \mchip.index [10] & ~_02523_;
	assign _02525_ = _01304_ | _02984_;
	assign _02526_ = _02525_ | _02097_;
	assign _02527_ = _02526_ | \mchip.index [8];
	assign _02528_ = _02527_ | _07758_;
	assign _02530_ = \mchip.index [10] & ~_02528_;
	assign _02531_ = _01502_ | \mchip.index [7];
	assign _02532_ = _02531_ | _04648_;
	assign _02533_ = _02532_ | \mchip.index [9];
	assign _02534_ = _01986_ & ~_02533_;
	assign _02535_ = _01505_ | _07758_;
	assign _02536_ = \mchip.index [10] & ~_02535_;
	assign _02537_ = _01198_ | _04648_;
	assign _02538_ = _02537_ | \mchip.index [9];
	assign _02539_ = _01986_ & ~_02538_;
	assign _02542_ = _04871_ | _02984_;
	assign _02543_ = _02542_ | \mchip.index [7];
	assign _02544_ = _02543_ | _04648_;
	assign _02545_ = _02544_ | _07758_;
	assign _02546_ = _01986_ & ~_02545_;
	assign _02547_ = _01477_ | _04648_;
	assign _02548_ = _07758_ & ~_02547_;
	assign _02549_ = _01249_ | \mchip.index [7];
	assign _02550_ = _02549_ | \mchip.index [9];
	assign _02551_ = _01875_ & ~_02550_;
	assign _02553_ = _00879_ | \mchip.index [5];
	assign _02554_ = _02553_ | \mchip.index [6];
	assign _02555_ = _02554_ | _02097_;
	assign _02556_ = _02555_ | \mchip.index [8];
	assign _02557_ = _02556_ | \mchip.index [9];
	assign _02558_ = \mchip.index [10] & ~_02557_;
	assign _02559_ = _02094_ | _07758_;
	assign _02560_ = _01875_ & ~_02559_;
	assign _02561_ = _03206_ | _07758_;
	assign _02562_ = _02561_ | \mchip.index [10];
	assign _02564_ = \mchip.index [11] & ~_02562_;
	assign _02565_ = _04871_ | _05424_;
	assign _02566_ = _02565_ | _02984_;
	assign _02567_ = _02566_ | _07758_;
	assign _02568_ = \mchip.index [10] & ~_02567_;
	assign _02569_ = _00593_ | _02097_;
	assign _02570_ = _02569_ | _04648_;
	assign _02571_ = _02570_ | \mchip.index [9];
	assign _02572_ = _01986_ & ~_02571_;
	assign _02573_ = _00856_ | \mchip.index [5];
	assign _02575_ = _02573_ | _02984_;
	assign _02576_ = _02575_ | \mchip.index [7];
	assign _02577_ = _02576_ | _04648_;
	assign _02578_ = _02577_ | _07758_;
	assign _02579_ = \mchip.index [10] & ~_02578_;
	assign _02580_ = _04205_ | \mchip.index [6];
	assign _02581_ = _02580_ | _02097_;
	assign _02582_ = _02581_ | \mchip.index [8];
	assign _02583_ = _02582_ | \mchip.index [9];
	assign _02584_ = _02583_ | _01986_;
	assign _02586_ = _01875_ & ~_02584_;
	assign _02587_ = _01680_ | _04648_;
	assign _02588_ = _07758_ & ~_02587_;
	assign _02589_ = _07311_ | \mchip.index [7];
	assign _02590_ = _02589_ | _04648_;
	assign _02591_ = _02590_ | \mchip.index [9];
	assign _02592_ = _01986_ & ~_02591_;
	assign _02593_ = _00879_ | \mchip.index [6];
	assign _02594_ = _02593_ | _02097_;
	assign _02595_ = _02594_ | _04648_;
	assign _02597_ = _02595_ | _07758_;
	assign _02598_ = _02597_ | _01986_;
	assign _02599_ = _01875_ & ~_02598_;
	assign _02600_ = _07798_ | \mchip.index [5];
	assign _02601_ = _02600_ | _02984_;
	assign _02602_ = _02601_ | _02097_;
	assign _02603_ = _02602_ | _04648_;
	assign _02604_ = _02603_ | \mchip.index [9];
	assign _02605_ = _01875_ & ~_02604_;
	assign _02606_ = _01848_ | \mchip.index [6];
	assign _02608_ = _02606_ | \mchip.index [7];
	assign _02609_ = _02608_ | _04648_;
	assign _02610_ = _02609_ | \mchip.index [9];
	assign _02611_ = \mchip.index [10] & ~_02610_;
	assign _02612_ = _01586_ | _02097_;
	assign _02613_ = _02612_ | _04648_;
	assign _02614_ = _02613_ | _01986_;
	assign _02615_ = _01875_ & ~_02614_;
	assign _02616_ = _01153_ | _04648_;
	assign _02617_ = _02616_ | \mchip.index [9];
	assign _02619_ = \mchip.index [11] & ~_02617_;
	assign _02620_ = _00684_ | \mchip.index [6];
	assign _02621_ = _02620_ | \mchip.index [7];
	assign _02622_ = _02621_ | \mchip.index [8];
	assign _02623_ = \mchip.index [11] & ~_02622_;
	assign _02624_ = \mchip.index [11] & ~_02570_;
	assign _02625_ = _01000_ | \mchip.index [5];
	assign _02626_ = _02625_ | \mchip.index [6];
	assign _02627_ = _02626_ | _02097_;
	assign _02628_ = _02627_ | _01986_;
	assign _02630_ = \mchip.index [11] & ~_02628_;
	assign _02631_ = _00299_ | _02097_;
	assign _02632_ = _02631_ | \mchip.index [9];
	assign _02633_ = _02632_ | \mchip.index [10];
	assign _02634_ = _01875_ & ~_02633_;
	assign _02635_ = _01824_ | _02097_;
	assign _02636_ = _02635_ | \mchip.index [8];
	assign _02637_ = _02636_ | \mchip.index [9];
	assign _02638_ = \mchip.index [10] & ~_02637_;
	assign _02639_ = _01390_ | \mchip.index [9];
	assign _02641_ = _02639_ | \mchip.index [10];
	assign _02642_ = _01875_ & ~_02641_;
	assign _02643_ = ~(_02729_ & \mchip.index [9]);
	assign _02644_ = \mchip.index [11] & ~_02643_;
	assign _02645_ = \mchip.index [11] & ~_01906_;
	assign _02646_ = _00884_ | _02097_;
	assign _02647_ = _02646_ | \mchip.index [9];
	assign _02648_ = _01875_ & ~_02647_;
	assign _02649_ = _07773_ | \mchip.index [5];
	assign _02650_ = _02649_ | \mchip.index [6];
	assign _02653_ = _02650_ | _07758_;
	assign _02654_ = \mchip.index [11] & ~_02653_;
	assign _02655_ = _01196_ | _05424_;
	assign _02656_ = _02655_ | \mchip.index [6];
	assign _02657_ = _02097_ & ~_02656_;
	assign _02658_ = _02029_ | _02097_;
	assign _02659_ = _02658_ | \mchip.index [9];
	assign _02660_ = \mchip.index [10] & ~_02659_;
	assign _02661_ = _01823_ | \mchip.index [5];
	assign _02662_ = _02661_ | \mchip.index [7];
	assign _02664_ = _02662_ | _04648_;
	assign _02665_ = _02664_ | _07758_;
	assign _02666_ = _02665_ | _01986_;
	assign _02667_ = _01875_ & ~_02666_;
	assign _02668_ = _05070_ | _02097_;
	assign _02669_ = _02668_ | _04648_;
	assign _02670_ = _02669_ | _07758_;
	assign _02671_ = _01986_ & ~_02670_;
	assign _02672_ = _01230_ | _02984_;
	assign _02673_ = _02672_ | \mchip.index [8];
	assign _02675_ = _02673_ | _07758_;
	assign _02676_ = \mchip.index [11] & ~_02675_;
	assign _02677_ = _01428_ | \mchip.index [6];
	assign _02678_ = _02677_ | _02097_;
	assign _02679_ = _02678_ | _04648_;
	assign _02680_ = \mchip.index [11] & ~_02679_;
	assign _02681_ = _01547_ | \mchip.index [6];
	assign _02682_ = _02681_ | _04648_;
	assign _02683_ = _01986_ & ~_02682_;
	assign _02684_ = _01600_ | _07758_;
	assign _02686_ = _02684_ | \mchip.index [10];
	assign _02687_ = \mchip.index [11] & ~_02686_;
	assign _02688_ = _01262_ | _04648_;
	assign _02689_ = _02688_ | \mchip.index [9];
	assign _02690_ = \mchip.index [10] & ~_02689_;
	assign _02691_ = _01255_ | \mchip.index [7];
	assign _02692_ = _02691_ | \mchip.index [8];
	assign _02693_ = _01875_ & ~_02692_;
	assign _02694_ = _04882_ | \mchip.index [6];
	assign _02695_ = _02694_ | \mchip.index [7];
	assign _02697_ = _02695_ | \mchip.index [8];
	assign _02698_ = _07758_ & ~_02697_;
	assign _02699_ = _00345_ | \mchip.index [6];
	assign _02700_ = _02699_ | _02097_;
	assign _02701_ = _02700_ | \mchip.index [8];
	assign _02702_ = _02701_ | \mchip.index [9];
	assign _02703_ = _01875_ & ~_02702_;
	assign _02704_ = _00380_ | \mchip.index [7];
	assign _02705_ = _02704_ | \mchip.index [8];
	assign _02706_ = _02705_ | \mchip.index [10];
	assign _02708_ = _01875_ & ~_02706_;
	assign _02709_ = _00353_ | _02097_;
	assign _02710_ = _02709_ | \mchip.index [9];
	assign _02711_ = _02710_ | \mchip.index [10];
	assign _02712_ = _01875_ & ~_02711_;
	assign _02713_ = _00856_ | _02984_;
	assign _02714_ = _02713_ | _02097_;
	assign _02715_ = _02714_ | \mchip.index [8];
	assign _02716_ = _02715_ | \mchip.index [9];
	assign _02717_ = \mchip.index [10] & ~_02716_;
	assign _02719_ = _01343_ | _02984_;
	assign _02720_ = _02719_ | _04648_;
	assign _02721_ = _02720_ | \mchip.index [9];
	assign _02722_ = _02721_ | \mchip.index [10];
	assign _02723_ = _01875_ & ~_02722_;
	assign _02724_ = _01147_ | _02984_;
	assign _02725_ = _02724_ | \mchip.index [7];
	assign _02726_ = _02725_ | \mchip.index [10];
	assign _02727_ = \mchip.index [11] & ~_02726_;
	assign _02728_ = _01551_ | \mchip.index [6];
	assign _02730_ = _02728_ | \mchip.index [7];
	assign _02731_ = _02730_ | _07758_;
	assign _02732_ = \mchip.index [11] & ~_02731_;
	assign _02733_ = _07310_ | \mchip.index [8];
	assign _02734_ = _02733_ | _07758_;
	assign _02735_ = _02734_ | \mchip.index [10];
	assign _02736_ = _01875_ & ~_02735_;
	assign _02737_ = _02719_ | _02097_;
	assign _02738_ = _02737_ | _01986_;
	assign _02739_ = \mchip.index [11] & ~_02738_;
	assign _02741_ = _01250_ | _04648_;
	assign _02742_ = \mchip.index [10] & ~_02741_;
	assign _02743_ = _01908_ | \mchip.index [6];
	assign _02744_ = _02743_ | \mchip.index [7];
	assign _02745_ = _02744_ | _04648_;
	assign _02746_ = _02745_ | \mchip.index [9];
	assign _02747_ = _01986_ & ~_02746_;
	assign _02748_ = _01333_ | \mchip.index [8];
	assign _02749_ = \mchip.index [10] & ~_02748_;
	assign _02750_ = _01892_ | _02984_;
	assign _02752_ = _02750_ | _02097_;
	assign _02753_ = _02752_ | \mchip.index [8];
	assign _02754_ = _07758_ & ~_02753_;
	assign _02755_ = _01892_ | \mchip.index [7];
	assign _02756_ = _02755_ | _07758_;
	assign _02757_ = _01875_ & ~_02756_;
	assign _02758_ = _01461_ | \mchip.index [6];
	assign _02759_ = _02758_ | _07758_;
	assign _02760_ = _02759_ | \mchip.index [10];
	assign _02761_ = _01875_ & ~_02760_;
	assign _02764_ = _01387_ | \mchip.index [8];
	assign _02765_ = _02764_ | \mchip.index [9];
	assign _02766_ = \mchip.index [10] & ~_02765_;
	assign _02767_ = _02694_ | _02097_;
	assign _02768_ = _02767_ | _04648_;
	assign _02769_ = \mchip.index [10] & ~_02768_;
	assign _02770_ = _02209_ | _02097_;
	assign _02771_ = _02770_ | _07758_;
	assign _02772_ = _02771_ | \mchip.index [10];
	assign _02773_ = \mchip.index [11] & ~_02772_;
	assign _02775_ = _00837_ | _02984_;
	assign _02776_ = _02775_ | \mchip.index [7];
	assign _02777_ = _02776_ | _04648_;
	assign _02778_ = _02777_ | _07758_;
	assign _02779_ = _01875_ & ~_02778_;
	assign _02780_ = _04482_ | _05424_;
	assign _02781_ = _02097_ & ~_02780_;
	assign _02782_ = _01774_ | \mchip.index [7];
	assign _02783_ = _02782_ | _04648_;
	assign _02784_ = _07758_ & ~_02783_;
	assign _02786_ = _00429_ | \mchip.index [6];
	assign _02787_ = _02786_ | \mchip.index [7];
	assign _02788_ = _02787_ | \mchip.index [9];
	assign _02789_ = _01875_ & ~_02788_;
	assign _02790_ = _00559_ | \mchip.index [5];
	assign _02791_ = _02790_ | _02984_;
	assign _02792_ = _02791_ | \mchip.index [7];
	assign _02793_ = _02792_ | _01986_;
	assign _02794_ = \mchip.index [11] & ~_02793_;
	assign _02795_ = _01501_ | _02984_;
	assign _02797_ = _02795_ | _02097_;
	assign _02798_ = _02797_ | \mchip.index [9];
	assign _02799_ = \mchip.index [11] & ~_02798_;
	assign _02800_ = _00380_ | \mchip.index [6];
	assign _02801_ = _02800_ | \mchip.index [8];
	assign _02802_ = _02801_ | _07758_;
	assign _02803_ = _02802_ | \mchip.index [10];
	assign _02804_ = _01875_ & ~_02803_;
	assign _02805_ = _01796_ | \mchip.index [7];
	assign _02806_ = _02805_ | _04648_;
	assign _02808_ = _02806_ | \mchip.index [9];
	assign _02809_ = \mchip.index [10] & ~_02808_;
	assign _02810_ = _01904_ | \mchip.index [6];
	assign _02811_ = _02810_ | _02097_;
	assign _02812_ = _02811_ | \mchip.index [9];
	assign _02813_ = \mchip.index [10] & ~_02812_;
	assign _02814_ = _01802_ | \mchip.index [9];
	assign _02815_ = \mchip.index [11] & ~_02814_;
	assign _02816_ = _01106_ | _07758_;
	assign _02817_ = \mchip.index [10] & ~_02816_;
	assign _02819_ = _01111_ | _05424_;
	assign _02820_ = _02819_ | _02097_;
	assign _02821_ = _02820_ | _07758_;
	assign _02822_ = _01875_ & ~_02821_;
	assign _02823_ = _01230_ | _02097_;
	assign _02824_ = _02823_ | \mchip.index [8];
	assign _02825_ = _02824_ | \mchip.index [9];
	assign _02826_ = _02825_ | \mchip.index [10];
	assign _02827_ = _01875_ & ~_02826_;
	assign _02828_ = _00351_ | _02097_;
	assign _02830_ = _02828_ | \mchip.index [8];
	assign _02831_ = _02830_ | _07758_;
	assign _02832_ = _02831_ | \mchip.index [10];
	assign _02833_ = \mchip.index [11] & ~_02832_;
	assign _02834_ = _01814_ | \mchip.index [9];
	assign _02835_ = \mchip.index [10] & ~_02834_;
	assign _02836_ = _01748_ | _02097_;
	assign _02837_ = _02836_ | _04648_;
	assign _02838_ = _02837_ | _07758_;
	assign _02839_ = _01986_ & ~_02838_;
	assign _02841_ = _05868_ | _05424_;
	assign _02842_ = _02841_ | _02984_;
	assign _02843_ = _02842_ | \mchip.index [7];
	assign _02844_ = _02843_ | _04648_;
	assign _02845_ = _01875_ & ~_02844_;
	assign _02846_ = _02087_ | _02984_;
	assign _02847_ = _02846_ | \mchip.index [7];
	assign _02848_ = _02847_ | _04648_;
	assign _02849_ = \mchip.index [10] & ~_02848_;
	assign _02850_ = _01476_ | _05424_;
	assign _02852_ = _02850_ | \mchip.index [7];
	assign _02853_ = _02852_ | _04648_;
	assign _02854_ = \mchip.index [11] & ~_02853_;
	assign _02855_ = _07675_ | \mchip.index [4];
	assign _02856_ = _02855_ | \mchip.index [6];
	assign _02857_ = _02856_ | \mchip.index [7];
	assign _02858_ = _02857_ | _07758_;
	assign _02859_ = _02858_ | \mchip.index [10];
	assign _02860_ = \mchip.index [11] & ~_02859_;
	assign _02861_ = _07773_ | \mchip.index [7];
	assign _02863_ = _02861_ | _07758_;
	assign _02864_ = _01986_ & ~_02863_;
	assign _02865_ = \mchip.index [10] & ~_02643_;
	assign _02866_ = _00406_ | _02097_;
	assign _02867_ = _02866_ | \mchip.index [8];
	assign _02868_ = \mchip.index [10] & ~_02867_;
	assign _02869_ = _03040_ | _02097_;
	assign _02870_ = _02869_ | \mchip.index [9];
	assign _02871_ = _02870_ | \mchip.index [10];
	assign _02872_ = _01875_ & ~_02871_;
	assign _02875_ = _00453_ | _02097_;
	assign _02876_ = _02875_ | _04648_;
	assign _02877_ = _02876_ | _07758_;
	assign _02878_ = _02877_ | _01986_;
	assign _02879_ = _01875_ & ~_02878_;
	assign _02880_ = _02088_ | _02097_;
	assign _02881_ = _02880_ | _04648_;
	assign _02882_ = _02881_ | _07758_;
	assign _02883_ = \mchip.index [10] & ~_02882_;
	assign _02884_ = _01290_ | \mchip.index [6];
	assign _02886_ = _02884_ | _02097_;
	assign _02887_ = _02886_ | \mchip.index [8];
	assign _02888_ = _02887_ | \mchip.index [9];
	assign _02889_ = _01986_ & ~_02888_;
	assign _02890_ = _07088_ | _05424_;
	assign _02891_ = _02890_ | _04648_;
	assign _02892_ = _02891_ | _07758_;
	assign _02893_ = _02892_ | _01986_;
	assign _02894_ = _01875_ & ~_02893_;
	assign _02895_ = _01943_ | \mchip.index [5];
	assign _02897_ = _02895_ | _02097_;
	assign _02898_ = _02897_ | _04648_;
	assign _02899_ = _02898_ | \mchip.index [10];
	assign _02900_ = _01875_ & ~_02899_;
	assign _02901_ = _01104_ | _04648_;
	assign _02902_ = _02901_ | \mchip.index [10];
	assign _02903_ = \mchip.index [11] & ~_02902_;
	assign _02904_ = _01607_ | _01986_;
	assign _02905_ = \mchip.index [11] & ~_02904_;
	assign _02906_ = _02856_ | _02097_;
	assign _02908_ = _02906_ | _04648_;
	assign _02909_ = _02908_ | \mchip.index [9];
	assign _02910_ = \mchip.index [10] & ~_02909_;
	assign _02911_ = _03029_ | \mchip.index [6];
	assign _02912_ = _02911_ | \mchip.index [7];
	assign _02913_ = _02912_ | \mchip.index [8];
	assign _02914_ = _02913_ | \mchip.index [9];
	assign _02915_ = \mchip.index [10] & ~_02914_;
	assign _02916_ = _01535_ | \mchip.index [8];
	assign _02917_ = _02916_ | _07758_;
	assign _02919_ = _02917_ | \mchip.index [10];
	assign _02920_ = _01875_ & ~_02919_;
	assign _02921_ = _01904_ | _04648_;
	assign _02922_ = _02921_ | _07758_;
	assign _02923_ = _02922_ | _01986_;
	assign _02924_ = _01875_ & ~_02923_;
	assign _02925_ = _02419_ | \mchip.index [5];
	assign _02926_ = _02925_ | \mchip.index [6];
	assign _02927_ = _02926_ | _02097_;
	assign _02928_ = _02927_ | _04648_;
	assign _02930_ = \mchip.index [11] & ~_02928_;
	assign _02931_ = _01376_ | \mchip.index [6];
	assign _02932_ = _02931_ | _02097_;
	assign _02933_ = _02932_ | _04648_;
	assign _02934_ = _02933_ | \mchip.index [9];
	assign _02935_ = \mchip.index [10] & ~_02934_;
	assign _02936_ = _07824_ | _05424_;
	assign _02937_ = _02097_ & ~_02936_;
	assign _02938_ = _01379_ | \mchip.index [8];
	assign _02939_ = _02938_ | \mchip.index [10];
	assign _02941_ = _01875_ & ~_02939_;
	assign _02942_ = _07671_ | _02984_;
	assign _02943_ = _02942_ | _02097_;
	assign _02944_ = _02943_ | _04648_;
	assign _02945_ = _02944_ | \mchip.index [10];
	assign _02946_ = \mchip.index [11] & ~_02945_;
	assign _02947_ = _01253_ | \mchip.index [6];
	assign _02948_ = _02947_ | \mchip.index [7];
	assign _02949_ = _02948_ | \mchip.index [9];
	assign _02950_ = \mchip.index [10] & ~_02949_;
	assign _02952_ = _02088_ | \mchip.index [6];
	assign _02953_ = _02952_ | \mchip.index [7];
	assign _02954_ = _02953_ | \mchip.index [10];
	assign _02955_ = \mchip.index [11] & ~_02954_;
	assign _02956_ = _02087_ | \mchip.index [6];
	assign _02957_ = _02956_ | _02097_;
	assign _02958_ = _02957_ | _04648_;
	assign _02959_ = \mchip.index [10] & ~_02958_;
	assign _02960_ = _05059_ | \mchip.index [5];
	assign _02961_ = _02960_ | _02984_;
	assign _02963_ = _02961_ | \mchip.index [7];
	assign _02964_ = _02963_ | _01986_;
	assign _02965_ = \mchip.index [11] & ~_02964_;
	assign _02966_ = _01231_ | \mchip.index [7];
	assign _02967_ = _02966_ | _07758_;
	assign _02968_ = _02967_ | _01986_;
	assign _02969_ = _01875_ & ~_02968_;
	assign _02970_ = _00469_ | _02984_;
	assign _02971_ = _02970_ | \mchip.index [7];
	assign _02972_ = _02971_ | _01986_;
	assign _02974_ = \mchip.index [11] & ~_02972_;
	assign _02975_ = _03240_ | \mchip.index [5];
	assign _02976_ = _02975_ | _02097_;
	assign _02977_ = _02976_ | \mchip.index [8];
	assign _02978_ = _02977_ | \mchip.index [9];
	assign _02979_ = _01875_ & ~_02978_;
	assign _02980_ = _01863_ | _02984_;
	assign _02981_ = _02980_ | \mchip.index [7];
	assign _02982_ = _02981_ | \mchip.index [9];
	assign _02983_ = \mchip.index [11] & ~_02982_;
	assign _02986_ = _02677_ | \mchip.index [7];
	assign _02987_ = _02986_ | _07758_;
	assign _02988_ = _01986_ & ~_02987_;
	assign _02989_ = _01461_ | \mchip.index [5];
	assign _02990_ = _02989_ | _02984_;
	assign _02991_ = _02990_ | \mchip.index [7];
	assign _02992_ = _02991_ | \mchip.index [8];
	assign _02993_ = _02992_ | \mchip.index [9];
	assign _02994_ = \mchip.index [11] & ~_02993_;
	assign _02995_ = _01347_ | _02984_;
	assign _02997_ = _02995_ | _02097_;
	assign _02998_ = _02997_ | \mchip.index [8];
	assign _02999_ = _02998_ | \mchip.index [9];
	assign _03000_ = _02999_ | \mchip.index [10];
	assign _03001_ = _01875_ & ~_03000_;
	assign _03002_ = _04882_ | _02097_;
	assign _03003_ = _03002_ | \mchip.index [9];
	assign _03004_ = \mchip.index [11] & ~_03003_;
	assign _03005_ = _00770_ | _04648_;
	assign _03006_ = _03005_ | _07758_;
	assign _03008_ = _03006_ | _01986_;
	assign _03009_ = _01875_ & ~_03008_;
	assign _03010_ = _00209_ | _05424_;
	assign _03011_ = _03010_ | _02097_;
	assign _03012_ = \mchip.index [11] & ~_03011_;
	assign _03013_ = _01398_ | _02097_;
	assign _03014_ = _03013_ | _01986_;
	assign _03015_ = \mchip.index [11] & ~_03014_;
	assign _03016_ = _01196_ | \mchip.index [5];
	assign _03017_ = _03016_ | _02984_;
	assign _03019_ = _03017_ | _02097_;
	assign _03020_ = _03019_ | _07758_;
	assign _03021_ = _03020_ | _01986_;
	assign _03022_ = _01875_ & ~_03021_;
	assign _03023_ = _01167_ | _01986_;
	assign _03024_ = \mchip.index [11] & ~_03023_;
	assign _03025_ = _01749_ | _07758_;
	assign _03026_ = _03025_ | \mchip.index [10];
	assign _03027_ = _01875_ & ~_03026_;
	assign _03028_ = _00816_ | \mchip.index [6];
	assign _03030_ = _03028_ | \mchip.index [7];
	assign _03031_ = _03030_ | \mchip.index [10];
	assign _03032_ = _01875_ & ~_03031_;
	assign _03033_ = _07773_ | _02097_;
	assign _03034_ = \mchip.index [11] & ~_03033_;
	assign _03035_ = _02191_ | _02984_;
	assign _03036_ = _03035_ | _04648_;
	assign _03037_ = _03036_ | \mchip.index [9];
	assign _03038_ = \mchip.index [11] & ~_03037_;
	assign _03039_ = _01681_ | \mchip.index [7];
	assign _03041_ = _03039_ | _07758_;
	assign _03042_ = \mchip.index [11] & ~_03041_;
	assign _03043_ = _01253_ | _02097_;
	assign _03044_ = _03043_ | \mchip.index [8];
	assign _03045_ = \mchip.index [11] & ~_03044_;
	assign _03046_ = _04471_ & ~_01875_;
	assign _03047_ = _00384_ | _05424_;
	assign _03048_ = _03047_ | _02097_;
	assign _03049_ = _03048_ | _04648_;
	assign _03050_ = \mchip.index [10] & ~_03049_;
	assign _03052_ = _04848_ | \mchip.index [8];
	assign _03053_ = _03052_ | \mchip.index [9];
	assign _03054_ = \mchip.index [10] & ~_03053_;
	assign _03055_ = _01558_ | \mchip.index [8];
	assign _03056_ = \mchip.index [9] & ~_03055_;
	assign _03057_ = _07399_ | _02984_;
	assign _03058_ = _03057_ | _02097_;
	assign _03059_ = _03058_ | _04648_;
	assign _03060_ = _03059_ | \mchip.index [9];
	assign _03061_ = _01875_ & ~_03060_;
	assign _03063_ = _01398_ | _02984_;
	assign _03064_ = _03063_ | _01986_;
	assign _03065_ = \mchip.index [11] & ~_03064_;
	assign _03066_ = _01253_ | \mchip.index [7];
	assign _03067_ = _03066_ | \mchip.index [9];
	assign _03068_ = \mchip.index [11] & ~_03067_;
	assign _03069_ = _01918_ | \mchip.index [7];
	assign _03070_ = _03069_ | _04648_;
	assign _03071_ = \mchip.index [9] & ~_03070_;
	assign _03072_ = _03071_ & ~\mchip.index [10];
	assign _03074_ = _01324_ | _02984_;
	assign _03075_ = _03074_ | _02097_;
	assign _03076_ = _03075_ | _04648_;
	assign _03077_ = _03076_ | _07758_;
	assign _03078_ = _03077_ | _01986_;
	assign _03079_ = _01875_ & ~_03078_;
	assign _03080_ = _01104_ | \mchip.index [6];
	assign _03081_ = _03080_ | _02097_;
	assign _03082_ = _07758_ & ~_03081_;
	assign _03083_ = _02149_ | _02097_;
	assign _03085_ = _03083_ | \mchip.index [8];
	assign _03086_ = _03085_ | \mchip.index [9];
	assign _03087_ = \mchip.index [11] & ~_03086_;
	assign _03088_ = _03080_ | \mchip.index [7];
	assign _03089_ = _04648_ & ~_03088_;
	assign _03090_ = _03089_ & ~_07758_;
	assign _03091_ = _06389_ | _02984_;
	assign _03092_ = _03091_ | _04648_;
	assign _03093_ = _03092_ | \mchip.index [9];
	assign _03094_ = \mchip.index [10] & ~_03093_;
	assign _03097_ = _01901_ | \mchip.index [8];
	assign _03098_ = _03097_ | _07758_;
	assign _03099_ = _01875_ & ~_03098_;
	assign _03100_ = _06346_ | \mchip.index [6];
	assign _03101_ = _03100_ | _02097_;
	assign _03102_ = _07758_ & ~_03101_;
	assign _03103_ = _01355_ | \mchip.index [9];
	assign _03104_ = _03103_ | \mchip.index [10];
	assign _03105_ = _01875_ & ~_03104_;
	assign _03106_ = _03080_ | _04648_;
	assign _03108_ = _03106_ | \mchip.index [9];
	assign _03109_ = \mchip.index [10] & ~_03108_;
	assign _03110_ = _01502_ | \mchip.index [5];
	assign _03111_ = _03110_ | \mchip.index [6];
	assign _03112_ = _03111_ | _02097_;
	assign _03113_ = _03112_ | _07758_;
	assign _03114_ = \mchip.index [11] & ~_03113_;
	assign _03115_ = _02840_ | \mchip.index [5];
	assign _03116_ = _03115_ | _02097_;
	assign _03117_ = _03116_ | _04648_;
	assign _03119_ = _03117_ | _07758_;
	assign _03120_ = _01986_ & ~_03119_;
	assign _03121_ = _00895_ | _07758_;
	assign _03122_ = _03121_ | \mchip.index [10];
	assign _03123_ = \mchip.index [11] & ~_03122_;
	assign _03124_ = _02842_ | _04648_;
	assign _03125_ = _03124_ | \mchip.index [10];
	assign _03126_ = _01875_ & ~_03125_;
	assign _03127_ = _02087_ | \mchip.index [7];
	assign _03128_ = _03127_ | _04648_;
	assign _03130_ = _03128_ | _07758_;
	assign _03131_ = _03130_ | _01986_;
	assign _03132_ = _01875_ & ~_03131_;
	assign _03133_ = _00000_ | \mchip.index [6];
	assign _03134_ = _03133_ | \mchip.index [8];
	assign _03135_ = _03134_ | \mchip.index [9];
	assign _03136_ = _03135_ | \mchip.index [10];
	assign _03137_ = _01875_ & ~_03136_;
	assign _03138_ = _01110_ | \mchip.index [6];
	assign _03139_ = _03138_ | _02097_;
	assign _03141_ = _03139_ | _04648_;
	assign _03142_ = \mchip.index [9] & ~_03141_;
	assign _03143_ = _04882_ | \mchip.index [7];
	assign _03144_ = _03143_ | _04648_;
	assign _03145_ = _03144_ | _07758_;
	assign _03146_ = _03145_ | _01986_;
	assign _03147_ = _01875_ & ~_03146_;
	assign _03148_ = _00785_ | \mchip.index [7];
	assign _03149_ = _03148_ | _04648_;
	assign _03150_ = _07758_ & ~_03149_;
	assign _03152_ = _00004_ | _04648_;
	assign _03153_ = _07758_ & ~_03152_;
	assign _03154_ = _01949_ | \mchip.index [5];
	assign _03155_ = _03154_ | _02984_;
	assign _03156_ = _03155_ | \mchip.index [8];
	assign _03157_ = _03156_ | _07758_;
	assign _03158_ = \mchip.index [10] & ~_03157_;
	assign _03159_ = _06589_ | \mchip.index [7];
	assign _03160_ = _03159_ | _04648_;
	assign _03161_ = _03160_ | \mchip.index [9];
	assign _03163_ = _03161_ | \mchip.index [10];
	assign _03164_ = _01875_ & ~_03163_;
	assign _03165_ = _00472_ | \mchip.index [6];
	assign _03166_ = _03165_ | _04648_;
	assign _03167_ = _03166_ | \mchip.index [9];
	assign _03168_ = \mchip.index [10] & ~_03167_;
	assign _03169_ = _00577_ | \mchip.index [8];
	assign _03170_ = _03169_ | \mchip.index [10];
	assign _03171_ = _01875_ & ~_03170_;
	assign _03172_ = _00471_ | \mchip.index [8];
	assign _03174_ = _03172_ | \mchip.index [9];
	assign _03175_ = \mchip.index [10] & ~_03174_;
	assign _03176_ = _02087_ | _02097_;
	assign _03177_ = _03176_ | _04648_;
	assign _03178_ = _03177_ | \mchip.index [9];
	assign _03179_ = _03178_ | \mchip.index [10];
	assign _03180_ = _01875_ & ~_03179_;
	assign _03181_ = _01914_ | \mchip.index [7];
	assign _03182_ = _03181_ | _04648_;
	assign _03183_ = _01986_ & ~_03182_;
	assign _03185_ = _01737_ | _02984_;
	assign _03186_ = _03185_ | \mchip.index [7];
	assign _03187_ = _03186_ | \mchip.index [8];
	assign _03188_ = _03187_ | \mchip.index [9];
	assign _03189_ = _01986_ & ~_03188_;
	assign _03190_ = _02177_ | \mchip.index [8];
	assign _03191_ = _03190_ | \mchip.index [9];
	assign _03192_ = \mchip.index [10] & ~_03191_;
	assign _03193_ = _01671_ | \mchip.index [8];
	assign _03194_ = \mchip.index [10] & ~_03193_;
	assign _03196_ = _01189_ | \mchip.index [7];
	assign _03197_ = _03196_ | \mchip.index [9];
	assign _03198_ = _03197_ | \mchip.index [10];
	assign _03199_ = _01875_ & ~_03198_;
	assign _03200_ = _00463_ | \mchip.index [5];
	assign _03201_ = _03200_ | _02984_;
	assign _03202_ = _03201_ | _02097_;
	assign _03203_ = _03202_ | _04648_;
	assign _03204_ = _03203_ | _07758_;
	assign _03205_ = _01986_ & ~_03204_;
	assign _03208_ = \mchip.index [11] & ~_02054_;
	assign _03209_ = _02542_ | _02097_;
	assign _03210_ = _03209_ | \mchip.index [10];
	assign _03211_ = \mchip.index [11] & ~_03210_;
	assign _03212_ = _02431_ | _02097_;
	assign _03213_ = _03212_ | \mchip.index [10];
	assign _03214_ = \mchip.index [11] & ~_03213_;
	assign _03215_ = _00561_ | \mchip.index [9];
	assign _03216_ = _03215_ | \mchip.index [10];
	assign _03217_ = _01875_ & ~_03216_;
	assign _03219_ = _02500_ | \mchip.index [7];
	assign _03220_ = _03219_ | _04648_;
	assign _03221_ = _03220_ | \mchip.index [10];
	assign _03222_ = \mchip.index [11] & ~_03221_;
	assign _03223_ = _00395_ | _02097_;
	assign _03224_ = _03223_ | \mchip.index [8];
	assign _03225_ = _03224_ | _07758_;
	assign _03226_ = \mchip.index [10] & ~_03225_;
	assign _03227_ = _00530_ | \mchip.index [7];
	assign _03228_ = _03227_ | \mchip.index [8];
	assign _03230_ = _03228_ | _07758_;
	assign _03231_ = \mchip.index [10] & ~_03230_;
	assign _03232_ = _01792_ | \mchip.index [9];
	assign _03233_ = _01986_ & ~_03232_;
	assign _03234_ = _00559_ | _02097_;
	assign _03235_ = _03234_ | _04648_;
	assign _03236_ = _03235_ | _07758_;
	assign _03237_ = _01986_ & ~_03236_;
	assign _03238_ = _01551_ | _02097_;
	assign _03239_ = _03238_ | _04648_;
	assign _03241_ = _03239_ | _01986_;
	assign _03242_ = _01875_ & ~_03241_;
	assign _03243_ = _01708_ | _02984_;
	assign _03244_ = _03243_ | \mchip.index [7];
	assign _03245_ = _03244_ | _07758_;
	assign _03246_ = _03245_ | _01986_;
	assign _03247_ = _01875_ & ~_03246_;
	assign _03248_ = _02801_ | \mchip.index [9];
	assign _03249_ = \mchip.index [11] & ~_03248_;
	assign _03250_ = ~(_05037_ & _01986_);
	assign _03252_ = _01875_ & ~_03250_;
	assign _03253_ = _01687_ | \mchip.index [6];
	assign _03254_ = _03253_ | \mchip.index [7];
	assign _03255_ = _03254_ | \mchip.index [9];
	assign _03256_ = _03255_ | \mchip.index [10];
	assign _03257_ = _01875_ & ~_03256_;
	assign _03258_ = _03002_ | _04648_;
	assign _03259_ = \mchip.index [11] & ~_03258_;
	assign _03260_ = _01152_ | \mchip.index [6];
	assign _03261_ = _03260_ | _02097_;
	assign _03263_ = _03261_ | _07758_;
	assign _03264_ = _03263_ | \mchip.index [10];
	assign _03265_ = \mchip.index [11] & ~_03264_;
	assign _03266_ = _01481_ | _04648_;
	assign _03267_ = _03266_ | _07758_;
	assign _03268_ = _01986_ & ~_03267_;
	assign _03269_ = _07828_ | _02984_;
	assign _03270_ = _03269_ | \mchip.index [8];
	assign _03271_ = _03270_ | \mchip.index [9];
	assign _03272_ = \mchip.index [10] & ~_03271_;
	assign _03274_ = _03916_ | \mchip.index [7];
	assign _03275_ = _03274_ | \mchip.index [8];
	assign _03276_ = _03275_ | \mchip.index [9];
	assign _03277_ = \mchip.index [10] & ~_03276_;
	assign _03278_ = _00110_ | _02984_;
	assign _03279_ = _03278_ | \mchip.index [7];
	assign _03280_ = _03279_ | _04648_;
	assign _03281_ = _03280_ | \mchip.index [10];
	assign _03282_ = \mchip.index [11] & ~_03281_;
	assign _03283_ = _07721_ | _02984_;
	assign _03285_ = _03283_ | \mchip.index [8];
	assign _03286_ = _03285_ | _07758_;
	assign _03287_ = _01986_ & ~_03286_;
	assign _03288_ = _01586_ | \mchip.index [8];
	assign _03289_ = _03288_ | \mchip.index [9];
	assign _03290_ = \mchip.index [10] & ~_03289_;
	assign _03291_ = _01353_ | \mchip.index [7];
	assign _03292_ = _03291_ | _04648_;
	assign _03293_ = _03292_ | \mchip.index [9];
	assign _03294_ = \mchip.index [10] & ~_03293_;
	assign _03296_ = _07455_ | _02097_;
	assign _03297_ = _03296_ | \mchip.index [8];
	assign _03298_ = \mchip.index [9] & ~_03297_;
	assign _03299_ = _07746_ | _04648_;
	assign _03300_ = _03299_ | \mchip.index [9];
	assign _03301_ = \mchip.index [10] & ~_03300_;
	assign _03302_ = _01716_ | \mchip.index [7];
	assign _03303_ = _03302_ | \mchip.index [8];
	assign _03304_ = \mchip.index [9] & ~_03303_;
	assign _03305_ = _03562_ | \mchip.index [10];
	assign _03307_ = _01875_ & ~_03305_;
	assign _03308_ = _01485_ | _02097_;
	assign _03309_ = _03308_ | _04648_;
	assign _03310_ = _03309_ | \mchip.index [10];
	assign _03311_ = _01875_ & ~_03310_;
	assign _03312_ = _01486_ | \mchip.index [8];
	assign _03313_ = \mchip.index [9] & ~_03312_;
	assign _03314_ = _01133_ | _02097_;
	assign _03315_ = _03314_ | _04648_;
	assign _03316_ = _03315_ | _07758_;
	assign _03319_ = _01875_ & ~_03316_;
	assign _03320_ = _07653_ | \mchip.index [6];
	assign _03321_ = _03320_ | \mchip.index [7];
	assign _03322_ = _03321_ | _04648_;
	assign _03323_ = _03322_ | _07758_;
	assign _03324_ = _01986_ & ~_03323_;
	assign _03325_ = _01153_ | _02097_;
	assign _03326_ = _03325_ | _04648_;
	assign _03327_ = _03326_ | _07758_;
	assign _03328_ = _01986_ & ~_03327_;
	assign _03330_ = _01542_ | \mchip.index [8];
	assign _03331_ = _03330_ | \mchip.index [9];
	assign _03332_ = \mchip.index [10] & ~_03331_;
	assign _03333_ = _01133_ | \mchip.index [8];
	assign _03334_ = _03333_ | _07758_;
	assign _03335_ = \mchip.index [10] & ~_03334_;
	assign _03336_ = _06378_ | _02984_;
	assign _03337_ = _03336_ | _02097_;
	assign _03338_ = _03337_ | _04648_;
	assign _03339_ = _03338_ | \mchip.index [9];
	assign _03341_ = \mchip.index [10] & ~_03339_;
	assign _03342_ = _07675_ | _05424_;
	assign _03343_ = _03342_ | _02097_;
	assign _03344_ = _03343_ | \mchip.index [9];
	assign _03345_ = _01986_ & ~_03344_;
	assign _03346_ = _02419_ | _02097_;
	assign _03347_ = _03346_ | \mchip.index [8];
	assign _03348_ = _03347_ | \mchip.index [9];
	assign _03349_ = \mchip.index [10] & ~_03348_;
	assign _03350_ = _01309_ | \mchip.index [8];
	assign _03352_ = _03350_ | _07758_;
	assign _03353_ = \mchip.index [10] & ~_03352_;
	assign _03354_ = _01384_ | \mchip.index [7];
	assign _03355_ = _03354_ | _04648_;
	assign _03356_ = _01986_ & ~_03355_;
	assign _03357_ = _00411_ | _02097_;
	assign _03358_ = _03357_ | _01986_;
	assign _03359_ = \mchip.index [11] & ~_03358_;
	assign _03360_ = _02707_ | \mchip.index [7];
	assign _03361_ = _03360_ | _04648_;
	assign _03363_ = _03361_ | \mchip.index [9];
	assign _03364_ = \mchip.index [11] & ~_03363_;
	assign _03365_ = _02602_ | \mchip.index [8];
	assign _03366_ = \mchip.index [11] & ~_03365_;
	assign _03367_ = _01629_ | _02097_;
	assign _03368_ = _03367_ | _04648_;
	assign _03369_ = _03368_ | \mchip.index [9];
	assign _03370_ = _01986_ & ~_03369_;
	assign _03371_ = _01189_ | \mchip.index [6];
	assign _03372_ = _03371_ | \mchip.index [7];
	assign _03374_ = _03372_ | \mchip.index [8];
	assign _03375_ = _07758_ & ~_03374_;
	assign _03376_ = _01259_ | _07758_;
	assign _03377_ = \mchip.index [10] & ~_03376_;
	assign _03378_ = _04893_ | _02097_;
	assign _03379_ = _04648_ & ~_03378_;
	assign _03380_ = _07768_ | \mchip.index [6];
	assign _03381_ = _03380_ | \mchip.index [7];
	assign _03382_ = _03381_ | _07758_;
	assign _03383_ = _03382_ | \mchip.index [10];
	assign _03385_ = \mchip.index [11] & ~_03383_;
	assign _03386_ = _02134_ | _04648_;
	assign _03387_ = _03386_ | _07758_;
	assign _03388_ = _01986_ & ~_03387_;
	assign _03389_ = _07828_ | _05424_;
	assign _03390_ = _03389_ | \mchip.index [6];
	assign _03391_ = _03390_ | _02097_;
	assign _03392_ = \mchip.index [11] & ~_03391_;
	assign _03393_ = _00879_ | _02984_;
	assign _03394_ = _03393_ | \mchip.index [7];
	assign _03396_ = _03394_ | \mchip.index [8];
	assign _03397_ = _03396_ | \mchip.index [9];
	assign _03398_ = \mchip.index [10] & ~_03397_;
	assign _03399_ = _01305_ | \mchip.index [7];
	assign _03400_ = _03399_ | _04648_;
	assign _03401_ = \mchip.index [11] & ~_03400_;
	assign _03402_ = _01943_ | _07758_;
	assign _03403_ = _03402_ | \mchip.index [10];
	assign _03404_ = \mchip.index [11] & ~_03403_;
	assign _03405_ = _01168_ | _07758_;
	assign _03407_ = \mchip.index [11] & ~_03405_;
	assign _03408_ = _01849_ | \mchip.index [6];
	assign _03409_ = _03408_ | _02097_;
	assign _03410_ = _03409_ | \mchip.index [8];
	assign _03411_ = _03410_ | \mchip.index [9];
	assign _03412_ = \mchip.index [10] & ~_03411_;
	assign _03413_ = _07768_ | _02984_;
	assign _03414_ = _03413_ | \mchip.index [7];
	assign _03415_ = _03414_ | \mchip.index [8];
	assign _03416_ = _03415_ | \mchip.index [9];
	assign _03418_ = \mchip.index [11] & ~_03416_;
	assign _03419_ = _07843_ | \mchip.index [6];
	assign _03420_ = _03419_ | \mchip.index [7];
	assign _03421_ = _03420_ | _01986_;
	assign _03422_ = \mchip.index [11] & ~_03421_;
	assign _03423_ = ~(_00338_ & _07758_);
	assign _03424_ = _03423_ | \mchip.index [10];
	assign _03425_ = _01875_ & ~_03424_;
	assign _03426_ = _02057_ | _02097_;
	assign _03427_ = _03426_ | \mchip.index [9];
	assign _03430_ = _03427_ | \mchip.index [10];
	assign _03431_ = \mchip.index [11] & ~_03430_;
	assign _03432_ = _02157_ | \mchip.index [7];
	assign _03433_ = _03432_ | _04648_;
	assign _03434_ = \mchip.index [11] & ~_03433_;
	assign _03435_ = _01528_ | \mchip.index [7];
	assign _03436_ = _03435_ | _04648_;
	assign _03437_ = _03436_ | _01986_;
	assign _03438_ = _01875_ & ~_03437_;
	assign _03439_ = _01874_ | \mchip.index [7];
	assign _03441_ = _03439_ | _04648_;
	assign _03442_ = _03441_ | _07758_;
	assign _03443_ = _01986_ & ~_03442_;
	assign _03444_ = _01245_ | \mchip.index [7];
	assign _03445_ = _03444_ | _04648_;
	assign _03446_ = _03445_ | _07758_;
	assign _03447_ = _03446_ | _01986_;
	assign _03448_ = _01875_ & ~_03447_;
	assign _03449_ = _01943_ | _02984_;
	assign _03450_ = _03449_ | \mchip.index [8];
	assign _03452_ = _03450_ | _07758_;
	assign _03453_ = \mchip.index [10] & ~_03452_;
	assign _03454_ = _07720_ | _05424_;
	assign _03455_ = _03454_ | _02097_;
	assign _03456_ = _03455_ | \mchip.index [8];
	assign _03457_ = \mchip.index [9] & ~_03456_;
	assign _03458_ = _03095_ | _02097_;
	assign _03459_ = _03458_ | \mchip.index [8];
	assign _03460_ = _03459_ | _07758_;
	assign _03461_ = \mchip.index [11] & ~_03460_;
	assign _03463_ = _00571_ | _02984_;
	assign _03464_ = _03463_ | \mchip.index [7];
	assign _03465_ = _03464_ | _04648_;
	assign _03466_ = _03465_ | \mchip.index [9];
	assign _03467_ = \mchip.index [10] & ~_03466_;
	assign _03468_ = _01840_ | \mchip.index [8];
	assign _03469_ = _03468_ | \mchip.index [9];
	assign _03470_ = \mchip.index [11] & ~_03469_;
	assign _03471_ = _02015_ | _02097_;
	assign _03472_ = _03471_ | _04648_;
	assign _03474_ = _03472_ | \mchip.index [9];
	assign _03475_ = \mchip.index [11] & ~_03474_;
	assign _03476_ = _03235_ | \mchip.index [9];
	assign _03477_ = \mchip.index [10] & ~_03476_;
	assign _03478_ = _01278_ | \mchip.index [8];
	assign _03479_ = _03478_ | _07758_;
	assign _03480_ = \mchip.index [10] & ~_03479_;
	assign _03481_ = _00527_ | \mchip.index [7];
	assign _03482_ = _03481_ | \mchip.index [8];
	assign _03483_ = \mchip.index [11] & ~_03482_;
	assign _03485_ = _06545_ | \mchip.index [5];
	assign _03486_ = _03485_ | _02984_;
	assign _03487_ = _03486_ | \mchip.index [7];
	assign _03488_ = _03487_ | _01986_;
	assign _03489_ = \mchip.index [11] & ~_03488_;
	assign _03490_ = _03489_ | _03483_;
	assign _03491_ = _03490_ | _03480_;
	assign _03492_ = _03491_ | _03477_;
	assign _03493_ = _03492_ | _03475_;
	assign _03494_ = _03493_ | _03470_;
	assign _03496_ = _03494_ | _03467_;
	assign _03497_ = _03496_ | _03461_;
	assign _03498_ = _03497_ | _03457_;
	assign _03499_ = _03498_ | _03453_;
	assign _03500_ = _03499_ | _03448_;
	assign _03501_ = _03500_ | _03443_;
	assign _03502_ = _03501_ | _03438_;
	assign _03503_ = _03502_ | _03434_;
	assign _03504_ = _03503_ | _03431_;
	assign _03505_ = _03504_ | _03425_;
	assign _03507_ = _03505_ | _03422_;
	assign _03508_ = _03507_ | _03418_;
	assign _03509_ = _03508_ | _03412_;
	assign _03510_ = _03509_ | _03407_;
	assign _03511_ = _03510_ | _03404_;
	assign _03512_ = _03511_ | _03401_;
	assign _03513_ = _03512_ | _03398_;
	assign _03514_ = _03513_ | _03392_;
	assign _03515_ = _03514_ | _03388_;
	assign _03516_ = _03515_ | _03385_;
	assign _03518_ = _03516_ | _03379_;
	assign _03519_ = _03518_ | _03377_;
	assign _03520_ = _03519_ | _03375_;
	assign _03521_ = _03520_ | _03370_;
	assign _03522_ = _03521_ | _03366_;
	assign _03523_ = _03522_ | _03364_;
	assign _03524_ = _03523_ | _03359_;
	assign _03525_ = _03524_ | _03356_;
	assign _03526_ = _03525_ | _03353_;
	assign _03527_ = _03526_ | _03349_;
	assign _03529_ = _03527_ | _03345_;
	assign _03530_ = _03529_ | _03341_;
	assign _03531_ = _03530_ | _03335_;
	assign _03532_ = _03531_ | _03332_;
	assign _03533_ = _03532_ | _03328_;
	assign _03534_ = _03533_ | _03324_;
	assign _03535_ = _03534_ | _03319_;
	assign _03536_ = _03535_ | _03313_;
	assign _03537_ = _03536_ | _03311_;
	assign _03538_ = _03537_ | _03307_;
	assign _03541_ = _03538_ | _03304_;
	assign _03542_ = _03541_ | _03301_;
	assign _03543_ = _03542_ | _03298_;
	assign _03544_ = _03543_ | _03294_;
	assign _03545_ = _03544_ | _03290_;
	assign _03546_ = _03545_ | _03287_;
	assign _03547_ = _03546_ | _03282_;
	assign _03548_ = _03547_ | _03277_;
	assign _03549_ = _03548_ | _03272_;
	assign _03550_ = _03549_ | _03268_;
	assign _03552_ = _03550_ | _03265_;
	assign _03553_ = _03552_ | _03259_;
	assign _03554_ = _03553_ | _03257_;
	assign _03555_ = _03554_ | _03252_;
	assign _03556_ = _03555_ | _03249_;
	assign _03557_ = _03556_ | _03247_;
	assign _03558_ = _03557_ | _03242_;
	assign _03559_ = _03558_ | _03237_;
	assign _03560_ = _03559_ | _03233_;
	assign _03561_ = _03560_ | _03231_;
	assign _03563_ = _03561_ | _03226_;
	assign _03564_ = _03563_ | _03222_;
	assign _03565_ = _03564_ | _03217_;
	assign _03566_ = _03565_ | _03214_;
	assign _03567_ = _03566_ | _03211_;
	assign _03568_ = _03567_ | _03208_;
	assign _03569_ = _03568_ | _03205_;
	assign _03570_ = _03569_ | _03199_;
	assign _03571_ = _03570_ | _03194_;
	assign _03572_ = _03571_ | _03192_;
	assign _03574_ = _03572_ | _03189_;
	assign _03575_ = _03574_ | _03183_;
	assign _03576_ = _03575_ | _03180_;
	assign _03577_ = _03576_ | _03175_;
	assign _03578_ = _03577_ | _03171_;
	assign _03579_ = _03578_ | _03168_;
	assign _03580_ = _03579_ | _03164_;
	assign _03581_ = _03580_ | _03158_;
	assign _03582_ = _03581_ | _03153_;
	assign _03583_ = _03582_ | _03150_;
	assign _03585_ = _03583_ | _03147_;
	assign _03586_ = _03585_ | _03142_;
	assign _03587_ = _03586_ | _03137_;
	assign _03588_ = _03587_ | _03132_;
	assign _03589_ = _03588_ | _03126_;
	assign _03590_ = _03589_ | _03123_;
	assign _03591_ = _03590_ | _03120_;
	assign _03592_ = _03591_ | _03114_;
	assign _03593_ = _03592_ | _03109_;
	assign _03594_ = _03593_ | _03105_;
	assign _03596_ = _03594_ | _03102_;
	assign _03597_ = _03596_ | _03099_;
	assign _03598_ = _03597_ | _03094_;
	assign _03599_ = _03598_ | _03090_;
	assign _03600_ = _03599_ | _03087_;
	assign _03601_ = _03600_ | _03082_;
	assign _03602_ = _03601_ | _03079_;
	assign _03603_ = _03602_ | _03072_;
	assign _03604_ = _03603_ | _03068_;
	assign _03605_ = _03604_ | _03065_;
	assign _03607_ = _03605_ | _03061_;
	assign _03608_ = _03607_ | _03056_;
	assign _03609_ = _03608_ | _03054_;
	assign _03610_ = _03609_ | _03050_;
	assign _03611_ = _03610_ | _03046_;
	assign _03612_ = _03611_ | _03045_;
	assign _03613_ = _03612_ | _03042_;
	assign _03614_ = _03613_ | _03038_;
	assign _03615_ = _03614_ | _03034_;
	assign _03616_ = _03615_ | _03032_;
	assign _03618_ = _03616_ | _03027_;
	assign _03619_ = _03618_ | _03024_;
	assign _03620_ = _03619_ | _03022_;
	assign _03621_ = _03620_ | _03015_;
	assign _03622_ = _03621_ | _03012_;
	assign _03623_ = _03622_ | _03009_;
	assign _03624_ = _03623_ | _03004_;
	assign _03625_ = _03624_ | _03001_;
	assign _03626_ = _03625_ | _02994_;
	assign _03627_ = _03626_ | _02988_;
	assign _03629_ = _03627_ | _02983_;
	assign _03630_ = _03629_ | _02979_;
	assign _03631_ = _03630_ | _02974_;
	assign _03632_ = _03631_ | _02969_;
	assign _03633_ = _03632_ | _02965_;
	assign _03634_ = _03633_ | _02959_;
	assign _03635_ = _03634_ | _02955_;
	assign _03636_ = _03635_ | _02950_;
	assign _03637_ = _03636_ | _02946_;
	assign _03638_ = _03637_ | _02941_;
	assign _03640_ = _03638_ | _02937_;
	assign _03641_ = _03640_ | _02935_;
	assign _03642_ = _03641_ | _02930_;
	assign _03643_ = _03642_ | _02924_;
	assign _03644_ = _03643_ | _02920_;
	assign _03645_ = _03644_ | _02915_;
	assign _03646_ = _03645_ | _02910_;
	assign _03647_ = _03646_ | _02905_;
	assign _03648_ = _03647_ | _02903_;
	assign _03649_ = _03648_ | _02900_;
	assign _03652_ = _03649_ | _02894_;
	assign _03653_ = _03652_ | _02889_;
	assign _03654_ = _03653_ | _02883_;
	assign _03655_ = _03654_ | _02879_;
	assign _03656_ = _03655_ | _02872_;
	assign _03657_ = _03656_ | _02868_;
	assign _03658_ = _03657_ | _02865_;
	assign _03659_ = _03658_ | _02864_;
	assign _03660_ = _03659_ | _02860_;
	assign _03661_ = _03660_ | _02854_;
	assign _03663_ = _03661_ | _02849_;
	assign _03664_ = _03663_ | _02845_;
	assign _03665_ = _03664_ | _02839_;
	assign _03666_ = _03665_ | _02835_;
	assign _03667_ = _03666_ | _02833_;
	assign _03668_ = _03667_ | _02827_;
	assign _03669_ = _03668_ | _02822_;
	assign _03670_ = _03669_ | _02817_;
	assign _03671_ = _03670_ | _02815_;
	assign _03672_ = _03671_ | _02813_;
	assign _03674_ = _03672_ | _02809_;
	assign _03675_ = _03674_ | _02804_;
	assign _03676_ = _03675_ | _02799_;
	assign _03677_ = _03676_ | _02794_;
	assign _03678_ = _03677_ | _02789_;
	assign _03679_ = _03678_ | _02784_;
	assign _03680_ = _03679_ | _02781_;
	assign _03681_ = _03680_ | _02779_;
	assign _03682_ = _03681_ | _02773_;
	assign _03683_ = _03682_ | _02769_;
	assign _03685_ = _03683_ | _02766_;
	assign _03686_ = _03685_ | _02761_;
	assign _03687_ = _03686_ | _02757_;
	assign _03688_ = _03687_ | _02754_;
	assign _03689_ = _03688_ | _02749_;
	assign _03690_ = _03689_ | _02747_;
	assign _03691_ = _03690_ | _02742_;
	assign _03692_ = _03691_ | _02739_;
	assign _03693_ = _03692_ | _02736_;
	assign _03694_ = _03693_ | _02732_;
	assign _03696_ = _03694_ | _02727_;
	assign _03697_ = _03696_ | _02723_;
	assign _03698_ = _03697_ | _02717_;
	assign _03699_ = _03698_ | _02712_;
	assign _03700_ = _03699_ | _02708_;
	assign _03701_ = _03700_ | _02703_;
	assign _03702_ = _03701_ | _02698_;
	assign _03703_ = _03702_ | _02693_;
	assign _03704_ = _03703_ | _02690_;
	assign _03705_ = _03704_ | _02687_;
	assign _03707_ = _03705_ | _02683_;
	assign _03708_ = _03707_ | _02680_;
	assign _03709_ = _03708_ | _02676_;
	assign _03710_ = _03709_ | _02671_;
	assign _03711_ = _03710_ | _02667_;
	assign _03712_ = _03711_ | _02660_;
	assign _03713_ = _03712_ | _02657_;
	assign _03714_ = _03713_ | _02654_;
	assign _03715_ = _03714_ | _02648_;
	assign _03716_ = _03715_ | _02645_;
	assign _03718_ = _03716_ | _02644_;
	assign _03719_ = _03718_ | _02642_;
	assign _03720_ = _03719_ | _02638_;
	assign _03721_ = _03720_ | _02634_;
	assign _03722_ = _03721_ | _02630_;
	assign _03723_ = _03722_ | _02624_;
	assign _03724_ = _03723_ | _02623_;
	assign _03725_ = _03724_ | _02619_;
	assign _03726_ = _03725_ | _02615_;
	assign _03727_ = _03726_ | _02611_;
	assign _03729_ = _03727_ | _02605_;
	assign _03730_ = _03729_ | _02599_;
	assign _03731_ = _03730_ | _02592_;
	assign _03732_ = _03731_ | _02588_;
	assign _03733_ = _03732_ | _02586_;
	assign _03734_ = _03733_ | _02579_;
	assign _03735_ = _03734_ | _02572_;
	assign _03736_ = _03735_ | _02568_;
	assign _03737_ = _03736_ | _02564_;
	assign _03738_ = _03737_ | _02560_;
	assign _03740_ = _03738_ | _02558_;
	assign _03741_ = _03740_ | _02551_;
	assign _03742_ = _03741_ | _02548_;
	assign _03743_ = _03742_ | _02546_;
	assign _03744_ = _03743_ | _02539_;
	assign _03745_ = _03744_ | _02536_;
	assign _03746_ = _03745_ | _02534_;
	assign _03747_ = _03746_ | _02530_;
	assign _03748_ = _03747_ | _02524_;
	assign _03749_ = _03748_ | _02522_;
	assign _03751_ = _03749_ | _02517_;
	assign _03752_ = _03751_ | _02515_;
	assign _03753_ = _03752_ | _02509_;
	assign _03754_ = _03753_ | _02504_;
	assign _03755_ = _03754_ | _02499_;
	assign _03756_ = _03755_ | _02494_;
	assign _03757_ = _03756_ | _02491_;
	assign _03758_ = _03757_ | _02490_;
	assign _03759_ = _03758_ | _02484_;
	assign _03760_ = _03759_ | _02480_;
	assign _03763_ = _03760_ | _02476_;
	assign _03764_ = _03763_ | _02471_;
	assign _03765_ = _03764_ | _02468_;
	assign _03766_ = _03765_ | _02466_;
	assign _03767_ = _03766_ | _02460_;
	assign _03768_ = _03767_ | _02457_;
	assign _03769_ = _03768_ | _02454_;
	assign _03770_ = _03769_ | _02451_;
	assign _03771_ = _03770_ | _02448_;
	assign \mchip.val [3] = _03771_ | _02443_;
	assign _03773_ = _00822_ | \mchip.index [6];
	assign _03774_ = _03773_ | \mchip.index [7];
	assign _03775_ = _03774_ | \mchip.index [8];
	assign _03776_ = \mchip.index [11] & ~_03775_;
	assign _03777_ = _01354_ | \mchip.index [9];
	assign _03778_ = _03777_ | \mchip.index [10];
	assign _03779_ = _01875_ & ~_03778_;
	assign _03780_ = _01379_ | _02097_;
	assign _03781_ = _03780_ | _04648_;
	assign _03782_ = _07758_ & ~_03781_;
	assign _03784_ = _07725_ | _02984_;
	assign _03785_ = _03784_ | \mchip.index [7];
	assign _03786_ = _03785_ | _07758_;
	assign _03787_ = \mchip.index [11] & ~_03786_;
	assign _03788_ = _07792_ | _02097_;
	assign _03789_ = _03788_ | \mchip.index [8];
	assign _03790_ = _03789_ | \mchip.index [9];
	assign _03791_ = \mchip.index [11] & ~_03790_;
	assign _03792_ = _02681_ | _07758_;
	assign _03793_ = _01875_ & ~_03792_;
	assign _03795_ = _01806_ | _04648_;
	assign _03796_ = _03795_ | _07758_;
	assign _03797_ = _01986_ & ~_03796_;
	assign _03798_ = _05447_ | \mchip.index [9];
	assign _03799_ = \mchip.index [10] & ~_03798_;
	assign _03800_ = _06600_ | _04648_;
	assign _03801_ = _07758_ & ~_03800_;
	assign _03802_ = _00607_ | _02097_;
	assign _03803_ = _03802_ | \mchip.index [9];
	assign _03804_ = \mchip.index [10] & ~_03803_;
	assign _03806_ = _07804_ | \mchip.index [6];
	assign _03807_ = _03806_ | _02097_;
	assign _03808_ = _03807_ | \mchip.index [8];
	assign _03809_ = _03808_ | \mchip.index [9];
	assign _03810_ = _01986_ & ~_03809_;
	assign _03811_ = _02580_ | \mchip.index [7];
	assign _03812_ = _03811_ | \mchip.index [8];
	assign _03813_ = _03812_ | _01986_;
	assign _03814_ = _01875_ & ~_03813_;
	assign _03815_ = _01326_ | _02097_;
	assign _03817_ = _03815_ | \mchip.index [8];
	assign _03818_ = _03817_ | \mchip.index [9];
	assign _03819_ = _03818_ | \mchip.index [10];
	assign _03820_ = \mchip.index [11] & ~_03819_;
	assign _03821_ = _02840_ | \mchip.index [7];
	assign _03822_ = _03821_ | _04648_;
	assign _03823_ = _03822_ | \mchip.index [9];
	assign _03824_ = \mchip.index [10] & ~_03823_;
	assign _03825_ = _02961_ | _02097_;
	assign _03826_ = _03825_ | _04648_;
	assign _03828_ = _03826_ | _07758_;
	assign _03829_ = _03828_ | _01986_;
	assign _03830_ = _01875_ & ~_03829_;
	assign _03831_ = _02730_ | _04648_;
	assign _03832_ = \mchip.index [9] & ~_03831_;
	assign _03833_ = _03219_ | \mchip.index [8];
	assign _03834_ = \mchip.index [9] & ~_03833_;
	assign _03835_ = _01147_ | _04648_;
	assign _03836_ = _03835_ | \mchip.index [9];
	assign _03837_ = \mchip.index [10] & ~_03836_;
	assign _03839_ = _01944_ | \mchip.index [8];
	assign _03840_ = _03839_ | _07758_;
	assign _03841_ = \mchip.index [10] & ~_03840_;
	assign _03842_ = _01104_ | \mchip.index [7];
	assign _03843_ = _03842_ | \mchip.index [8];
	assign _03844_ = \mchip.index [9] & ~_03843_;
	assign _03845_ = _01104_ | _01986_;
	assign _03846_ = \mchip.index [11] & ~_03845_;
	assign _03847_ = _01501_ | \mchip.index [6];
	assign _03848_ = _03847_ | \mchip.index [9];
	assign _03850_ = _03848_ | \mchip.index [10];
	assign _03851_ = _01875_ & ~_03850_;
	assign _03852_ = _00255_ | _05424_;
	assign _03853_ = _02984_ & ~_03852_;
	assign _03854_ = _03706_ | _04648_;
	assign _03855_ = _03854_ | \mchip.index [10];
	assign _03856_ = \mchip.index [11] & ~_03855_;
	assign _03857_ = _00484_ | \mchip.index [6];
	assign _03858_ = _03857_ | \mchip.index [7];
	assign _03859_ = _03858_ | \mchip.index [9];
	assign _03861_ = _03859_ | \mchip.index [10];
	assign _03862_ = _01875_ & ~_03861_;
	assign _03863_ = _04993_ | \mchip.index [5];
	assign _03864_ = _03863_ | _02984_;
	assign _03865_ = _03864_ | \mchip.index [7];
	assign _03866_ = _03865_ | \mchip.index [8];
	assign _03867_ = _03866_ | _07758_;
	assign _03868_ = \mchip.index [10] & ~_03867_;
	assign _03869_ = _05180_ | _01098_;
	assign _03870_ = _03869_ | _02984_;
	assign _03873_ = _03870_ | _02097_;
	assign _03874_ = _03873_ | _04648_;
	assign _03875_ = _03874_ | \mchip.index [10];
	assign _03876_ = \mchip.index [11] & ~_03875_;
	assign _03877_ = _05979_ | _05424_;
	assign _03878_ = _03877_ | \mchip.index [8];
	assign _03879_ = _03878_ | \mchip.index [10];
	assign _03880_ = _01875_ & ~_03879_;
	assign _03881_ = _00687_ | \mchip.index [7];
	assign _03882_ = _03881_ | \mchip.index [8];
	assign _03884_ = \mchip.index [9] & ~_03882_;
	assign _03885_ = _03927_ | _02097_;
	assign _03886_ = _03885_ | \mchip.index [8];
	assign _03887_ = \mchip.index [9] & ~_03886_;
	assign _03888_ = _02625_ | _02984_;
	assign _03889_ = _03888_ | \mchip.index [8];
	assign _03890_ = _03889_ | _07758_;
	assign _03891_ = \mchip.index [10] & ~_03890_;
	assign _03892_ = \mchip.index [10] & ~_01683_;
	assign _03893_ = _01494_ | _04648_;
	assign _03895_ = _03893_ | _07758_;
	assign _03896_ = _01986_ & ~_03895_;
	assign _03897_ = _01202_ | \mchip.index [8];
	assign _03898_ = _03897_ | _07758_;
	assign _03899_ = _03898_ | \mchip.index [10];
	assign _03900_ = _01875_ & ~_03899_;
	assign _03901_ = _01197_ | \mchip.index [8];
	assign _03902_ = _03901_ | _07758_;
	assign _03903_ = _03902_ | \mchip.index [10];
	assign _03904_ = _01875_ & ~_03903_;
	assign _03906_ = _00835_ | \mchip.index [5];
	assign _03907_ = _03906_ | \mchip.index [6];
	assign _03908_ = _03907_ | _02097_;
	assign _03909_ = _03908_ | _07758_;
	assign _03910_ = \mchip.index [11] & ~_03909_;
	assign _03911_ = _03378_ | _07758_;
	assign _03912_ = _03911_ | _01986_;
	assign _03913_ = _01875_ & ~_03912_;
	assign _03914_ = _01179_ | \mchip.index [9];
	assign _03915_ = _03914_ | \mchip.index [10];
	assign _03917_ = _01875_ & ~_03915_;
	assign _03918_ = _01629_ | \mchip.index [9];
	assign _03919_ = \mchip.index [11] & ~_03918_;
	assign _03920_ = _02851_ | _02097_;
	assign _03921_ = \mchip.index [11] & ~_03920_;
	assign _03922_ = _02461_ | _02097_;
	assign _03923_ = _03922_ | _04648_;
	assign _03924_ = _03923_ | \mchip.index [10];
	assign _03925_ = _01875_ & ~_03924_;
	assign _03926_ = _01943_ | _02097_;
	assign _03928_ = \mchip.index [11] & ~_03926_;
	assign _03929_ = _00531_ | _02097_;
	assign _03930_ = _03929_ | _07758_;
	assign _03931_ = \mchip.index [11] & ~_03930_;
	assign _03932_ = _01848_ | _02984_;
	assign _03933_ = _03932_ | \mchip.index [8];
	assign _03934_ = _03933_ | \mchip.index [9];
	assign _03935_ = _03934_ | \mchip.index [10];
	assign _03936_ = _01875_ & ~_03935_;
	assign _03937_ = _01492_ | \mchip.index [6];
	assign _03939_ = _03937_ | _02097_;
	assign _03940_ = _03939_ | _04648_;
	assign _03941_ = _03940_ | \mchip.index [9];
	assign _03942_ = _01875_ & ~_03941_;
	assign _03943_ = _00835_ | _02984_;
	assign _03944_ = _03943_ | \mchip.index [7];
	assign _03945_ = _03944_ | _04648_;
	assign _03946_ = _03945_ | _07758_;
	assign _03947_ = _03946_ | _01986_;
	assign _03948_ = _01875_ & ~_03947_;
	assign _03950_ = _03408_ | \mchip.index [7];
	assign _03951_ = _03950_ | \mchip.index [8];
	assign _03952_ = _03951_ | _07758_;
	assign _03953_ = \mchip.index [11] & ~_03952_;
	assign _03954_ = _01376_ | _05424_;
	assign _03955_ = _03954_ | _02097_;
	assign _03956_ = _03955_ | \mchip.index [8];
	assign _03957_ = \mchip.index [10] & ~_03956_;
	assign _03958_ = _03885_ | _04648_;
	assign _03959_ = \mchip.index [11] & ~_03958_;
	assign _03961_ = _03932_ | _02097_;
	assign _03962_ = _03961_ | \mchip.index [8];
	assign _03963_ = _03962_ | _07758_;
	assign _03964_ = \mchip.index [10] & ~_03963_;
	assign _03965_ = _00494_ & ~_01875_;
	assign _03966_ = _02661_ | _02984_;
	assign _03967_ = _03966_ | \mchip.index [8];
	assign _03968_ = _03967_ | _07758_;
	assign _03969_ = _01875_ & ~_03968_;
	assign _03970_ = _02685_ | _02984_;
	assign _03972_ = _03970_ | _02097_;
	assign _03973_ = _03972_ | _04648_;
	assign _03974_ = _03973_ | \mchip.index [9];
	assign _03975_ = _03974_ | \mchip.index [10];
	assign _03976_ = _01875_ & ~_03975_;
	assign _03977_ = _00811_ | \mchip.index [6];
	assign _03978_ = _03977_ | _02097_;
	assign _03979_ = _03978_ | _04648_;
	assign _03980_ = _03979_ | _07758_;
	assign _03981_ = _01986_ & ~_03980_;
	assign _03984_ = _01561_ | \mchip.index [6];
	assign _03985_ = _03984_ | \mchip.index [7];
	assign _03986_ = _03985_ | _01986_;
	assign _03987_ = \mchip.index [11] & ~_03986_;
	assign _03988_ = _02947_ | _02097_;
	assign _03989_ = _03988_ | _07758_;
	assign _03990_ = \mchip.index [10] & ~_03989_;
	assign _03991_ = _03095_ | \mchip.index [6];
	assign _03992_ = _03991_ | _02097_;
	assign _03993_ = _03992_ | _07758_;
	assign _03995_ = _01986_ & ~_03993_;
	assign _03996_ = _03033_ | \mchip.index [8];
	assign _03997_ = \mchip.index [10] & ~_03996_;
	assign _03998_ = _00684_ | \mchip.index [7];
	assign _03999_ = _03998_ | \mchip.index [8];
	assign _04000_ = \mchip.index [9] & ~_03999_;
	assign _04001_ = _00662_ | \mchip.index [6];
	assign _04002_ = _04001_ | _02097_;
	assign _04003_ = _04002_ | \mchip.index [10];
	assign _04004_ = _01875_ & ~_04003_;
	assign _04006_ = _02319_ | _05424_;
	assign _04007_ = _04006_ | \mchip.index [7];
	assign _04008_ = _04007_ | _04648_;
	assign _04009_ = _04008_ | \mchip.index [9];
	assign _04010_ = \mchip.index [10] & ~_04009_;
	assign _04011_ = _00022_ | \mchip.index [7];
	assign _04012_ = _04011_ | _01986_;
	assign _04013_ = \mchip.index [11] & ~_04012_;
	assign _04014_ = _02002_ | \mchip.index [8];
	assign _04015_ = \mchip.index [9] & ~_04014_;
	assign _04017_ = _00759_ | _02097_;
	assign _04018_ = _04017_ | _04648_;
	assign _04019_ = _04018_ | \mchip.index [10];
	assign _04020_ = _01875_ & ~_04019_;
	assign _04021_ = \mchip.index [8] & ~_02138_;
	assign _04022_ = _04871_ | \mchip.index [7];
	assign _04023_ = _04022_ | \mchip.index [8];
	assign _04024_ = _04023_ | \mchip.index [10];
	assign _04025_ = _01875_ & ~_04024_;
	assign _04026_ = _03811_ | \mchip.index [9];
	assign _04028_ = _04026_ | \mchip.index [10];
	assign _04029_ = \mchip.index [11] & ~_04028_;
	assign _04030_ = _01875_ & ~_01757_;
	assign _04031_ = _01379_ | _02984_;
	assign _04032_ = _04031_ | \mchip.index [9];
	assign _04033_ = \mchip.index [11] & ~_04032_;
	assign _04034_ = _02996_ | _02097_;
	assign _04035_ = _04034_ | _04648_;
	assign _04036_ = _04035_ | _07758_;
	assign _04037_ = _01875_ & ~_04036_;
	assign _04039_ = _01842_ | _02984_;
	assign _04040_ = _04039_ | \mchip.index [7];
	assign _04041_ = _04040_ | \mchip.index [8];
	assign _04042_ = _04041_ | _07758_;
	assign _04043_ = \mchip.index [10] & ~_04042_;
	assign _04044_ = _02397_ & ~_01875_;
	assign _04045_ = _01875_ & ~_03181_;
	assign _04046_ = _00337_ | _02097_;
	assign _04047_ = _04046_ | _04648_;
	assign _04048_ = _04047_ | _07758_;
	assign _04050_ = _01986_ & ~_04048_;
	assign _04051_ = _01875_ & ~_01505_;
	assign _04052_ = _01476_ | _02984_;
	assign _04053_ = _04052_ | \mchip.index [7];
	assign _04054_ = \mchip.index [10] & ~_04053_;
	assign _04055_ = _01731_ | \mchip.index [6];
	assign _04056_ = _04055_ | _02097_;
	assign _04057_ = _04056_ | _04648_;
	assign _04058_ = _04057_ | \mchip.index [9];
	assign _04059_ = _01875_ & ~_04058_;
	assign _04061_ = _03261_ | \mchip.index [9];
	assign _04062_ = _04061_ | \mchip.index [10];
	assign _04063_ = _01875_ & ~_04062_;
	assign _04064_ = _02176_ | \mchip.index [7];
	assign _04065_ = _04064_ | _07758_;
	assign _04066_ = _01875_ & ~_04065_;
	assign _04067_ = _03209_ | _04648_;
	assign _04068_ = _04067_ | _07758_;
	assign _04069_ = _01986_ & ~_04068_;
	assign _04070_ = _05004_ | _05424_;
	assign _04072_ = _04070_ | \mchip.index [9];
	assign _04073_ = \mchip.index [11] & ~_04072_;
	assign _04074_ = _03240_ | \mchip.index [8];
	assign _04075_ = _04074_ | \mchip.index [9];
	assign _04076_ = _01986_ & ~_04075_;
	assign _04077_ = _04076_ & ~\mchip.index [11];
	assign _04078_ = _02182_ | \mchip.index [9];
	assign _04079_ = \mchip.index [10] & ~_04078_;
	assign _04080_ = _01875_ & ~_02843_;
	assign _04081_ = _03916_ | \mchip.index [6];
	assign _04083_ = _04081_ | _04648_;
	assign _04084_ = _04083_ | _07758_;
	assign _04085_ = _01875_ & ~_04084_;
	assign _04086_ = _02601_ | \mchip.index [8];
	assign _04087_ = _04086_ | \mchip.index [9];
	assign _04088_ = \mchip.index [11] & ~_04087_;
	assign _04089_ = _07588_ | _05424_;
	assign _04090_ = _04089_ | _04648_;
	assign _04091_ = _01875_ & ~_04090_;
	assign _04092_ = _04006_ | \mchip.index [6];
	assign _04095_ = _04092_ | \mchip.index [8];
	assign _04096_ = _04095_ | _07758_;
	assign _04097_ = \mchip.index [10] & ~_04096_;
	assign _04098_ = _00759_ | _04648_;
	assign _04099_ = _04098_ | _07758_;
	assign _04100_ = _01986_ & ~_04099_;
	assign _04101_ = _02320_ | _05424_;
	assign _04102_ = _04101_ | _02984_;
	assign _04103_ = \mchip.index [8] & ~_04102_;
	assign _04104_ = _02565_ | _02097_;
	assign _04106_ = \mchip.index [9] & ~_04104_;
	assign _04107_ = _01569_ | \mchip.index [7];
	assign _04108_ = _04107_ | _07758_;
	assign _04109_ = _01875_ & ~_04108_;
	assign _04110_ = _04052_ | _04648_;
	assign _04111_ = _04110_ | _07758_;
	assign _04112_ = \mchip.index [10] & ~_04111_;
	assign _04113_ = _04304_ | _02984_;
	assign _04114_ = _04113_ | \mchip.index [7];
	assign _04115_ = _04114_ | _07758_;
	assign _04117_ = \mchip.index [11] & ~_04115_;
	assign _04118_ = _04460_ | _04648_;
	assign _04119_ = _04118_ | _07758_;
	assign _04120_ = \mchip.index [10] & ~_04119_;
	assign _04121_ = _00506_ | \mchip.index [6];
	assign _04122_ = _04121_ | _02097_;
	assign _04123_ = _04122_ | \mchip.index [8];
	assign _04124_ = _04123_ | \mchip.index [9];
	assign _04125_ = \mchip.index [11] & ~_04124_;
	assign _04126_ = _01979_ | \mchip.index [9];
	assign _04128_ = _01875_ & ~_04126_;
	assign _04129_ = _00692_ | _01986_;
	assign _04130_ = \mchip.index [11] & ~_04129_;
	assign _04131_ = _07835_ | \mchip.index [7];
	assign _04132_ = _04131_ | \mchip.index [8];
	assign _04133_ = _07758_ & ~_04132_;
	assign _04134_ = _00689_ & ~\mchip.index [10];
	assign _04135_ = _04382_ | \mchip.index [4];
	assign _04136_ = _04135_ | \mchip.index [5];
	assign _04137_ = _04136_ | _02984_;
	assign _04139_ = _04137_ | _02097_;
	assign _04140_ = _04139_ | \mchip.index [8];
	assign _04141_ = _04140_ | \mchip.index [9];
	assign _04142_ = \mchip.index [11] & ~_04141_;
	assign _04143_ = _07769_ | \mchip.index [4];
	assign _04144_ = _04143_ | \mchip.index [5];
	assign _04145_ = _04144_ | \mchip.index [6];
	assign _04146_ = _04145_ | _02097_;
	assign _04147_ = _04146_ | \mchip.index [8];
	assign _04148_ = _04147_ | \mchip.index [9];
	assign _04150_ = \mchip.index [10] & ~_04148_;
	assign _04151_ = _02051_ | _04648_;
	assign _04152_ = \mchip.index [11] & ~_04151_;
	assign _04153_ = _07715_ | _04648_;
	assign _04154_ = _04153_ | \mchip.index [9];
	assign _04155_ = \mchip.index [10] & ~_04154_;
	assign _04156_ = _00261_ | \mchip.index [7];
	assign _04157_ = _04156_ | _04648_;
	assign _04158_ = _04157_ | \mchip.index [10];
	assign _04159_ = _01875_ & ~_04158_;
	assign _04161_ = _02718_ | \mchip.index [7];
	assign _04162_ = _04161_ | _07758_;
	assign _04163_ = _01986_ & ~_04162_;
	assign _04164_ = _07864_ | _02097_;
	assign _04165_ = _04164_ | \mchip.index [8];
	assign _04166_ = _04165_ | _07758_;
	assign _04167_ = _01986_ & ~_04166_;
	assign _04168_ = _01364_ | _07758_;
	assign _04169_ = \mchip.index [11] & ~_04168_;
	assign _04170_ = _03110_ | _02097_;
	assign _04172_ = _04170_ | \mchip.index [9];
	assign _04173_ = _01986_ & ~_04172_;
	assign _04174_ = _02718_ | _02097_;
	assign _04175_ = _04174_ | \mchip.index [9];
	assign _04176_ = \mchip.index [11] & ~_04175_;
	assign _04177_ = _04249_ | \mchip.index [6];
	assign _04178_ = _04177_ | \mchip.index [8];
	assign _04179_ = _04178_ | \mchip.index [9];
	assign _04180_ = _04179_ | \mchip.index [10];
	assign _04181_ = _01875_ & ~_04180_;
	assign _04183_ = _01501_ | \mchip.index [5];
	assign _04184_ = _04183_ | _02984_;
	assign _04185_ = _04184_ | \mchip.index [7];
	assign _04186_ = _04185_ | _07758_;
	assign _04187_ = \mchip.index [11] & ~_04186_;
	assign _04188_ = _01232_ | _05424_;
	assign _04189_ = _04188_ | \mchip.index [6];
	assign _04190_ = _02097_ & ~_04189_;
	assign _04191_ = _02890_ | _02097_;
	assign _04192_ = _04191_ | _07758_;
	assign _04194_ = _01986_ & ~_04192_;
	assign _04195_ = _03869_ | \mchip.index [6];
	assign _04196_ = _04195_ | _02097_;
	assign _04197_ = _04196_ | \mchip.index [8];
	assign _04198_ = _04197_ | _07758_;
	assign _04199_ = \mchip.index [11] & ~_04198_;
	assign _04200_ = _00785_ | _02097_;
	assign _04201_ = _04200_ | \mchip.index [9];
	assign _04202_ = \mchip.index [11] & ~_04201_;
	assign _04203_ = _02167_ | \mchip.index [7];
	assign _04206_ = _04203_ | \mchip.index [8];
	assign _04207_ = _07758_ & ~_04206_;
	assign _04208_ = _03033_ | \mchip.index [9];
	assign _04209_ = \mchip.index [11] & ~_04208_;
	assign _04210_ = _01155_ | _04648_;
	assign _04211_ = \mchip.index [11] & ~_04210_;
	assign _04212_ = _01245_ | \mchip.index [8];
	assign _04213_ = _07758_ & ~_04212_;
	assign _04214_ = _02932_ | _01986_;
	assign _04215_ = \mchip.index [11] & ~_04214_;
	assign _04217_ = _00945_ | _02097_;
	assign _04218_ = _04217_ | \mchip.index [8];
	assign _04219_ = _04218_ | \mchip.index [9];
	assign _04220_ = _04219_ | _01986_;
	assign _04221_ = _01875_ & ~_04220_;
	assign _04222_ = _02364_ | _02984_;
	assign _04223_ = _04222_ | \mchip.index [8];
	assign _04224_ = _04223_ | _07758_;
	assign _04225_ = \mchip.index [11] & ~_04224_;
	assign _04226_ = _00822_ | \mchip.index [7];
	assign _04228_ = _04226_ | \mchip.index [8];
	assign _04229_ = _04228_ | \mchip.index [9];
	assign _04230_ = \mchip.index [11] & ~_04229_;
	assign _04231_ = _01105_ | \mchip.index [7];
	assign _04232_ = \mchip.index [11] & ~_04231_;
	assign _04233_ = _05347_ | _04648_;
	assign _04234_ = _04233_ | \mchip.index [9];
	assign _04235_ = _04234_ | \mchip.index [10];
	assign _04236_ = _01875_ & ~_04235_;
	assign _04237_ = _01147_ | \mchip.index [6];
	assign _04239_ = _04237_ | _04648_;
	assign _04240_ = _04239_ | _07758_;
	assign _04241_ = _01875_ & ~_04240_;
	assign _04242_ = _00869_ | _02097_;
	assign _04243_ = _04242_ | _01986_;
	assign _04244_ = \mchip.index [11] & ~_04243_;
	assign _04245_ = _01528_ | \mchip.index [9];
	assign _04246_ = _04245_ | _01986_;
	assign _04247_ = _01875_ & ~_04246_;
	assign _04248_ = _01986_ & ~_01735_;
	assign _04250_ = _01905_ | _04648_;
	assign _04251_ = _01875_ & ~_04250_;
	assign _04252_ = _07658_ | \mchip.index [6];
	assign _04253_ = _04252_ | _02097_;
	assign _04254_ = _04253_ | _04648_;
	assign _04255_ = \mchip.index [10] & ~_04254_;
	assign _04256_ = _00715_ | \mchip.index [8];
	assign _04257_ = _04256_ | \mchip.index [9];
	assign _04258_ = _04257_ | \mchip.index [10];
	assign _04259_ = _01875_ & ~_04258_;
	assign _04261_ = _00479_ | \mchip.index [8];
	assign _04262_ = \mchip.index [9] & ~_04261_;
	assign _04263_ = _01573_ | _04648_;
	assign _04264_ = _04263_ | _07758_;
	assign _04265_ = _04264_ | _01986_;
	assign _04266_ = _01875_ & ~_04265_;
	assign _04267_ = _02823_ | \mchip.index [9];
	assign _04268_ = \mchip.index [10] & ~_04267_;
	assign _04269_ = _01451_ | \mchip.index [8];
	assign _04270_ = _04269_ | _07758_;
	assign _04272_ = _01986_ & ~_04270_;
	assign _04273_ = _01438_ | \mchip.index [7];
	assign _04274_ = _04273_ | _04648_;
	assign _04275_ = \mchip.index [11] & ~_04274_;
	assign _04276_ = _01290_ | \mchip.index [7];
	assign _04277_ = _04276_ | _04648_;
	assign _04278_ = _04277_ | _07758_;
	assign _04279_ = _01986_ & ~_04278_;
	assign _04280_ = _07783_ | \mchip.index [7];
	assign _04281_ = _04280_ | \mchip.index [8];
	assign _04283_ = \mchip.index [11] & ~_04281_;
	assign _04284_ = _01983_ | \mchip.index [8];
	assign _04285_ = _04284_ | \mchip.index [9];
	assign _04286_ = \mchip.index [11] & ~_04285_;
	assign _04287_ = _02890_ | \mchip.index [6];
	assign _04288_ = _04287_ | \mchip.index [8];
	assign _04289_ = \mchip.index [11] & ~_04288_;
	assign _04290_ = _07714_ | \mchip.index [4];
	assign _04291_ = _04290_ | \mchip.index [5];
	assign _04292_ = _04291_ | \mchip.index [6];
	assign _04294_ = _04292_ | _04648_;
	assign _04295_ = _04294_ | \mchip.index [9];
	assign _04296_ = \mchip.index [11] & ~_04295_;
	assign _04297_ = _04031_ | \mchip.index [7];
	assign _04298_ = _04297_ | \mchip.index [8];
	assign _04299_ = \mchip.index [10] & ~_04298_;
	assign _04300_ = _07750_ | _04648_;
	assign _04301_ = _04300_ | _07758_;
	assign _04302_ = _04301_ | _01986_;
	assign _04303_ = _01875_ & ~_04302_;
	assign _04305_ = _01325_ | _02097_;
	assign _04306_ = _04305_ | _04648_;
	assign _04307_ = _04306_ | _07758_;
	assign _04308_ = _04307_ | _01986_;
	assign _04309_ = _01875_ & ~_04308_;
	assign _04310_ = _01178_ | \mchip.index [6];
	assign _04311_ = _04310_ | _02097_;
	assign _04312_ = _04311_ | _04648_;
	assign _04313_ = _01875_ & ~_04312_;
	assign _04314_ = _00255_ | \mchip.index [7];
	assign _04317_ = _04314_ | \mchip.index [8];
	assign _04318_ = _04317_ | \mchip.index [10];
	assign _04319_ = _01875_ & ~_04318_;
	assign _04320_ = _00320_ | \mchip.index [6];
	assign _04321_ = _04320_ | _02097_;
	assign _04322_ = _04321_ | \mchip.index [8];
	assign _04323_ = _04322_ | _07758_;
	assign _04324_ = \mchip.index [11] & ~_04323_;
	assign _04325_ = _04006_ | _02984_;
	assign _04326_ = _04325_ | \mchip.index [7];
	assign _04328_ = _04326_ | _07758_;
	assign _04329_ = _01986_ & ~_04328_;
	assign _04330_ = \mchip.index [11] & ~_02952_;
	assign _04331_ = _01924_ | _04648_;
	assign _04332_ = _04331_ | \mchip.index [10];
	assign _04333_ = \mchip.index [11] & ~_04332_;
	assign _04334_ = _00566_ | _02984_;
	assign _04335_ = _04334_ | \mchip.index [7];
	assign _04336_ = _04335_ | _04648_;
	assign _04337_ = _04336_ | \mchip.index [9];
	assign _04339_ = \mchip.index [11] & ~_04337_;
	assign _04340_ = _06135_ | \mchip.index [5];
	assign _04341_ = _04340_ | _02097_;
	assign _04342_ = _04341_ | _04648_;
	assign _04343_ = _04342_ | \mchip.index [9];
	assign _04344_ = \mchip.index [10] & ~_04343_;
	assign _04345_ = _01510_ | \mchip.index [8];
	assign _04346_ = _04345_ | \mchip.index [9];
	assign _04347_ = _01875_ & ~_04346_;
	assign _04348_ = _01742_ | \mchip.index [6];
	assign _04350_ = _04348_ | \mchip.index [7];
	assign _04351_ = _04350_ | _04648_;
	assign _04352_ = \mchip.index [11] & ~_04351_;
	assign _04353_ = _00430_ | \mchip.index [7];
	assign _04354_ = _04353_ | _04648_;
	assign _04355_ = \mchip.index [10] & ~_04354_;
	assign _04356_ = _03944_ | \mchip.index [8];
	assign _04357_ = _04356_ | \mchip.index [9];
	assign _04358_ = \mchip.index [11] & ~_04357_;
	assign _04359_ = _03244_ | \mchip.index [9];
	assign _04361_ = _04359_ | \mchip.index [10];
	assign _04362_ = _01875_ & ~_04361_;
	assign _04363_ = _00633_ | _07758_;
	assign _04364_ = _01875_ & ~_04363_;
	assign _04365_ = _03454_ | _02984_;
	assign _04366_ = _04365_ | \mchip.index [8];
	assign _04367_ = _01875_ & ~_04366_;
	assign _04368_ = _00476_ | \mchip.index [7];
	assign _04369_ = _04368_ | _07758_;
	assign _04370_ = _04369_ | _01986_;
	assign _04372_ = _01875_ & ~_04370_;
	assign _04373_ = _00856_ | \mchip.index [7];
	assign _04374_ = _04373_ | \mchip.index [8];
	assign _04375_ = _04374_ | _07758_;
	assign _04376_ = \mchip.index [10] & ~_04375_;
	assign _04377_ = _04237_ | _07758_;
	assign _04378_ = _04377_ | \mchip.index [10];
	assign _04379_ = _01875_ & ~_04378_;
	assign _04380_ = _03785_ | \mchip.index [8];
	assign _04381_ = _01986_ & ~_04380_;
	assign _04383_ = _02510_ | \mchip.index [7];
	assign _04384_ = _04383_ | _04648_;
	assign _04385_ = _04384_ | \mchip.index [9];
	assign _04386_ = \mchip.index [10] & ~_04385_;
	assign _04387_ = _01818_ | _04648_;
	assign _04388_ = _04387_ | \mchip.index [9];
	assign _04389_ = _01986_ & ~_04388_;
	assign _04390_ = _01391_ | \mchip.index [10];
	assign _04391_ = _01875_ & ~_04390_;
	assign _04392_ = _03200_ | \mchip.index [6];
	assign _04394_ = _04392_ | \mchip.index [8];
	assign _04395_ = _04394_ | \mchip.index [9];
	assign _04396_ = \mchip.index [10] & ~_04395_;
	assign _04397_ = _01320_ | \mchip.index [5];
	assign _04398_ = _04397_ | _02984_;
	assign _04399_ = _04398_ | _02097_;
	assign _04400_ = _04399_ | _01986_;
	assign _04401_ = \mchip.index [11] & ~_04400_;
	assign _04402_ = _01272_ | \mchip.index [6];
	assign _04403_ = \mchip.index [11] & ~_04402_;
	assign _04405_ = _01166_ | \mchip.index [7];
	assign _04406_ = _04405_ | _07758_;
	assign _04407_ = \mchip.index [11] & ~_04406_;
	assign _04408_ = _01708_ | _02097_;
	assign _04409_ = _04408_ | \mchip.index [8];
	assign _04410_ = _04409_ | _07758_;
	assign _04411_ = _04410_ | _01986_;
	assign _04412_ = _01875_ & ~_04411_;
	assign _04413_ = _05070_ | \mchip.index [8];
	assign _04414_ = _04413_ | \mchip.index [10];
	assign _04416_ = _01875_ & ~_04414_;
	assign _04417_ = _00398_ | \mchip.index [8];
	assign _04418_ = _04417_ | \mchip.index [9];
	assign _04419_ = \mchip.index [10] & ~_04418_;
	assign _04420_ = _00255_ | _02097_;
	assign _04421_ = _04420_ | \mchip.index [8];
	assign _04422_ = _04421_ | _07758_;
	assign _04423_ = \mchip.index [10] & ~_04422_;
	assign _04424_ = _03115_ | _02984_;
	assign _04425_ = _04424_ | _02097_;
	assign _04428_ = _04425_ | \mchip.index [8];
	assign _04429_ = _04428_ | \mchip.index [9];
	assign _04430_ = \mchip.index [10] & ~_04429_;
	assign _04431_ = _07774_ | \mchip.index [8];
	assign _04432_ = _07758_ & ~_04431_;
	assign _04433_ = _04759_ | _02984_;
	assign _04434_ = _04433_ | _02097_;
	assign _04435_ = _04434_ | _04648_;
	assign _04436_ = _04435_ | \mchip.index [9];
	assign _04437_ = \mchip.index [10] & ~_04436_;
	assign _04439_ = _02192_ | _02097_;
	assign _04440_ = _04439_ | _04648_;
	assign _04441_ = _04440_ | \mchip.index [10];
	assign _04442_ = \mchip.index [11] & ~_04441_;
	assign _04443_ = _07199_ | \mchip.index [7];
	assign _04444_ = _04443_ | _04648_;
	assign _04445_ = _04444_ | \mchip.index [9];
	assign _04446_ = _04445_ | \mchip.index [10];
	assign _04447_ = _01875_ & ~_04446_;
	assign _04448_ = _03773_ | _02097_;
	assign _04450_ = _04448_ | _04648_;
	assign _04451_ = _04450_ | _07758_;
	assign _04452_ = _01875_ & ~_04451_;
	assign _04453_ = _02810_ | _07758_;
	assign _04454_ = _01986_ & ~_04453_;
	assign _04455_ = _00516_ | \mchip.index [7];
	assign _04456_ = _04455_ | \mchip.index [9];
	assign _04457_ = _04456_ | \mchip.index [10];
	assign _04458_ = _01875_ & ~_04457_;
	assign _04459_ = _01343_ | \mchip.index [6];
	assign _04461_ = _04459_ | _04648_;
	assign _04462_ = _04461_ | \mchip.index [10];
	assign _04463_ = _01875_ & ~_04462_;
	assign _04464_ = _01562_ | _02097_;
	assign _04465_ = _04464_ | \mchip.index [8];
	assign _04466_ = _04465_ | \mchip.index [9];
	assign _04467_ = \mchip.index [10] & ~_04466_;
	assign _04468_ = _07835_ | \mchip.index [9];
	assign _04469_ = _04468_ | \mchip.index [10];
	assign _04470_ = _01875_ & ~_04469_;
	assign _04472_ = _02430_ | \mchip.index [6];
	assign _04473_ = _04472_ | \mchip.index [7];
	assign _04474_ = _04473_ | _04648_;
	assign _04475_ = _04474_ | _07758_;
	assign _04476_ = _01986_ & ~_04475_;
	assign _04477_ = _02167_ | \mchip.index [8];
	assign _04478_ = \mchip.index [10] & ~_04477_;
	assign _04479_ = _02149_ | \mchip.index [9];
	assign _04480_ = \mchip.index [10] & ~_04479_;
	assign _04481_ = _02797_ | \mchip.index [8];
	assign _04483_ = _07758_ & ~_04481_;
	assign _04484_ = _03110_ | _02984_;
	assign _04485_ = _04484_ | _04648_;
	assign _04486_ = _04485_ | \mchip.index [10];
	assign _04487_ = _01875_ & ~_04486_;
	assign _04488_ = _06346_ | _02097_;
	assign _04489_ = _04488_ | _07758_;
	assign _04490_ = \mchip.index [11] & ~_04489_;
	assign _04491_ = _00433_ | _02097_;
	assign _04492_ = _04491_ | _04648_;
	assign _04494_ = _04492_ | \mchip.index [9];
	assign _04495_ = \mchip.index [10] & ~_04494_;
	assign _04496_ = _02944_ | _07758_;
	assign _04497_ = _01986_ & ~_04496_;
	assign _04498_ = _05946_ | \mchip.index [6];
	assign _04499_ = _04498_ | _02097_;
	assign _04500_ = _04499_ | \mchip.index [8];
	assign _04501_ = _04500_ | _07758_;
	assign _04502_ = _01986_ & ~_04501_;
	assign _04503_ = _01986_ & ~_03059_;
	assign _04505_ = _02823_ | _04648_;
	assign _04506_ = _04505_ | _01986_;
	assign _04507_ = _01875_ & ~_04506_;
	assign _04508_ = _01242_ | _02984_;
	assign _04509_ = _04508_ | _04648_;
	assign _04510_ = _04509_ | \mchip.index [9];
	assign _04511_ = \mchip.index [10] & ~_04510_;
	assign _04512_ = _03035_ | _02097_;
	assign _04513_ = _04512_ | \mchip.index [8];
	assign _04514_ = _04513_ | \mchip.index [9];
	assign _04516_ = _01986_ & ~_04514_;
	assign _04517_ = _01509_ | \mchip.index [6];
	assign _04518_ = _04517_ | \mchip.index [8];
	assign _04519_ = _04518_ | \mchip.index [9];
	assign _04520_ = _04519_ | \mchip.index [10];
	assign _04521_ = _01875_ & ~_04520_;
	assign _04522_ = _01742_ | _02984_;
	assign _04523_ = _04522_ | _02097_;
	assign _04524_ = _04523_ | _07758_;
	assign _04525_ = \mchip.index [10] & ~_04524_;
	assign _04527_ = _01105_ | _07758_;
	assign _04528_ = \mchip.index [11] & ~_04527_;
	assign _04529_ = _02375_ | \mchip.index [7];
	assign _04530_ = _04529_ | \mchip.index [8];
	assign _04531_ = _04530_ | _07758_;
	assign _04532_ = \mchip.index [10] & ~_04531_;
	assign _04533_ = _04276_ | \mchip.index [8];
	assign _04534_ = _04533_ | \mchip.index [9];
	assign _04535_ = \mchip.index [10] & ~_04534_;
	assign _04536_ = _02364_ | \mchip.index [8];
	assign _04539_ = _04536_ | \mchip.index [9];
	assign _04540_ = _04539_ | \mchip.index [10];
	assign _04541_ = _01875_ & ~_04540_;
	assign _04542_ = _07666_ | \mchip.index [8];
	assign _04543_ = _04542_ | \mchip.index [10];
	assign _04544_ = _01875_ & ~_04543_;
	assign _04545_ = _02021_ | _02097_;
	assign _04546_ = _04545_ | \mchip.index [8];
	assign _04547_ = \mchip.index [9] & ~_04546_;
	assign _04548_ = _03971_ | \mchip.index [6];
	assign _04550_ = _04548_ | \mchip.index [7];
	assign _04551_ = _04550_ | _01986_;
	assign _04552_ = \mchip.index [11] & ~_04551_;
	assign _04553_ = _07721_ | \mchip.index [7];
	assign _04554_ = _04553_ | \mchip.index [8];
	assign _04555_ = _04554_ | \mchip.index [9];
	assign _04556_ = \mchip.index [10] & ~_04555_;
	assign _04557_ = _03932_ | \mchip.index [7];
	assign _04558_ = _04557_ | \mchip.index [8];
	assign _04559_ = _04558_ | \mchip.index [9];
	assign _04561_ = _01875_ & ~_04559_;
	assign _04562_ = _01190_ | _04648_;
	assign _04563_ = _04562_ | \mchip.index [9];
	assign _04564_ = _01986_ & ~_04563_;
	assign _04565_ = _02609_ | \mchip.index [10];
	assign _04566_ = \mchip.index [11] & ~_04565_;
	assign _04567_ = _02161_ | \mchip.index [8];
	assign _04568_ = _04567_ | _07758_;
	assign _04569_ = \mchip.index [10] & ~_04568_;
	assign _04570_ = \mchip.index [10] & ~_03999_;
	assign _04572_ = _00670_ | \mchip.index [7];
	assign _04573_ = _04572_ | \mchip.index [8];
	assign _04574_ = _04573_ | \mchip.index [9];
	assign _04575_ = \mchip.index [10] & ~_04574_;
	assign _04576_ = _07839_ | \mchip.index [5];
	assign _04577_ = _04576_ | _02984_;
	assign _04578_ = _04577_ | _02097_;
	assign _04579_ = _04578_ | _07758_;
	assign _04580_ = _01986_ & ~_04579_;
	assign _04581_ = _03454_ | \mchip.index [7];
	assign _04583_ = _07758_ & ~_04581_;
	assign _04584_ = \mchip.index [11] & ~_01474_;
	assign _04585_ = _01422_ | _02097_;
	assign _04586_ = _04585_ | _04648_;
	assign _04587_ = _04586_ | \mchip.index [9];
	assign _04588_ = _01875_ & ~_04587_;
	assign _04589_ = _03860_ | \mchip.index [6];
	assign _04590_ = _04589_ | \mchip.index [7];
	assign _04591_ = _04590_ | \mchip.index [9];
	assign _04592_ = _04591_ | \mchip.index [10];
	assign _04594_ = _01875_ & ~_04592_;
	assign _04595_ = _01457_ | \mchip.index [8];
	assign _04596_ = _04595_ | \mchip.index [9];
	assign _04597_ = \mchip.index [10] & ~_04596_;
	assign _04598_ = _02495_ | \mchip.index [7];
	assign _04599_ = _04598_ | _04648_;
	assign _04600_ = _07758_ & ~_04599_;
	assign _04601_ = _02661_ | \mchip.index [6];
	assign _04602_ = _04601_ | \mchip.index [7];
	assign _04603_ = _04602_ | _04648_;
	assign _04605_ = \mchip.index [10] & ~_04603_;
	assign _04606_ = _01548_ | \mchip.index [7];
	assign _04607_ = _07758_ & ~_04606_;
	assign _04608_ = _00255_ | \mchip.index [5];
	assign _04609_ = _04608_ | _02984_;
	assign _04610_ = _04609_ | \mchip.index [7];
	assign _04611_ = _04610_ | _01986_;
	assign _04612_ = \mchip.index [11] & ~_04611_;
	assign _04613_ = _01641_ | \mchip.index [7];
	assign _04614_ = _04613_ | _01986_;
	assign _04616_ = \mchip.index [11] & ~_04614_;
	assign _04617_ = _04205_ | _05424_;
	assign _04618_ = _04617_ | \mchip.index [6];
	assign _04619_ = _04618_ | _02097_;
	assign _04620_ = _04619_ | _07758_;
	assign _04621_ = \mchip.index [11] & ~_04620_;
	assign _04622_ = _01748_ | _02984_;
	assign _04623_ = _04622_ | \mchip.index [7];
	assign _04624_ = \mchip.index [10] & ~_04623_;
	assign _04625_ = \mchip.index [10] & ~_03442_;
	assign _04627_ = _01427_ | \mchip.index [7];
	assign _04628_ = _04627_ | _04648_;
	assign _04629_ = _04628_ | \mchip.index [9];
	assign _04630_ = \mchip.index [11] & ~_04629_;
	assign _04631_ = _00463_ | _02984_;
	assign _04632_ = _04631_ | \mchip.index [7];
	assign _04633_ = _04632_ | _04648_;
	assign _04634_ = _04633_ | \mchip.index [9];
	assign _04635_ = _01875_ & ~_04634_;
	assign _04636_ = _01929_ | _04648_;
	assign _04638_ = \mchip.index [10] & ~_04636_;
	assign _04639_ = _06135_ | _02984_;
	assign _04640_ = _04639_ | \mchip.index [7];
	assign _04641_ = _04640_ | _04648_;
	assign _04642_ = _04641_ | \mchip.index [9];
	assign _04643_ = _04642_ | \mchip.index [10];
	assign _04644_ = _01875_ & ~_04643_;
	assign _04645_ = _04682_ | _02984_;
	assign _04646_ = _04645_ | _02097_;
	assign _04647_ = _04646_ | _04648_;
	assign _04650_ = _04647_ | _07758_;
	assign _04651_ = _01986_ & ~_04650_;
	assign _04652_ = _01710_ | \mchip.index [7];
	assign _04653_ = _04652_ | _07758_;
	assign _04654_ = _04653_ | _01986_;
	assign _04655_ = _01875_ & ~_04654_;
	assign _04656_ = _02724_ | _02097_;
	assign _04657_ = _04656_ | \mchip.index [9];
	assign _04658_ = _01875_ & ~_04657_;
	assign _04659_ = _01153_ | _01986_;
	assign _04661_ = \mchip.index [11] & ~_04659_;
	assign _04662_ = _01133_ | _07758_;
	assign _04663_ = _04662_ | \mchip.index [10];
	assign _04664_ = \mchip.index [11] & ~_04663_;
	assign _04665_ = _00366_ | _02984_;
	assign _04666_ = _04665_ | _02097_;
	assign _04667_ = _04666_ | _04648_;
	assign _04668_ = _04667_ | \mchip.index [9];
	assign _04669_ = _04668_ | \mchip.index [10];
	assign _04670_ = _01875_ & ~_04669_;
	assign _04672_ = _00887_ | \mchip.index [7];
	assign _04673_ = _04672_ | _01986_;
	assign _04674_ = \mchip.index [11] & ~_04673_;
	assign _04675_ = \mchip.index [5] & ~_03860_;
	assign _04676_ = _03304_ & ~_01875_;
	assign _04677_ = _02439_ | _02097_;
	assign _04678_ = _04677_ | \mchip.index [9];
	assign _04679_ = \mchip.index [10] & ~_04678_;
	assign _04680_ = _01428_ | _02097_;
	assign _04681_ = _04680_ | _07758_;
	assign _04683_ = \mchip.index [10] & ~_04681_;
	assign _04684_ = _01503_ | \mchip.index [8];
	assign _04685_ = _04684_ | \mchip.index [9];
	assign _04686_ = \mchip.index [11] & ~_04685_;
	assign _04687_ = _07758_ & ~_04288_;
	assign _04688_ = _01600_ | _04648_;
	assign _04689_ = _04688_ | \mchip.index [9];
	assign _04690_ = \mchip.index [11] & ~_04689_;
	assign _04691_ = _02031_ | \mchip.index [6];
	assign _04692_ = _04691_ | _02097_;
	assign _04694_ = _04692_ | \mchip.index [8];
	assign _04695_ = \mchip.index [11] & ~_04694_;
	assign _04696_ = _02996_ | _04648_;
	assign _04697_ = _04696_ | \mchip.index [9];
	assign _04698_ = \mchip.index [10] & ~_04697_;
	assign _04699_ = _00505_ | \mchip.index [6];
	assign _04700_ = _04699_ | _02097_;
	assign _04701_ = _04700_ | _04648_;
	assign _04702_ = _04701_ | \mchip.index [9];
	assign _04703_ = \mchip.index [11] & ~_04702_;
	assign _04705_ = _07721_ | _05424_;
	assign _04706_ = \mchip.index [11] & ~_04705_;
	assign _04707_ = _07768_ | _02097_;
	assign _04708_ = _04707_ | _04648_;
	assign _04709_ = _04708_ | _07758_;
	assign _04710_ = _04709_ | _01986_;
	assign _04711_ = _01875_ & ~_04710_;
	assign _04712_ = _04193_ | _02984_;
	assign _04713_ = _04712_ | \mchip.index [7];
	assign _04714_ = _04713_ | _04648_;
	assign _04716_ = _04714_ | \mchip.index [9];
	assign _04717_ = _04716_ | \mchip.index [10];
	assign _04718_ = _01875_ & ~_04717_;
	assign _04719_ = _04522_ | _04648_;
	assign _04720_ = \mchip.index [9] & ~_04719_;
	assign _04721_ = _00837_ | _04648_;
	assign _04722_ = _04721_ | \mchip.index [10];
	assign _04723_ = _01875_ & ~_04722_;
	assign _04724_ = _02017_ | _01986_;
	assign _04725_ = _01875_ & ~_04724_;
	assign _04727_ = _07840_ | \mchip.index [8];
	assign _04728_ = _04727_ | _07758_;
	assign _04729_ = \mchip.index [11] & ~_04728_;
	assign _04730_ = _00632_ | _02097_;
	assign _04731_ = _04730_ | \mchip.index [8];
	assign _04732_ = _04731_ | \mchip.index [9];
	assign _04733_ = _01986_ & ~_04732_;
	assign _04734_ = _01208_ | \mchip.index [9];
	assign _04735_ = _04734_ | \mchip.index [10];
	assign _04736_ = _01875_ & ~_04735_;
	assign _04738_ = _07793_ | _04648_;
	assign _04739_ = _04738_ | \mchip.index [9];
	assign _04740_ = _01986_ & ~_04739_;
	assign _04741_ = _00560_ | \mchip.index [4];
	assign _04742_ = _04741_ | \mchip.index [5];
	assign _04743_ = _04742_ | \mchip.index [6];
	assign _04744_ = _04743_ | _02097_;
	assign _04745_ = _04744_ | _07758_;
	assign _04746_ = _04745_ | \mchip.index [10];
	assign _04747_ = _01875_ & ~_04746_;
	assign _04749_ = _00868_ & ~_01875_;
	assign _04750_ = _05048_ | _05424_;
	assign _04751_ = _01986_ & ~_04750_;
	assign _04752_ = _03371_ | _02097_;
	assign _04753_ = _04752_ | _07758_;
	assign _04754_ = _04753_ | _01986_;
	assign _04755_ = _01875_ & ~_04754_;
	assign _04756_ = _01389_ | _02984_;
	assign _04757_ = _04756_ | _02097_;
	assign _04758_ = _04757_ | \mchip.index [10];
	assign _04761_ = \mchip.index [11] & ~_04758_;
	assign _04762_ = _02960_ | \mchip.index [6];
	assign _04763_ = _04762_ | \mchip.index [7];
	assign _04764_ = _04763_ | _04648_;
	assign _04765_ = _04764_ | _01986_;
	assign _04766_ = _01875_ & ~_04765_;
	assign _04767_ = _03325_ | \mchip.index [8];
	assign _04768_ = \mchip.index [11] & ~_04767_;
	assign _04769_ = _02884_ | \mchip.index [8];
	assign _04770_ = _04769_ | _07758_;
	assign _04772_ = \mchip.index [10] & ~_04770_;
	assign _04773_ = _04593_ | _04648_;
	assign _04774_ = _04773_ | \mchip.index [9];
	assign _04775_ = \mchip.index [10] & ~_04774_;
	assign _04776_ = _04775_ | _04772_;
	assign _04777_ = _04776_ | _04768_;
	assign _04778_ = _04777_ | _04766_;
	assign _04779_ = _04778_ | _04761_;
	assign _04780_ = _04779_ | _04755_;
	assign _04781_ = _04780_ | _04751_;
	assign _04783_ = _04781_ | _04749_;
	assign _04784_ = _04783_ | _04747_;
	assign _04785_ = _04784_ | _04740_;
	assign _04786_ = _04785_ | _04736_;
	assign _04787_ = _04786_ | _04733_;
	assign _04788_ = _04787_ | _04729_;
	assign _04789_ = _04788_ | _04725_;
	assign _04790_ = _04789_ | _04723_;
	assign _04791_ = _04790_ | _04720_;
	assign _04792_ = _04791_ | _04718_;
	assign _04794_ = _04792_ | _04711_;
	assign _04795_ = _04794_ | _04706_;
	assign _04796_ = _04795_ | _04703_;
	assign _04797_ = _04796_ | _04698_;
	assign _04798_ = _04797_ | _04695_;
	assign _04799_ = _04798_ | _04690_;
	assign _04800_ = _04799_ | _04687_;
	assign _04801_ = _04800_ | _04686_;
	assign _04802_ = _04801_ | _04683_;
	assign _04803_ = _04802_ | _04679_;
	assign _04805_ = _04803_ | _04676_;
	assign _04806_ = _04805_ | _04675_;
	assign _04807_ = _04806_ | _03375_;
	assign _04808_ = _04807_ | _04674_;
	assign _04809_ = _04808_ | _04670_;
	assign _04810_ = _04809_ | _04664_;
	assign _04811_ = _04810_ | _04661_;
	assign _04812_ = _04811_ | _03366_;
	assign _04813_ = _04812_ | _04658_;
	assign _04814_ = _04813_ | _04655_;
	assign _04816_ = _04814_ | _04651_;
	assign _04817_ = _04816_ | _04644_;
	assign _04818_ = _04817_ | _04638_;
	assign _04819_ = _04818_ | _04635_;
	assign _04820_ = _04819_ | _04630_;
	assign _04821_ = _04820_ | _04625_;
	assign _04822_ = _04821_ | _04624_;
	assign _04823_ = _04822_ | _04621_;
	assign _04824_ = _04823_ | _04616_;
	assign _04825_ = _04824_ | _04612_;
	assign _04827_ = _04825_ | _04607_;
	assign _04828_ = _04827_ | _04605_;
	assign _04829_ = _04828_ | _04600_;
	assign _04830_ = _04829_ | _04597_;
	assign _04831_ = _04830_ | _04594_;
	assign _04832_ = _04831_ | _04588_;
	assign _04833_ = _04832_ | _04584_;
	assign _04834_ = _04833_ | _04583_;
	assign _04835_ = _04834_ | _04580_;
	assign _04836_ = _04835_ | _04575_;
	assign _04838_ = _04836_ | _01999_;
	assign _04839_ = _04838_ | _04570_;
	assign _04840_ = _04839_ | _04569_;
	assign _04841_ = _04840_ | _04566_;
	assign _04842_ = _04841_ | _04564_;
	assign _04843_ = _04842_ | _04561_;
	assign _04844_ = _04843_ | _04556_;
	assign _04845_ = _04844_ | _04552_;
	assign _04846_ = _04845_ | _04547_;
	assign _04847_ = _04846_ | _04544_;
	assign _04849_ = _04847_ | _04541_;
	assign _04850_ = _04849_ | _04535_;
	assign _04851_ = _04850_ | _04532_;
	assign _04852_ = _04851_ | _04528_;
	assign _04853_ = _04852_ | _04525_;
	assign _04854_ = _04853_ | _04521_;
	assign _04855_ = _04854_ | _04516_;
	assign _04856_ = _04855_ | _04511_;
	assign _04857_ = _04856_ | _04507_;
	assign _04858_ = _04857_ | _04503_;
	assign _04860_ = _04858_ | _04502_;
	assign _04861_ = _04860_ | _04497_;
	assign _04862_ = _04861_ | _04495_;
	assign _04863_ = _04862_ | _04490_;
	assign _04864_ = _04863_ | _04487_;
	assign _04865_ = _04864_ | _04483_;
	assign _04866_ = _04865_ | _04480_;
	assign _04867_ = _04866_ | _04478_;
	assign _04868_ = _04867_ | _04476_;
	assign _04869_ = _04868_ | _04470_;
	assign _04872_ = _04869_ | _04467_;
	assign _04873_ = _04872_ | _04463_;
	assign _04874_ = _04873_ | _04458_;
	assign _04875_ = _04874_ | _04454_;
	assign _04876_ = _04875_ | _04452_;
	assign _04877_ = _04876_ | _04447_;
	assign _04878_ = _04877_ | _04442_;
	assign _04879_ = _04878_ | _04437_;
	assign _04880_ = _04879_ | _04432_;
	assign _04881_ = _04880_ | _04430_;
	assign _04883_ = _04881_ | _04423_;
	assign _04884_ = _04883_ | _04419_;
	assign _04885_ = _04884_ | _04416_;
	assign _04886_ = _04885_ | _04412_;
	assign _04887_ = _04886_ | _04407_;
	assign _04888_ = _04887_ | _04403_;
	assign _04889_ = _04888_ | _04401_;
	assign _04890_ = _04889_ | _04396_;
	assign _04891_ = _04890_ | _04391_;
	assign _04892_ = _04891_ | _04389_;
	assign _04894_ = _04892_ | _04386_;
	assign _04895_ = _04894_ | _04381_;
	assign _04896_ = _04895_ | _04379_;
	assign _04897_ = _04896_ | _04376_;
	assign _04898_ = _04897_ | _04372_;
	assign _04899_ = _04898_ | _04367_;
	assign _04900_ = _04899_ | _04364_;
	assign _04901_ = _04900_ | _04362_;
	assign _04902_ = _04901_ | _04358_;
	assign _04903_ = _04902_ | _04355_;
	assign _04905_ = _04903_ | _04352_;
	assign _04906_ = _04905_ | _04347_;
	assign _04907_ = _04906_ | _04344_;
	assign _04908_ = _04907_ | _04339_;
	assign _04909_ = _04908_ | _03082_;
	assign _04910_ = _04909_ | _04333_;
	assign _04911_ = _04910_ | _04330_;
	assign _04912_ = _04911_ | _04329_;
	assign _04913_ = _04912_ | _04324_;
	assign _04914_ = _04913_ | _04319_;
	assign _04916_ = _04914_ | _04313_;
	assign _04917_ = _04916_ | _04309_;
	assign _04918_ = _04917_ | _04303_;
	assign _04919_ = _04918_ | _04299_;
	assign _04920_ = _04919_ | _04296_;
	assign _04921_ = _04920_ | _04289_;
	assign _04922_ = _04921_ | _04286_;
	assign _04923_ = _04922_ | _04283_;
	assign _04924_ = _04923_ | _04279_;
	assign _04925_ = _04924_ | _04275_;
	assign _04927_ = _04925_ | _04272_;
	assign _04928_ = _04927_ | _04268_;
	assign _04929_ = _04928_ | _04266_;
	assign _04930_ = _04929_ | _04262_;
	assign _04931_ = _04930_ | _04259_;
	assign _04932_ = _04931_ | _04255_;
	assign _04933_ = _04932_ | _04251_;
	assign _04934_ = _04933_ | _04248_;
	assign _04935_ = _04934_ | _04247_;
	assign _04936_ = _04935_ | _04244_;
	assign _04938_ = _04936_ | _02905_;
	assign _04939_ = _04938_ | _04241_;
	assign _04940_ = _04939_ | _04236_;
	assign _04941_ = _04940_ | _04232_;
	assign _04942_ = _04941_ | _04230_;
	assign _04943_ = _04942_ | _04225_;
	assign _04944_ = _04943_ | _04221_;
	assign _04945_ = _04944_ | _04215_;
	assign _04946_ = _04945_ | _04213_;
	assign _04947_ = _04946_ | _04211_;
	assign _04949_ = _04947_ | _04209_;
	assign _04950_ = _04949_ | _04207_;
	assign _04951_ = _04950_ | _04202_;
	assign _04952_ = _04951_ | _04199_;
	assign _04953_ = _04952_ | _04194_;
	assign _04954_ = _04953_ | _04190_;
	assign _04955_ = _04954_ | _04187_;
	assign _04956_ = _04955_ | _04181_;
	assign _04957_ = _04956_ | _04176_;
	assign _04958_ = _04957_ | _04173_;
	assign _04960_ = _04958_ | _04169_;
	assign _04961_ = _04960_ | _04167_;
	assign _04962_ = _04961_ | _04163_;
	assign _04963_ = _04962_ | _04159_;
	assign _04964_ = _04963_ | _04155_;
	assign _04965_ = _04964_ | _04152_;
	assign _04966_ = _04965_ | _04150_;
	assign _04967_ = _04966_ | _04142_;
	assign _04968_ = _04967_ | _04134_;
	assign _04969_ = _04968_ | _04133_;
	assign _04971_ = _04969_ | _04130_;
	assign _04972_ = _04971_ | _04128_;
	assign _04973_ = _04972_ | _04125_;
	assign _04974_ = _04973_ | _04120_;
	assign _04975_ = _04974_ | _04117_;
	assign _04976_ = _04975_ | _04112_;
	assign _04977_ = _04976_ | _02732_;
	assign _04978_ = _04977_ | _04109_;
	assign _04979_ = _04978_ | _04106_;
	assign _04980_ = _04979_ | _04103_;
	assign _04983_ = _04980_ | _04100_;
	assign _04984_ = _04983_ | _04097_;
	assign _04985_ = _04984_ | _04091_;
	assign _04986_ = _04985_ | _04088_;
	assign _04987_ = _04986_ | _04085_;
	assign _04988_ = _04987_ | _04080_;
	assign _04989_ = _04988_ | _04079_;
	assign _04990_ = _04989_ | _04077_;
	assign _04991_ = _04990_ | _04073_;
	assign _04992_ = _04991_ | _04069_;
	assign _04994_ = _04992_ | _04066_;
	assign _04995_ = _04994_ | _04063_;
	assign _04996_ = _04995_ | _04059_;
	assign _04997_ = _04996_ | _04054_;
	assign _04998_ = _04997_ | _04051_;
	assign _04999_ = _04998_ | _04050_;
	assign _05000_ = _04999_ | _04045_;
	assign _05001_ = _05000_ | _04044_;
	assign _05002_ = _05001_ | _04043_;
	assign _05003_ = _05002_ | _04037_;
	assign _05005_ = _05003_ | _04033_;
	assign _05006_ = _05005_ | _04030_;
	assign _05007_ = _05006_ | _04029_;
	assign _05008_ = _05007_ | _04025_;
	assign _05009_ = _05008_ | _04021_;
	assign _05010_ = _05009_ | _04020_;
	assign _05011_ = _05010_ | _02634_;
	assign _05012_ = _05011_ | _04015_;
	assign _05013_ = _05012_ | _04013_;
	assign _05014_ = _05013_ | _04010_;
	assign _05016_ = _05014_ | _04004_;
	assign _05017_ = _05016_ | _04000_;
	assign _05018_ = _05017_ | _03997_;
	assign _05019_ = _05018_ | _03995_;
	assign _05020_ = _05019_ | _03990_;
	assign _05021_ = _05020_ | _03987_;
	assign _05022_ = _05021_ | _03981_;
	assign _05023_ = _05022_ | _03976_;
	assign _05024_ = _05023_ | _03969_;
	assign _05025_ = _05024_ | _03965_;
	assign _05027_ = _05025_ | _03964_;
	assign _05028_ = _05027_ | _03959_;
	assign _05029_ = _05028_ | _03957_;
	assign _05030_ = _05029_ | _03953_;
	assign _05031_ = _05030_ | _03948_;
	assign _05032_ = _05031_ | _03942_;
	assign _05033_ = _05032_ | _03936_;
	assign _05034_ = _05033_ | _03931_;
	assign _05035_ = _05034_ | _03928_;
	assign _05036_ = _05035_ | _03925_;
	assign _05038_ = _05036_ | _03921_;
	assign _05039_ = _05038_ | _03919_;
	assign _05040_ = _05039_ | _03917_;
	assign _05041_ = _05040_ | _03913_;
	assign _05042_ = _05041_ | _03910_;
	assign _05043_ = _05042_ | _03904_;
	assign _05044_ = _05043_ | _03900_;
	assign _05045_ = _05044_ | _03896_;
	assign _05046_ = _05045_ | _03892_;
	assign _05047_ = _05046_ | _03891_;
	assign _05049_ = _05047_ | _03887_;
	assign _05050_ = _05049_ | _03884_;
	assign _05051_ = _05050_ | _03880_;
	assign _05052_ = _05051_ | _03876_;
	assign _05053_ = _05052_ | _03868_;
	assign _05054_ = _05053_ | _03862_;
	assign _05055_ = _05054_ | _03856_;
	assign _05056_ = _05055_ | _03853_;
	assign _05057_ = _05056_ | _03851_;
	assign _05058_ = _05057_ | _03846_;
	assign _05060_ = _05058_ | _03844_;
	assign _05061_ = _05060_ | _03841_;
	assign _05062_ = _05061_ | _03837_;
	assign _05063_ = _05062_ | _03834_;
	assign _05064_ = _05063_ | _03832_;
	assign _05065_ = _05064_ | _03830_;
	assign _05066_ = _05065_ | _03824_;
	assign _05067_ = _05066_ | _03820_;
	assign _05068_ = _05067_ | _03814_;
	assign _05069_ = _05068_ | _03810_;
	assign _05071_ = _05069_ | _03804_;
	assign _05072_ = _05071_ | _03801_;
	assign _05073_ = _05072_ | _03799_;
	assign _05074_ = _05073_ | _03797_;
	assign _05075_ = _05074_ | _03793_;
	assign _05076_ = _05075_ | _03791_;
	assign _05077_ = _05076_ | _03787_;
	assign _05078_ = _05077_ | _03782_;
	assign _05079_ = _05078_ | _03779_;
	assign _05080_ = _05079_ | _02448_;
	assign \mchip.val [2] = _05080_ | _03776_;
	assign _05082_ = _04666_ | \mchip.index [8];
	assign _05083_ = _05082_ | \mchip.index [9];
	assign _05084_ = _05083_ | \mchip.index [10];
	assign _05085_ = _01875_ & ~_05084_;
	assign _05086_ = _04656_ | _04648_;
	assign _05087_ = _05086_ | \mchip.index [9];
	assign _05088_ = _01875_ & ~_05087_;
	assign _05089_ = _01774_ | _02984_;
	assign _05090_ = _05089_ | _02097_;
	assign _05093_ = _05090_ | _07758_;
	assign _05094_ = _01986_ & ~_05093_;
	assign _05095_ = _02942_ | \mchip.index [7];
	assign _05096_ = _05095_ | \mchip.index [8];
	assign _05097_ = _05096_ | \mchip.index [9];
	assign _05098_ = _01986_ & ~_05097_;
	assign _05099_ = _02549_ | \mchip.index [8];
	assign _05100_ = _05099_ | \mchip.index [9];
	assign _05101_ = \mchip.index [10] & ~_05100_;
	assign _05102_ = _01399_ | _04648_;
	assign _05104_ = \mchip.index [11] & ~_05102_;
	assign _05105_ = _01387_ | _02097_;
	assign _05106_ = _05105_ | _04648_;
	assign _05107_ = _05106_ | \mchip.index [10];
	assign _05108_ = \mchip.index [11] & ~_05107_;
	assign _05109_ = \mchip.index [9] & ~_01800_;
	assign _05110_ = _01535_ | _04648_;
	assign _05111_ = _05110_ | \mchip.index [9];
	assign _05112_ = \mchip.index [10] & ~_05111_;
	assign _05113_ = _05868_ | \mchip.index [4];
	assign _05115_ = _05113_ | \mchip.index [5];
	assign _05116_ = _05115_ | _02984_;
	assign _05117_ = _05116_ | \mchip.index [7];
	assign _05118_ = _05117_ | \mchip.index [8];
	assign _05119_ = _05118_ | _07758_;
	assign _05120_ = \mchip.index [10] & ~_05119_;
	assign _05121_ = _07653_ | _05424_;
	assign _05122_ = _05121_ | _02984_;
	assign _05123_ = _05122_ | _02097_;
	assign _05124_ = _07758_ & ~_05123_;
	assign _05126_ = _07712_ | \mchip.index [6];
	assign _05127_ = _05126_ | _02097_;
	assign _05128_ = _05127_ | \mchip.index [8];
	assign _05129_ = _05128_ | _07758_;
	assign _05130_ = \mchip.index [10] & ~_05129_;
	assign _05131_ = _04380_ | \mchip.index [9];
	assign _05132_ = \mchip.index [11] & ~_05131_;
	assign _05133_ = _04522_ | \mchip.index [8];
	assign _05134_ = _05133_ | _07758_;
	assign _05135_ = \mchip.index [10] & ~_05134_;
	assign _05137_ = _07660_ | _04648_;
	assign _05138_ = _05137_ | _07758_;
	assign _05139_ = _05138_ | _01986_;
	assign _05140_ = _01875_ & ~_05139_;
	assign _05141_ = _02800_ | _02097_;
	assign _05142_ = _05141_ | \mchip.index [9];
	assign _05143_ = _05142_ | \mchip.index [10];
	assign _05144_ = _01875_ & ~_05143_;
	assign _05145_ = _01316_ | \mchip.index [5];
	assign _05146_ = _05145_ | \mchip.index [6];
	assign _05148_ = _05146_ | \mchip.index [7];
	assign _05149_ = _05148_ | _04648_;
	assign _05150_ = \mchip.index [9] & ~_05149_;
	assign _05151_ = _01179_ | _04648_;
	assign _05152_ = _05151_ | \mchip.index [9];
	assign _05153_ = _01875_ & ~_05152_;
	assign _05154_ = _01850_ | \mchip.index [8];
	assign _05155_ = _05154_ | \mchip.index [9];
	assign _05156_ = _05155_ | \mchip.index [10];
	assign _05157_ = _01875_ & ~_05156_;
	assign _05159_ = _02943_ | _07758_;
	assign _05160_ = _05159_ | _01986_;
	assign _05161_ = _01875_ & ~_05160_;
	assign _05162_ = _01823_ | _02984_;
	assign _05163_ = _05162_ | _01986_;
	assign _05164_ = \mchip.index [11] & ~_05163_;
	assign _05165_ = _00934_ | _02984_;
	assign _05166_ = _05165_ | \mchip.index [7];
	assign _05167_ = _05166_ | _04648_;
	assign _05168_ = _05167_ | \mchip.index [9];
	assign _05170_ = _05168_ | \mchip.index [10];
	assign _05171_ = \mchip.index [11] & ~_05170_;
	assign _05172_ = _06900_ | _02984_;
	assign _05173_ = _05172_ | _02097_;
	assign _05174_ = _05173_ | _04648_;
	assign _05175_ = _05174_ | _07758_;
	assign _05176_ = _01986_ & ~_05175_;
	assign _05177_ = _07848_ | _02984_;
	assign _05178_ = _05177_ | \mchip.index [8];
	assign _05179_ = _05178_ | _07758_;
	assign _05181_ = _05179_ | \mchip.index [10];
	assign _05182_ = _01875_ & ~_05181_;
	assign _05183_ = _04325_ | _02097_;
	assign _05184_ = _05183_ | \mchip.index [8];
	assign _05185_ = \mchip.index [11] & ~_05184_;
	assign _05186_ = _01099_ | \mchip.index [6];
	assign _05187_ = _05186_ | \mchip.index [7];
	assign _05188_ = _05187_ | _04648_;
	assign _05189_ = _05188_ | \mchip.index [9];
	assign _05190_ = _05189_ | _01986_;
	assign _05192_ = _01875_ & ~_05190_;
	assign _05193_ = _01869_ | \mchip.index [7];
	assign _05194_ = _05193_ | _01986_;
	assign _05195_ = \mchip.index [11] & ~_05194_;
	assign _05196_ = _01904_ | _02097_;
	assign _05197_ = _05196_ | _04648_;
	assign _05198_ = _01986_ & ~_05197_;
	assign _05199_ = _01184_ | \mchip.index [10];
	assign _05200_ = \mchip.index [11] & ~_05199_;
	assign _05201_ = _00713_ | \mchip.index [7];
	assign _05204_ = _05201_ | \mchip.index [8];
	assign _05205_ = _05204_ | \mchip.index [9];
	assign _05206_ = \mchip.index [11] & ~_05205_;
	assign _05207_ = _00600_ | \mchip.index [6];
	assign _05208_ = _05207_ | _02097_;
	assign _05209_ = _05208_ | _01986_;
	assign _05210_ = \mchip.index [11] & ~_05209_;
	assign _05211_ = _02998_ | _07758_;
	assign _05212_ = \mchip.index [10] & ~_05211_;
	assign _05213_ = _00476_ | _02097_;
	assign _05215_ = _05213_ | _04648_;
	assign _05216_ = _05215_ | \mchip.index [9];
	assign _05217_ = \mchip.index [10] & ~_05216_;
	assign _05218_ = _01431_ | \mchip.index [5];
	assign _05219_ = _05218_ | \mchip.index [6];
	assign _05220_ = _05219_ | _01986_;
	assign _05221_ = \mchip.index [11] & ~_05220_;
	assign _05222_ = _04193_ | \mchip.index [6];
	assign _05223_ = _05222_ | \mchip.index [7];
	assign _05224_ = _05223_ | \mchip.index [8];
	assign _05226_ = _05224_ | _07758_;
	assign _05227_ = _05226_ | \mchip.index [10];
	assign _05228_ = \mchip.index [11] & ~_05227_;
	assign _05229_ = _03278_ | _02097_;
	assign _05230_ = _05229_ | _01986_;
	assign _05231_ = \mchip.index [11] & ~_05230_;
	assign _05232_ = _01417_ | \mchip.index [6];
	assign _05233_ = _05232_ | _02097_;
	assign _05234_ = _05233_ | \mchip.index [8];
	assign _05235_ = _07758_ & ~_05234_;
	assign _05237_ = _01178_ | \mchip.index [7];
	assign _05238_ = _05237_ | \mchip.index [8];
	assign _05239_ = _05238_ | \mchip.index [9];
	assign _05240_ = _01875_ & ~_05239_;
	assign _05241_ = _00261_ | _02984_;
	assign _05242_ = _05241_ | _02097_;
	assign _05243_ = _05242_ | _04648_;
	assign _05244_ = _05243_ | _07758_;
	assign _05245_ = _01875_ & ~_05244_;
	assign _05246_ = _01490_ | _01098_;
	assign _05248_ = _05246_ | \mchip.index [5];
	assign _05249_ = _05248_ | \mchip.index [6];
	assign _05250_ = _05249_ | \mchip.index [7];
	assign _05251_ = _05250_ | _01986_;
	assign _05252_ = \mchip.index [11] & ~_05251_;
	assign _05253_ = _02540_ | \mchip.index [6];
	assign _05254_ = _05253_ | \mchip.index [7];
	assign _05255_ = _05254_ | \mchip.index [9];
	assign _05256_ = _05255_ | \mchip.index [10];
	assign _05257_ = _01875_ & ~_05256_;
	assign _05259_ = _00417_ | \mchip.index [8];
	assign _05260_ = _05259_ | \mchip.index [9];
	assign _05261_ = \mchip.index [10] & ~_05260_;
	assign _05262_ = _01380_ | \mchip.index [8];
	assign _05263_ = \mchip.index [11] & ~_05262_;
	assign _05264_ = _02895_ | _02984_;
	assign _05265_ = _05264_ | _04648_;
	assign _05266_ = _05265_ | _07758_;
	assign _05267_ = _01875_ & ~_05266_;
	assign _05268_ = _03984_ | \mchip.index [8];
	assign _05270_ = _05268_ | \mchip.index [9];
	assign _05271_ = \mchip.index [11] & ~_05270_;
	assign _05272_ = _06378_ | _05424_;
	assign _05273_ = _05272_ | _02984_;
	assign _05274_ = _05273_ | \mchip.index [9];
	assign _05275_ = \mchip.index [10] & ~_05274_;
	assign _05276_ = _00507_ | \mchip.index [6];
	assign _05277_ = _05276_ | \mchip.index [7];
	assign _05278_ = _05277_ | _01986_;
	assign _05279_ = \mchip.index [11] & ~_05278_;
	assign _05281_ = _03454_ | \mchip.index [6];
	assign _05282_ = _05281_ | _07758_;
	assign _05283_ = _01875_ & ~_05282_;
	assign _05284_ = _01750_ | _04648_;
	assign _05285_ = \mchip.index [10] & ~_05284_;
	assign _05286_ = _01342_ | _02097_;
	assign _05287_ = _05286_ | _04648_;
	assign _05288_ = _05287_ | _07758_;
	assign _05289_ = \mchip.index [10] & ~_05288_;
	assign _05290_ = _04633_ | _07758_;
	assign _05292_ = _01986_ & ~_05290_;
	assign _05293_ = _01576_ | \mchip.index [7];
	assign _05294_ = _05293_ | _04648_;
	assign _05295_ = _05294_ | _07758_;
	assign _05296_ = _05295_ | _01986_;
	assign _05297_ = _01875_ & ~_05296_;
	assign _05298_ = _01599_ | \mchip.index [7];
	assign _05299_ = _05298_ | _04648_;
	assign _05300_ = _05299_ | \mchip.index [9];
	assign _05301_ = _05300_ | \mchip.index [10];
	assign _05303_ = _01875_ & ~_05301_;
	assign _05304_ = _05680_ | _05424_;
	assign _05305_ = _05304_ | \mchip.index [7];
	assign _05306_ = _05305_ | \mchip.index [9];
	assign _05307_ = \mchip.index [10] & ~_05306_;
	assign _05308_ = _07733_ | \mchip.index [8];
	assign _05309_ = _05308_ | _07758_;
	assign _05310_ = _05309_ | \mchip.index [10];
	assign _05311_ = _01875_ & ~_05310_;
	assign _05312_ = _00261_ | \mchip.index [8];
	assign _05315_ = _05312_ | _07758_;
	assign _05316_ = _05315_ | \mchip.index [10];
	assign _05317_ = _01875_ & ~_05316_;
	assign _05318_ = _07355_ | _02097_;
	assign _05319_ = _05318_ | \mchip.index [8];
	assign _05320_ = _05319_ | _07758_;
	assign _05321_ = _05320_ | \mchip.index [10];
	assign _05322_ = _01875_ & ~_05321_;
	assign _05323_ = _00705_ | _02984_;
	assign _05324_ = _05323_ | \mchip.index [7];
	assign _05326_ = _05324_ | \mchip.index [9];
	assign _05327_ = \mchip.index [11] & ~_05326_;
	assign _05328_ = _05323_ | \mchip.index [8];
	assign _05329_ = _05328_ | _07758_;
	assign _05330_ = \mchip.index [10] & ~_05329_;
	assign _05331_ = _00687_ | _04648_;
	assign _05332_ = _05331_ | \mchip.index [10];
	assign _05333_ = \mchip.index [11] & ~_05332_;
	assign _05334_ = _05165_ | _02097_;
	assign _05335_ = _05334_ | \mchip.index [8];
	assign _05337_ = _05335_ | _07758_;
	assign _05338_ = _01986_ & ~_05337_;
	assign _05339_ = _01440_ | \mchip.index [9];
	assign _05340_ = \mchip.index [11] & ~_05339_;
	assign _05341_ = _01975_ | _02984_;
	assign _05342_ = _05341_ | _02097_;
	assign _05343_ = _05342_ | _04648_;
	assign _05344_ = _05343_ | _07758_;
	assign _05345_ = _05344_ | _01986_;
	assign _05346_ = \mchip.index [11] & ~_05345_;
	assign _05348_ = _07640_ | \mchip.index [7];
	assign _05349_ = _01875_ & ~_05348_;
	assign _05350_ = _01317_ | _02097_;
	assign _05351_ = _05350_ | \mchip.index [9];
	assign _05352_ = \mchip.index [11] & ~_05351_;
	assign _05353_ = _07783_ | _02097_;
	assign _05354_ = _05353_ | \mchip.index [8];
	assign _05355_ = _05354_ | \mchip.index [9];
	assign _05356_ = _01986_ & ~_05355_;
	assign _05357_ = _06445_ | _02984_;
	assign _05359_ = _05357_ | \mchip.index [7];
	assign _05360_ = _05359_ | \mchip.index [8];
	assign _05361_ = _05360_ | _07758_;
	assign _05362_ = _05361_ | \mchip.index [10];
	assign _05363_ = \mchip.index [11] & ~_05362_;
	assign _05364_ = _02850_ | \mchip.index [6];
	assign _05365_ = _05364_ | \mchip.index [7];
	assign _05366_ = _05365_ | _07758_;
	assign _05367_ = \mchip.index [11] & ~_05366_;
	assign _05368_ = _01113_ | _04648_;
	assign _05370_ = _05368_ | _07758_;
	assign _05371_ = _05370_ | _01986_;
	assign _05372_ = \mchip.index [11] & ~_05371_;
	assign _05373_ = _01839_ | _02097_;
	assign _05374_ = _05373_ | _04648_;
	assign _05375_ = _05374_ | \mchip.index [10];
	assign _05376_ = _01875_ & ~_05375_;
	assign _05377_ = _02948_ | \mchip.index [8];
	assign _05378_ = \mchip.index [10] & ~_05377_;
	assign _05379_ = _01799_ | _04648_;
	assign _05381_ = _05379_ | \mchip.index [9];
	assign _05382_ = \mchip.index [10] & ~_05381_;
	assign _05383_ = _03269_ | \mchip.index [7];
	assign _05384_ = _05383_ | _04648_;
	assign _05385_ = _05384_ | \mchip.index [9];
	assign _05386_ = _01875_ & ~_05385_;
	assign _05387_ = _02601_ | \mchip.index [7];
	assign _05388_ = _05387_ | _04648_;
	assign _05389_ = \mchip.index [11] & ~_05388_;
	assign _05390_ = _01311_ | \mchip.index [7];
	assign _05392_ = _05390_ | _04648_;
	assign _05393_ = _05392_ | \mchip.index [10];
	assign _05394_ = \mchip.index [11] & ~_05393_;
	assign _05395_ = _01389_ | \mchip.index [6];
	assign _05396_ = _05395_ | \mchip.index [7];
	assign _05397_ = \mchip.index [11] & ~_05396_;
	assign _05398_ = _01399_ | \mchip.index [9];
	assign _05399_ = _01986_ & ~_05398_;
	assign _05400_ = _01776_ | _02984_;
	assign _05401_ = _05400_ | \mchip.index [7];
	assign _05403_ = _05401_ | _04648_;
	assign _05404_ = _05403_ | \mchip.index [9];
	assign _05405_ = \mchip.index [10] & ~_05404_;
	assign _05406_ = _02039_ | \mchip.index [7];
	assign _05407_ = _05406_ | _07758_;
	assign _05408_ = _05407_ | _01986_;
	assign _05409_ = _01875_ & ~_05408_;
	assign _05410_ = _02100_ | \mchip.index [8];
	assign _05411_ = _05410_ | _07758_;
	assign _05412_ = _01875_ & ~_05411_;
	assign _05414_ = _07709_ | _02097_;
	assign _05415_ = _05414_ | _04648_;
	assign _05416_ = _05415_ | _07758_;
	assign _05417_ = _01986_ & ~_05416_;
	assign _05418_ = _01791_ | \mchip.index [7];
	assign _05419_ = _05418_ | _07758_;
	assign _05420_ = _05419_ | \mchip.index [10];
	assign _05421_ = \mchip.index [11] & ~_05420_;
	assign _05422_ = _07637_ | _05424_;
	assign _05423_ = _05422_ | \mchip.index [7];
	assign _05426_ = _05423_ | \mchip.index [8];
	assign _05427_ = _05426_ | _07758_;
	assign _05428_ = \mchip.index [10] & ~_05427_;
	assign _05429_ = _03154_ | \mchip.index [7];
	assign _05430_ = _05429_ | _04648_;
	assign _05431_ = _05430_ | \mchip.index [9];
	assign _05432_ = \mchip.index [10] & ~_05431_;
	assign _05433_ = _02408_ | _05424_;
	assign _05434_ = _05433_ | _02984_;
	assign _05435_ = _05434_ | _02097_;
	assign _05437_ = _05435_ | _04648_;
	assign _05438_ = \mchip.index [10] & ~_05437_;
	assign _05439_ = _00561_ | \mchip.index [8];
	assign _05440_ = _05439_ | _07758_;
	assign _05441_ = \mchip.index [10] & ~_05440_;
	assign _05442_ = _01971_ | \mchip.index [7];
	assign _05443_ = _05442_ | _07758_;
	assign _05444_ = \mchip.index [11] & ~_05443_;
	assign _05445_ = _07714_ | _05424_;
	assign _05446_ = _05445_ | _02984_;
	assign _05448_ = _05446_ | _07758_;
	assign _05449_ = \mchip.index [11] & ~_05448_;
	assign _05450_ = _00516_ | _02097_;
	assign _05451_ = _05450_ | \mchip.index [8];
	assign _05452_ = _05451_ | \mchip.index [9];
	assign _05453_ = _05452_ | \mchip.index [10];
	assign _05454_ = _01875_ & ~_05453_;
	assign _05455_ = _01749_ | _02097_;
	assign _05456_ = _05455_ | _04648_;
	assign _05457_ = \mchip.index [11] & ~_05456_;
	assign _05459_ = _03821_ | \mchip.index [8];
	assign _05460_ = _05459_ | \mchip.index [10];
	assign _05461_ = _01875_ & ~_05460_;
	assign _05462_ = _01230_ | _05424_;
	assign _05463_ = \mchip.index [7] & ~_05462_;
	assign _05464_ = _00110_ | _02097_;
	assign _05465_ = _05464_ | \mchip.index [8];
	assign _05466_ = _05465_ | \mchip.index [9];
	assign _05467_ = _05466_ | \mchip.index [10];
	assign _05468_ = _01875_ & ~_05467_;
	assign _05470_ = _03817_ | _07758_;
	assign _05471_ = _05470_ | _01986_;
	assign _05472_ = _01875_ & ~_05471_;
	assign _05473_ = _00484_ | _02984_;
	assign _05474_ = _05473_ | _02097_;
	assign _05475_ = _05474_ | \mchip.index [8];
	assign _05476_ = _05475_ | \mchip.index [9];
	assign _05477_ = \mchip.index [10] & ~_05476_;
	assign _05478_ = _00838_ | _02097_;
	assign _05479_ = _05478_ | \mchip.index [9];
	assign _05481_ = _01875_ & ~_05479_;
	assign _05482_ = _02076_ | _04648_;
	assign _05483_ = \mchip.index [10] & ~_05482_;
	assign _05484_ = _01110_ | \mchip.index [7];
	assign _05485_ = _05484_ | _04648_;
	assign _05486_ = _05485_ | _01986_;
	assign _05487_ = _01875_ & ~_05486_;
	assign _05488_ = ~(_01765_ & \mchip.index [9]);
	assign _05489_ = \mchip.index [10] & ~_05488_;
	assign _05490_ = _01191_ | \mchip.index [8];
	assign _05492_ = _05490_ | \mchip.index [10];
	assign _05493_ = _01875_ & ~_05492_;
	assign _05494_ = _01944_ | _07758_;
	assign _05495_ = \mchip.index [11] & ~_05494_;
	assign _05496_ = _01376_ | _02984_;
	assign _05497_ = _05496_ | _04648_;
	assign _05498_ = _05497_ | _07758_;
	assign _05499_ = _01986_ & ~_05498_;
	assign _05500_ = _04157_ | \mchip.index [9];
	assign _05501_ = \mchip.index [11] & ~_05500_;
	assign _05503_ = _02707_ | \mchip.index [8];
	assign _05504_ = _05503_ | _07758_;
	assign _05505_ = _05504_ | \mchip.index [10];
	assign _05506_ = _01875_ & ~_05505_;
	assign _05507_ = _01840_ | \mchip.index [9];
	assign _05508_ = _01875_ & ~_05507_;
	assign _05509_ = _02884_ | _04648_;
	assign _05510_ = _05509_ | _07758_;
	assign _05511_ = _01986_ & ~_05510_;
	assign _05512_ = _04071_ | \mchip.index [7];
	assign _05514_ = _05512_ | _01986_;
	assign _05515_ = \mchip.index [11] & ~_05514_;
	assign _05516_ = _04237_ | \mchip.index [8];
	assign _05517_ = _05516_ | _07758_;
	assign _05518_ = _05517_ | \mchip.index [10];
	assign _05519_ = _01875_ & ~_05518_;
	assign _05520_ = _00380_ | _02984_;
	assign _05521_ = _05520_ | _07758_;
	assign _05522_ = _05521_ | \mchip.index [10];
	assign _05523_ = \mchip.index [11] & ~_05522_;
	assign _05525_ = _01343_ | _02097_;
	assign _05526_ = _05525_ | _04648_;
	assign _05527_ = _05526_ | \mchip.index [9];
	assign _05528_ = \mchip.index [10] & ~_05527_;
	assign _05529_ = _02952_ | _04648_;
	assign _05530_ = _05529_ | _07758_;
	assign _05531_ = _01986_ & ~_05530_;
	assign _05532_ = _02069_ | _07758_;
	assign _05533_ = _05532_ | _01986_;
	assign _05534_ = _01875_ & ~_05533_;
	assign _05537_ = _03154_ | _02097_;
	assign _05538_ = _05537_ | \mchip.index [8];
	assign _05539_ = _05538_ | _07758_;
	assign _05540_ = \mchip.index [10] & ~_05539_;
	assign _05541_ = _02728_ | _02097_;
	assign _05542_ = _05541_ | \mchip.index [8];
	assign _05543_ = _05542_ | \mchip.index [9];
	assign _05544_ = \mchip.index [10] & ~_05543_;
	assign _05545_ = _00154_ | _02984_;
	assign _05546_ = _05545_ | \mchip.index [7];
	assign _05548_ = _05546_ | \mchip.index [8];
	assign _05549_ = _05548_ | \mchip.index [9];
	assign _05550_ = \mchip.index [10] & ~_05549_;
	assign _05551_ = _04294_ | \mchip.index [10];
	assign _05552_ = \mchip.index [11] & ~_05551_;
	assign _05553_ = _07758_ & ~_02958_;
	assign _05554_ = _06911_ | \mchip.index [7];
	assign _05555_ = _05554_ | \mchip.index [8];
	assign _05556_ = _05555_ | \mchip.index [9];
	assign _05557_ = \mchip.index [11] & ~_05556_;
	assign _05559_ = _01106_ | _01986_;
	assign _05560_ = _01875_ & ~_05559_;
	assign _05561_ = _07741_ | _02097_;
	assign _05562_ = _05561_ | _07758_;
	assign _05563_ = \mchip.index [11] & ~_05562_;
	assign _05564_ = _02505_ | _02097_;
	assign _05565_ = _05564_ | _01986_;
	assign _05566_ = \mchip.index [11] & ~_05565_;
	assign _05567_ = _04081_ | _02097_;
	assign _05568_ = _01986_ & ~_05567_;
	assign _05570_ = _03155_ | _02097_;
	assign _05571_ = _05570_ | \mchip.index [9];
	assign _05572_ = _05571_ | \mchip.index [10];
	assign _05573_ = _01875_ & ~_05572_;
	assign _05574_ = _00816_ | _02984_;
	assign _05575_ = _05574_ | _02097_;
	assign _05576_ = _05575_ | _04648_;
	assign _05577_ = _05576_ | \mchip.index [9];
	assign _05578_ = \mchip.index [10] & ~_05577_;
	assign _05579_ = _04222_ | _02097_;
	assign _05581_ = _05579_ | _04648_;
	assign _05582_ = _05581_ | _07758_;
	assign _05583_ = _01986_ & ~_05582_;
	assign _05584_ = _01300_ | _04648_;
	assign _05585_ = _05584_ | _01986_;
	assign _05586_ = _01875_ & ~_05585_;
	assign _05587_ = _02123_ | _07758_;
	assign _05588_ = _05587_ | \mchip.index [10];
	assign _05589_ = _01875_ & ~_05588_;
	assign _05590_ = _07701_ | _02984_;
	assign _05592_ = _05590_ | \mchip.index [7];
	assign _05593_ = _05592_ | _04648_;
	assign _05594_ = _05593_ | _07758_;
	assign _05595_ = _05594_ | \mchip.index [10];
	assign _05596_ = _01875_ & ~_05595_;
	assign _05597_ = _01325_ | \mchip.index [6];
	assign _05598_ = _05597_ | \mchip.index [7];
	assign _05599_ = _05598_ | _04648_;
	assign _05600_ = _05599_ | \mchip.index [9];
	assign _05601_ = _05600_ | \mchip.index [10];
	assign _05603_ = \mchip.index [11] & ~_05601_;
	assign _05604_ = _01379_ | _07758_;
	assign _05605_ = _01986_ & ~_05604_;
	assign _05606_ = _00324_ | \mchip.index [6];
	assign _05607_ = _05606_ | _02097_;
	assign _05608_ = _05607_ | _04648_;
	assign _05609_ = _05608_ | \mchip.index [10];
	assign _05610_ = _01875_ & ~_05609_;
	assign _05611_ = _01304_ | \mchip.index [7];
	assign _05612_ = _05611_ | _01986_;
	assign _05614_ = \mchip.index [11] & ~_05612_;
	assign _05615_ = _02116_ | \mchip.index [9];
	assign _05616_ = _05615_ | \mchip.index [10];
	assign _05617_ = \mchip.index [11] & ~_05616_;
	assign _05618_ = _02696_ | _05424_;
	assign _05619_ = _05618_ | _02984_;
	assign _05620_ = _05619_ | \mchip.index [7];
	assign _05621_ = \mchip.index [11] & ~_05620_;
	assign _05622_ = _00531_ | \mchip.index [7];
	assign _05623_ = _05622_ | \mchip.index [8];
	assign _05625_ = _05623_ | \mchip.index [9];
	assign _05626_ = \mchip.index [11] & ~_05625_;
	assign _05627_ = _00836_ | _02984_;
	assign _05628_ = _05627_ | \mchip.index [7];
	assign _05629_ = _05628_ | \mchip.index [8];
	assign _05630_ = _05629_ | _07758_;
	assign _05631_ = \mchip.index [10] & ~_05630_;
	assign _05632_ = _00461_ | _05424_;
	assign _05633_ = _05632_ | \mchip.index [6];
	assign _05634_ = _05633_ | \mchip.index [7];
	assign _05636_ = _05634_ | _01986_;
	assign _05637_ = \mchip.index [11] & ~_05636_;
	assign _05638_ = _05383_ | _07758_;
	assign _05639_ = \mchip.index [11] & ~_05638_;
	assign _05640_ = _05554_ | _04648_;
	assign _05641_ = _05640_ | _07758_;
	assign _05642_ = _01986_ & ~_05641_;
	assign _05643_ = _00402_ | _04648_;
	assign _05644_ = _05643_ | \mchip.index [9];
	assign _05645_ = _05644_ | \mchip.index [10];
	assign _05648_ = _01875_ & ~_05645_;
	assign _05649_ = _02007_ | \mchip.index [8];
	assign _05650_ = _05649_ | \mchip.index [9];
	assign _05651_ = \mchip.index [11] & ~_05650_;
	assign _05652_ = _05564_ | _04648_;
	assign _05653_ = _05652_ | \mchip.index [9];
	assign _05654_ = \mchip.index [10] & ~_05653_;
	assign _05655_ = _01629_ | \mchip.index [8];
	assign _05656_ = _05655_ | \mchip.index [9];
	assign _05657_ = _01986_ & ~_05656_;
	assign _05659_ = _05254_ | _01986_;
	assign _05660_ = \mchip.index [11] & ~_05659_;
	assign _05661_ = _02517_ & ~\mchip.index [7];
	assign _05662_ = _03954_ | \mchip.index [6];
	assign _05663_ = _05662_ | \mchip.index [8];
	assign _05664_ = _05663_ | \mchip.index [9];
	assign _05665_ = \mchip.index [10] & ~_05664_;
	assign _05666_ = _01552_ | _07758_;
	assign _05667_ = \mchip.index [11] & ~_05666_;
	assign _05668_ = _03040_ | \mchip.index [8];
	assign _05670_ = _05668_ | \mchip.index [9];
	assign _05671_ = \mchip.index [10] & ~_05670_;
	assign _05672_ = \mchip.index [10] & ~_03025_;
	assign _05673_ = _03884_ & ~_01986_;
	assign _05674_ = _01607_ | \mchip.index [8];
	assign _05675_ = \mchip.index [11] & ~_05674_;
	assign _05676_ = _06545_ | _02984_;
	assign _05677_ = _05676_ | _02097_;
	assign _05678_ = _05677_ | \mchip.index [9];
	assign _05679_ = _05678_ | \mchip.index [10];
	assign _05681_ = _01875_ & ~_05679_;
	assign _05682_ = _04639_ | _02097_;
	assign _05683_ = _05682_ | _04648_;
	assign _05684_ = _05683_ | \mchip.index [9];
	assign _05685_ = \mchip.index [10] & ~_05684_;
	assign _05686_ = _03825_ | \mchip.index [8];
	assign _05687_ = _05686_ | \mchip.index [9];
	assign _05688_ = \mchip.index [10] & ~_05687_;
	assign _05689_ = _01341_ | \mchip.index [7];
	assign _05690_ = _05689_ | _04648_;
	assign _05692_ = _05690_ | \mchip.index [9];
	assign _05693_ = _05692_ | \mchip.index [10];
	assign _05694_ = _01875_ & ~_05693_;
	assign _05695_ = _04601_ | _02097_;
	assign _05696_ = _05695_ | _04648_;
	assign _05697_ = _05696_ | _07758_;
	assign _05698_ = _01986_ & ~_05697_;
	assign _05699_ = _01818_ | \mchip.index [9];
	assign _05700_ = _05699_ | \mchip.index [10];
	assign _05701_ = _01875_ & ~_05700_;
	assign _05703_ = _02100_ | \mchip.index [7];
	assign _05704_ = _05703_ | _04648_;
	assign _05705_ = _05704_ | \mchip.index [9];
	assign _05706_ = \mchip.index [11] & ~_05705_;
	assign _05707_ = _02458_ | \mchip.index [8];
	assign _05708_ = _05707_ | _07758_;
	assign _05709_ = \mchip.index [10] & ~_05708_;
	assign _05710_ = _01159_ | _01986_;
	assign _05711_ = \mchip.index [11] & ~_05710_;
	assign _05712_ = _01297_ | _02097_;
	assign _05714_ = _05712_ | _01986_;
	assign _05715_ = \mchip.index [11] & ~_05714_;
	assign _05716_ = _04576_ | \mchip.index [6];
	assign _05717_ = _05716_ | \mchip.index [7];
	assign _05718_ = _05717_ | _07758_;
	assign _05719_ = _05718_ | _01986_;
	assign _05720_ = _01875_ & ~_05719_;
	assign _05721_ = _01384_ | _04648_;
	assign _05722_ = _05721_ | _07758_;
	assign _05723_ = _05722_ | _01986_;
	assign _05725_ = _01875_ & ~_05723_;
	assign _05726_ = _01097_ | \mchip.index [7];
	assign _05727_ = _05726_ | _04648_;
	assign _05728_ = _05727_ | _07758_;
	assign _05729_ = _01986_ & ~_05728_;
	assign _05730_ = _03773_ | _04648_;
	assign _05731_ = _05730_ | _07758_;
	assign _05732_ = _05731_ | _01986_;
	assign _05733_ = _01875_ & ~_05732_;
	assign _05734_ = _01635_ | _07758_;
	assign _05736_ = _01986_ & ~_05734_;
	assign _05737_ = _02713_ | \mchip.index [7];
	assign _05738_ = _05737_ | _07758_;
	assign _05739_ = _05738_ | \mchip.index [10];
	assign _05740_ = \mchip.index [11] & ~_05739_;
	assign _05741_ = _07671_ | _05424_;
	assign _05742_ = _05741_ | \mchip.index [6];
	assign _05743_ = _02097_ & ~_05742_;
	assign _05744_ = _07675_ | _02984_;
	assign _05745_ = _05744_ | \mchip.index [7];
	assign _05747_ = _05745_ | _04648_;
	assign _05748_ = _05747_ | \mchip.index [9];
	assign _05749_ = \mchip.index [10] & ~_05748_;
	assign _05750_ = _04432_ & ~_01875_;
	assign _05751_ = \mchip.index [11] & ~_03367_;
	assign _05752_ = _04626_ | \mchip.index [6];
	assign _05753_ = _05752_ | \mchip.index [8];
	assign _05754_ = _05753_ | \mchip.index [9];
	assign _05755_ = \mchip.index [11] & ~_05754_;
	assign _05756_ = _07774_ | _04648_;
	assign _05759_ = _05756_ | \mchip.index [9];
	assign _05760_ = \mchip.index [10] & ~_05759_;
	assign _05761_ = \mchip.index [6] & ~_02780_;
	assign _05762_ = _01481_ | \mchip.index [7];
	assign _05763_ = _05762_ | \mchip.index [9];
	assign _05764_ = \mchip.index [10] & ~_05763_;
	assign _05765_ = _07676_ | _02097_;
	assign _05766_ = _05765_ | \mchip.index [9];
	assign _05767_ = \mchip.index [11] & ~_05766_;
	assign _05768_ = _04321_ | _04648_;
	assign _05770_ = _05768_ | \mchip.index [10];
	assign _05771_ = \mchip.index [11] & ~_05770_;
	assign _05772_ = _02022_ | \mchip.index [9];
	assign _05773_ = _05772_ | \mchip.index [10];
	assign _05774_ = _01875_ & ~_05773_;
	assign _05775_ = _00268_ | \mchip.index [7];
	assign _05776_ = _05775_ | \mchip.index [8];
	assign _05777_ = _05776_ | _07758_;
	assign _05778_ = \mchip.index [11] & ~_05777_;
	assign _05779_ = _02855_ | \mchip.index [5];
	assign _05781_ = _05779_ | _02984_;
	assign _05782_ = _05781_ | _02097_;
	assign _05783_ = _05782_ | \mchip.index [9];
	assign _05784_ = _05783_ | \mchip.index [10];
	assign _05785_ = _01875_ & ~_05784_;
	assign _05786_ = _06378_ | \mchip.index [6];
	assign _05787_ = _05786_ | \mchip.index [8];
	assign _05788_ = _05787_ | \mchip.index [9];
	assign _05789_ = _05788_ | \mchip.index [10];
	assign _05790_ = _01875_ & ~_05789_;
	assign _05792_ = _04482_ | _02984_;
	assign _05793_ = _05792_ | _02097_;
	assign _05794_ = _05793_ | _07758_;
	assign _05795_ = _05794_ | \mchip.index [10];
	assign _05796_ = \mchip.index [11] & ~_05795_;
	assign _05797_ = _01581_ | \mchip.index [7];
	assign _05798_ = _05797_ | \mchip.index [8];
	assign _05799_ = _05798_ | \mchip.index [9];
	assign _05800_ = \mchip.index [10] & ~_05799_;
	assign _05801_ = _01738_ | \mchip.index [7];
	assign _05803_ = _05801_ | _04648_;
	assign _05804_ = \mchip.index [11] & ~_05803_;
	assign _05805_ = _02192_ | \mchip.index [8];
	assign _05806_ = _05805_ | \mchip.index [10];
	assign _05807_ = _01875_ & ~_05806_;
	assign _05808_ = _00397_ | _02097_;
	assign _05809_ = _05808_ | _04648_;
	assign _05810_ = _05809_ | _07758_;
	assign _05811_ = _01986_ & ~_05810_;
	assign _05812_ = _02150_ | _04648_;
	assign _05814_ = _05812_ | _07758_;
	assign _05815_ = _01875_ & ~_05814_;
	assign _05816_ = _01899_ | \mchip.index [7];
	assign _05817_ = _05816_ | _07758_;
	assign _05818_ = _05817_ | \mchip.index [10];
	assign _05819_ = \mchip.index [11] & ~_05818_;
	assign _05820_ = _01607_ | _07758_;
	assign _05821_ = \mchip.index [11] & ~_05820_;
	assign _05822_ = _03839_ | \mchip.index [9];
	assign _05823_ = \mchip.index [10] & ~_05822_;
	assign _05825_ = _05478_ | _04648_;
	assign _05826_ = _01875_ & ~_05825_;
	assign _05827_ = _07828_ | \mchip.index [6];
	assign _05828_ = _05827_ | _02097_;
	assign _05829_ = _05828_ | _04648_;
	assign _05830_ = \mchip.index [11] & ~_05829_;
	assign _05831_ = _01588_ | _04648_;
	assign _05832_ = _01986_ & ~_05831_;
	assign _05833_ = _00431_ | \mchip.index [9];
	assign _05834_ = \mchip.index [10] & ~_05833_;
	assign _05836_ = _04449_ | _07758_;
	assign _05837_ = \mchip.index [11] & ~_05836_;
	assign _05838_ = _01387_ | _02984_;
	assign _05839_ = _05838_ | _02097_;
	assign _05840_ = _05839_ | \mchip.index [9];
	assign _05841_ = \mchip.index [11] & ~_05840_;
	assign _05842_ = _02127_ | \mchip.index [8];
	assign _05843_ = _05842_ | \mchip.index [9];
	assign _05844_ = \mchip.index [11] & ~_05843_;
	assign _05845_ = _04334_ | _02097_;
	assign _05847_ = \mchip.index [11] & ~_05845_;
	assign _05848_ = _01914_ | _02097_;
	assign _05849_ = _05848_ | \mchip.index [8];
	assign _05850_ = \mchip.index [10] & ~_05849_;
	assign _05851_ = _03342_ | _07758_;
	assign _05852_ = _01986_ & ~_05851_;
	assign _05853_ = _06545_ | _02097_;
	assign _05854_ = _05853_ | \mchip.index [8];
	assign _05855_ = _05854_ | _07758_;
	assign _05856_ = \mchip.index [11] & ~_05855_;
	assign _05858_ = _07831_ | \mchip.index [8];
	assign _05859_ = \mchip.index [10] & ~_05858_;
	assign _05860_ = _02209_ | _05424_;
	assign _05861_ = \mchip.index [7] & ~_05860_;
	assign _05862_ = _01191_ | \mchip.index [7];
	assign _05863_ = _05862_ | _04648_;
	assign _05864_ = \mchip.index [10] & ~_05863_;
	assign _05865_ = _01237_ | \mchip.index [8];
	assign _05866_ = _05865_ | \mchip.index [10];
	assign _05867_ = _01875_ & ~_05866_;
	assign _05870_ = _02167_ | _02097_;
	assign _05871_ = _05870_ | \mchip.index [10];
	assign _05872_ = _01875_ & ~_05871_;
	assign _05873_ = _02672_ | \mchip.index [7];
	assign _05874_ = _05873_ | \mchip.index [8];
	assign _05875_ = _05874_ | _07758_;
	assign _05876_ = \mchip.index [10] & ~_05875_;
	assign _05877_ = _03360_ | \mchip.index [8];
	assign _05878_ = _05877_ | \mchip.index [9];
	assign _05879_ = \mchip.index [10] & ~_05878_;
	assign _05881_ = _01277_ | _04648_;
	assign _05882_ = _05881_ | \mchip.index [9];
	assign _05883_ = \mchip.index [11] & ~_05882_;
	assign _05884_ = _03091_ | \mchip.index [7];
	assign _05885_ = _05884_ | \mchip.index [9];
	assign _05886_ = \mchip.index [10] & ~_05885_;
	assign _05887_ = _03084_ | _02984_;
	assign _05888_ = _05887_ | _02097_;
	assign _05889_ = _05888_ | _04648_;
	assign _05890_ = _05889_ | \mchip.index [9];
	assign _05892_ = \mchip.index [11] & ~_05890_;
	assign _05893_ = _06445_ | \mchip.index [6];
	assign _05894_ = _05893_ | _02097_;
	assign _05895_ = _05894_ | _04648_;
	assign _05896_ = _05895_ | \mchip.index [9];
	assign _05897_ = _05896_ | _01986_;
	assign _05898_ = _01875_ & ~_05897_;
	assign _05899_ = _01651_ | _07758_;
	assign _05900_ = _01875_ & ~_05899_;
	assign _05901_ = _04484_ | \mchip.index [8];
	assign _05903_ = _05901_ | \mchip.index [9];
	assign _05904_ = \mchip.index [10] & ~_05903_;
	assign _05905_ = _05418_ | \mchip.index [8];
	assign _05906_ = _05905_ | \mchip.index [9];
	assign _05907_ = \mchip.index [10] & ~_05906_;
	assign _05908_ = _01986_ & ~_03088_;
	assign _05909_ = _05590_ | \mchip.index [8];
	assign _05910_ = _05909_ | \mchip.index [9];
	assign _05911_ = _05910_ | \mchip.index [10];
	assign _05912_ = _01875_ & ~_05911_;
	assign _05914_ = _04757_ | _04648_;
	assign _05915_ = \mchip.index [11] & ~_05914_;
	assign _05916_ = _04249_ | _05424_;
	assign _05917_ = _05916_ | _02097_;
	assign _05918_ = _05917_ | _01986_;
	assign _05919_ = \mchip.index [11] & ~_05918_;
	assign _05920_ = _01256_ | _01986_;
	assign _05921_ = _01875_ & ~_05920_;
	assign _05922_ = _01508_ | \mchip.index [7];
	assign _05923_ = _05922_ | \mchip.index [8];
	assign _05925_ = _05923_ | _07758_;
	assign _05926_ = \mchip.index [10] & ~_05925_;
	assign _05927_ = _01349_ | _01986_;
	assign _05928_ = \mchip.index [11] & ~_05927_;
	assign _05929_ = _01924_ | \mchip.index [8];
	assign _05930_ = _05929_ | _07758_;
	assign _05931_ = \mchip.index [10] & ~_05930_;
	assign _05932_ = _03389_ | _07758_;
	assign _05933_ = \mchip.index [11] & ~_05932_;
	assign _05934_ = _06578_ | \mchip.index [6];
	assign _05936_ = _05934_ | \mchip.index [8];
	assign _05937_ = _05936_ | _07758_;
	assign _05938_ = \mchip.index [10] & ~_05937_;
	assign _05939_ = _03236_ | _01986_;
	assign _05940_ = _01875_ & ~_05939_;
	assign _05941_ = _03239_ | _07758_;
	assign _05942_ = _01986_ & ~_05941_;
	assign _05943_ = _04508_ | \mchip.index [7];
	assign _05944_ = _05943_ | \mchip.index [8];
	assign _05945_ = _05944_ | \mchip.index [9];
	assign _05947_ = \mchip.index [11] & ~_05945_;
	assign _05948_ = _03381_ | \mchip.index [8];
	assign _05949_ = _05948_ | _07758_;
	assign _05950_ = \mchip.index [10] & ~_05949_;
	assign _05951_ = _05891_ | \mchip.index [10];
	assign _05952_ = \mchip.index [11] & ~_05951_;
	assign _05953_ = _01875_ & ~_02036_;
	assign _05954_ = _02770_ | \mchip.index [9];
	assign _05955_ = \mchip.index [11] & ~_05954_;
	assign _05956_ = _03444_ | \mchip.index [9];
	assign _05958_ = \mchip.index [10] & ~_05956_;
	assign _05959_ = _01842_ | \mchip.index [6];
	assign _05960_ = _05959_ | \mchip.index [7];
	assign _05961_ = _05960_ | \mchip.index [8];
	assign _05962_ = _05961_ | _07758_;
	assign _05963_ = \mchip.index [10] & ~_05962_;
	assign _05964_ = _02758_ | _02097_;
	assign _05965_ = _05964_ | \mchip.index [8];
	assign _05966_ = _05965_ | _07758_;
	assign _05967_ = _01986_ & ~_05966_;
	assign _05969_ = _03449_ | _02097_;
	assign _05970_ = _05969_ | _04648_;
	assign _05971_ = _01986_ & ~_05970_;
	assign _05972_ = _01783_ | _04648_;
	assign _05973_ = _05972_ | \mchip.index [9];
	assign _05974_ = _01986_ & ~_05973_;
	assign _05975_ = \mchip.index [9] & ~_02154_;
	assign _05976_ = _01316_ | _02097_;
	assign _05977_ = _05976_ | _04648_;
	assign _05978_ = _05977_ | \mchip.index [10];
	assign _05981_ = \mchip.index [11] & ~_05978_;
	assign _05982_ = _04484_ | _02097_;
	assign _05983_ = _05982_ | \mchip.index [8];
	assign _05984_ = \mchip.index [10] & ~_05983_;
	assign _05985_ = _01440_ | _07758_;
	assign _05986_ = \mchip.index [10] & ~_05985_;
	assign _05987_ = _03212_ | \mchip.index [8];
	assign _05988_ = _05987_ | \mchip.index [10];
	assign _05989_ = _01875_ & ~_05988_;
	assign _05990_ = _00631_ | \mchip.index [7];
	assign _05992_ = _05990_ | \mchip.index [8];
	assign _05993_ = \mchip.index [9] & ~_05992_;
	assign _05994_ = _02581_ | _04648_;
	assign _05995_ = _05994_ | _07758_;
	assign _05996_ = _05995_ | _01986_;
	assign _05997_ = \mchip.index [11] & ~_05996_;
	assign _05998_ = _05113_ | \mchip.index [6];
	assign _05999_ = _05998_ | \mchip.index [7];
	assign _06000_ = _05999_ | \mchip.index [8];
	assign _06001_ = _06000_ | \mchip.index [9];
	assign _06003_ = \mchip.index [11] & ~_06001_;
	assign _06004_ = _00836_ | _05424_;
	assign _06005_ = _06004_ | _02984_;
	assign _06006_ = _06005_ | _07758_;
	assign _06007_ = \mchip.index [11] & ~_06006_;
	assign _06008_ = _00302_ | _02984_;
	assign _06009_ = _06008_ | _02097_;
	assign _06010_ = _06009_ | \mchip.index [8];
	assign _06011_ = _06010_ | \mchip.index [9];
	assign _06012_ = \mchip.index [11] & ~_06011_;
	assign _06014_ = _02932_ | _07758_;
	assign _06015_ = _06014_ | \mchip.index [10];
	assign _06016_ = \mchip.index [11] & ~_06015_;
	assign _06017_ = _01173_ | _04648_;
	assign _06018_ = _01986_ & ~_06017_;
	assign _06019_ = _06556_ | \mchip.index [7];
	assign _06020_ = _06019_ | \mchip.index [8];
	assign _06021_ = \mchip.index [9] & ~_06020_;
	assign _06022_ = _02887_ | _07758_;
	assign _06023_ = \mchip.index [10] & ~_06022_;
	assign _06025_ = ~(_07711_ & \mchip.index [9]);
	assign _06026_ = \mchip.index [11] & ~_06025_;
	assign _06027_ = _00708_ | _04648_;
	assign _06028_ = _06027_ | _07758_;
	assign _06029_ = _06028_ | _01986_;
	assign _06030_ = _01875_ & ~_06029_;
	assign _06031_ = _01702_ | _04648_;
	assign _06032_ = _01986_ & ~_06031_;
	assign _06033_ = _07299_ | \mchip.index [7];
	assign _06034_ = _06033_ | \mchip.index [8];
	assign _06036_ = _06034_ | _07758_;
	assign _06037_ = \mchip.index [11] & ~_06036_;
	assign _06038_ = \mchip.index [10] & ~_01921_;
	assign _06039_ = _03540_ | _02984_;
	assign _06040_ = _06039_ | \mchip.index [7];
	assign _06041_ = _06040_ | _04648_;
	assign _06042_ = _06041_ | \mchip.index [9];
	assign _06043_ = \mchip.index [10] & ~_06042_;
	assign _06044_ = _04057_ | _01986_;
	assign _06045_ = _01875_ & ~_06044_;
	assign _06047_ = _06045_ | _06043_;
	assign _06048_ = _06047_ | _06038_;
	assign _06049_ = _06048_ | _06037_;
	assign _06050_ = _06049_ | _06032_;
	assign _06051_ = _06050_ | _03461_;
	assign _06052_ = _06051_ | _06030_;
	assign _06053_ = _06052_ | _06026_;
	assign _06054_ = _06053_ | _06023_;
	assign _06055_ = _06054_ | _06021_;
	assign _06056_ = _06055_ | _06018_;
	assign _06058_ = _06056_ | _06016_;
	assign _06059_ = _06058_ | _06012_;
	assign _06060_ = _06059_ | _06007_;
	assign _06061_ = _06060_ | _06003_;
	assign _06062_ = _06061_ | _02110_;
	assign _06063_ = _06062_ | _05997_;
	assign _06064_ = _06063_ | _05993_;
	assign _06065_ = _06064_ | _05989_;
	assign _06066_ = _06065_ | _05986_;
	assign _06067_ = _06066_ | _05984_;
	assign _06069_ = _06067_ | _05981_;
	assign _06070_ = _06069_ | _05975_;
	assign _06071_ = _06070_ | _05974_;
	assign _06072_ = _06071_ | _05971_;
	assign _06073_ = _06072_ | _05967_;
	assign _06074_ = _06073_ | _05963_;
	assign _06075_ = _06074_ | _05958_;
	assign _06076_ = _06075_ | _05955_;
	assign _06077_ = _06076_ | _05953_;
	assign _06078_ = _06077_ | _05952_;
	assign _06080_ = _06078_ | _05950_;
	assign _06081_ = _06080_ | _05947_;
	assign _06082_ = _06081_ | _05942_;
	assign _06083_ = _06082_ | _05940_;
	assign _06084_ = _06083_ | _05938_;
	assign _06085_ = _06084_ | _05933_;
	assign _06086_ = _06085_ | _05931_;
	assign _06087_ = _06086_ | _05928_;
	assign _06088_ = _06087_ | _05926_;
	assign _06089_ = _06088_ | _05921_;
	assign _06092_ = _06089_ | _05919_;
	assign _06093_ = _06092_ | _05915_;
	assign _06094_ = _06093_ | _05912_;
	assign _06095_ = _06094_ | _05908_;
	assign _06096_ = _06095_ | _03301_;
	assign _06097_ = _06096_ | _05907_;
	assign _06098_ = _06097_ | _05904_;
	assign _06099_ = _06098_ | _05900_;
	assign _06100_ = _06099_ | _05898_;
	assign _06101_ = _06100_ | _05892_;
	assign _06103_ = _06101_ | _05886_;
	assign _06104_ = _06103_ | _05883_;
	assign _06105_ = _06104_ | _05879_;
	assign _06106_ = _06105_ | _05876_;
	assign _06107_ = _06106_ | _05872_;
	assign _06108_ = _06107_ | _05867_;
	assign _06109_ = _06108_ | _05864_;
	assign _06110_ = _06109_ | _07694_;
	assign _06111_ = _06110_ | _05861_;
	assign _06112_ = _06111_ | _05859_;
	assign _06114_ = _06112_ | _05856_;
	assign _06115_ = _06114_ | _05852_;
	assign _06116_ = _06115_ | _05850_;
	assign _06117_ = _06116_ | _05847_;
	assign _06118_ = _06117_ | _05844_;
	assign _06119_ = _06118_ | _05841_;
	assign _06120_ = _06119_ | _05837_;
	assign _06121_ = _06120_ | _05834_;
	assign _06122_ = _06121_ | _05832_;
	assign _06123_ = _06122_ | _05830_;
	assign _06125_ = _06123_ | _05826_;
	assign _06126_ = _06125_ | _05823_;
	assign _06127_ = _06126_ | _05821_;
	assign _06128_ = _06127_ | _01907_;
	assign _06129_ = _06128_ | _05819_;
	assign _06130_ = _06129_ | _05815_;
	assign _06131_ = _06130_ | _05811_;
	assign _06132_ = _06131_ | _05807_;
	assign _06133_ = _06132_ | _05804_;
	assign _06134_ = _06133_ | _05800_;
	assign _06136_ = _06134_ | _05796_;
	assign _06137_ = _06136_ | _05790_;
	assign _06138_ = _06137_ | _05785_;
	assign _06139_ = _06138_ | _05778_;
	assign _06140_ = _06139_ | _05774_;
	assign _06141_ = _06140_ | _05771_;
	assign _06142_ = _06141_ | _05767_;
	assign _06143_ = _06142_ | _05764_;
	assign _06144_ = _06143_ | _05761_;
	assign _06145_ = _06144_ | _05760_;
	assign _06147_ = _06145_ | _05755_;
	assign _06148_ = _06147_ | _05751_;
	assign _06149_ = _06148_ | _05750_;
	assign _06150_ = _06149_ | _05749_;
	assign _06151_ = _06150_ | _05743_;
	assign _06152_ = _06151_ | _05740_;
	assign _06153_ = _06152_ | _05736_;
	assign _06154_ = _06153_ | _05733_;
	assign _06155_ = _06154_ | _05729_;
	assign _06156_ = _06155_ | _05725_;
	assign _06158_ = _06156_ | _05720_;
	assign _06159_ = _06158_ | _05715_;
	assign _06160_ = _06159_ | _05711_;
	assign _06161_ = _06160_ | _05709_;
	assign _06162_ = _06161_ | _05706_;
	assign _06163_ = _06162_ | _05701_;
	assign _06164_ = _06163_ | _05698_;
	assign _06165_ = _06164_ | _05694_;
	assign _06166_ = _06165_ | _05688_;
	assign _06167_ = _06166_ | _05685_;
	assign _06169_ = _06167_ | _05681_;
	assign _06170_ = _06169_ | _04299_;
	assign _06171_ = _06170_ | _05675_;
	assign _06172_ = _06171_ | _05673_;
	assign _06173_ = _06172_ | _05672_;
	assign _06174_ = _06173_ | _05671_;
	assign _06175_ = _06174_ | _05667_;
	assign _06176_ = _06175_ | _05665_;
	assign _06177_ = _06176_ | _05661_;
	assign _06178_ = _06177_ | _05660_;
	assign _06180_ = _06178_ | _05657_;
	assign _06181_ = _06180_ | _05654_;
	assign _06182_ = _06181_ | _05651_;
	assign _06183_ = _06182_ | _05648_;
	assign _06184_ = _06183_ | _05642_;
	assign _06185_ = _06184_ | _05639_;
	assign _06186_ = _06185_ | _05637_;
	assign _06187_ = _06186_ | _05631_;
	assign _06188_ = _06187_ | _05626_;
	assign _06189_ = _06188_ | _05621_;
	assign _06191_ = _06189_ | _05617_;
	assign _06192_ = _06191_ | _05614_;
	assign _06193_ = _06192_ | _05610_;
	assign _06194_ = _06193_ | _05605_;
	assign _06195_ = _06194_ | _05603_;
	assign _06196_ = _06195_ | _05596_;
	assign _06197_ = _06196_ | _05589_;
	assign _06198_ = _06197_ | _05586_;
	assign _06199_ = _06198_ | _05583_;
	assign _06200_ = _06199_ | _01707_;
	assign _06203_ = _06200_ | _05578_;
	assign _06204_ = _06203_ | _05573_;
	assign _06205_ = _06204_ | _05568_;
	assign _06206_ = _06205_ | _05566_;
	assign _06207_ = _06206_ | _05563_;
	assign _06208_ = _06207_ | _01660_;
	assign _06209_ = _06208_ | _05560_;
	assign _06210_ = _06209_ | _05557_;
	assign _06211_ = _06210_ | _05553_;
	assign _06212_ = _06211_ | _05552_;
	assign _06214_ = _06212_ | _05550_;
	assign _06215_ = _06214_ | _05544_;
	assign _06216_ = _06215_ | _05540_;
	assign _06217_ = _06216_ | _05534_;
	assign _06218_ = _06217_ | _05531_;
	assign _06219_ = _06218_ | _05528_;
	assign _06220_ = _06219_ | _05523_;
	assign _06221_ = _06220_ | _05519_;
	assign _06222_ = _06221_ | _05515_;
	assign _06223_ = _06222_ | _05511_;
	assign _06225_ = _06223_ | _05508_;
	assign _06226_ = _06225_ | _05506_;
	assign _06227_ = _06226_ | _05501_;
	assign _06228_ = _06227_ | _05499_;
	assign _06229_ = _06228_ | _05495_;
	assign _06230_ = _06229_ | _05493_;
	assign _06231_ = _06230_ | _05489_;
	assign _06232_ = _06231_ | _05487_;
	assign _06233_ = _06232_ | _01557_;
	assign _06234_ = _06233_ | _05483_;
	assign _06236_ = _06234_ | _05481_;
	assign _06237_ = _06236_ | _05477_;
	assign _06238_ = _06237_ | _05472_;
	assign _06239_ = _06238_ | _05468_;
	assign _06240_ = _06239_ | _05463_;
	assign _06241_ = _06240_ | _05461_;
	assign _06242_ = _06241_ | _05457_;
	assign _06243_ = _06242_ | _05454_;
	assign _06244_ = _06243_ | _05449_;
	assign _06245_ = _06244_ | _05444_;
	assign _06247_ = _06245_ | _05441_;
	assign _06248_ = _06247_ | _05438_;
	assign _06249_ = _06248_ | _05432_;
	assign _06250_ = _06249_ | _05428_;
	assign _06251_ = _06250_ | _05421_;
	assign _06252_ = _06251_ | _05417_;
	assign _06253_ = _06252_ | _05412_;
	assign _06254_ = _06253_ | _05409_;
	assign _06255_ = _06254_ | _05405_;
	assign _06256_ = _06255_ | _05399_;
	assign _06258_ = _06256_ | _05397_;
	assign _06259_ = _06258_ | _05394_;
	assign _06260_ = _06259_ | _05389_;
	assign _06261_ = _06260_ | _04059_;
	assign _06262_ = _06261_ | _05386_;
	assign _06263_ = _06262_ | _05382_;
	assign _06264_ = _06263_ | _05378_;
	assign _06265_ = _06264_ | _05376_;
	assign _06266_ = _06265_ | _04050_;
	assign _06267_ = _06266_ | _05372_;
	assign _06269_ = _06267_ | _05367_;
	assign _06270_ = _06269_ | _05363_;
	assign _06271_ = _06270_ | _05356_;
	assign _06272_ = _06271_ | _05352_;
	assign _06273_ = _06272_ | _05349_;
	assign _06274_ = _06273_ | _05346_;
	assign _06275_ = _06274_ | _05340_;
	assign _06276_ = _06275_ | _05338_;
	assign _06277_ = _06276_ | _05333_;
	assign _06278_ = _06277_ | _05330_;
	assign _06280_ = _06278_ | _05327_;
	assign _06281_ = _06280_ | _05322_;
	assign _06282_ = _06281_ | _05317_;
	assign _06283_ = _06282_ | _05311_;
	assign _06284_ = _06283_ | _01396_;
	assign _06285_ = _06284_ | _05307_;
	assign _06286_ = _06285_ | _05303_;
	assign _06287_ = _06286_ | _05297_;
	assign _06288_ = _06287_ | _05292_;
	assign _06289_ = _06288_ | _05289_;
	assign _06291_ = _06289_ | _05285_;
	assign _06292_ = _06291_ | _05283_;
	assign _06293_ = _06292_ | _05279_;
	assign _06294_ = _06293_ | _05275_;
	assign _06295_ = _06294_ | _05271_;
	assign _06296_ = _06295_ | _05267_;
	assign _06297_ = _06296_ | _05263_;
	assign _06298_ = _06297_ | _05261_;
	assign _06299_ = _06298_ | _05257_;
	assign _06300_ = _06299_ | _05252_;
	assign _06302_ = _06300_ | _05245_;
	assign _06303_ = _06302_ | _05240_;
	assign _06304_ = _06303_ | _05235_;
	assign _06305_ = _06304_ | _05231_;
	assign _06306_ = _06305_ | _05228_;
	assign _06307_ = _06306_ | _05221_;
	assign _06308_ = _06307_ | _05217_;
	assign _06309_ = _06308_ | _05212_;
	assign _06310_ = _06309_ | _05210_;
	assign _06311_ = _06310_ | _05206_;
	assign _06314_ = _06311_ | _05200_;
	assign _06315_ = _06314_ | _05198_;
	assign _06316_ = _06315_ | _05195_;
	assign _06317_ = _06316_ | _05192_;
	assign _06318_ = _06317_ | _05185_;
	assign _06319_ = _06318_ | _05182_;
	assign _06320_ = _06319_ | _05176_;
	assign _06321_ = _06320_ | _05171_;
	assign _06322_ = _06321_ | _05164_;
	assign _06323_ = _06322_ | _02483_;
	assign _06325_ = _06323_ | _05161_;
	assign _06326_ = _06325_ | _03089_;
	assign _06327_ = _06326_ | _05157_;
	assign _06328_ = _06327_ | _05153_;
	assign _06329_ = _06328_ | _05150_;
	assign _06330_ = _06329_ | _05144_;
	assign _06331_ = _06330_ | _05140_;
	assign _06332_ = _06331_ | _05135_;
	assign _06333_ = _06332_ | _05132_;
	assign _06334_ = _06333_ | _05130_;
	assign _06336_ = _06334_ | _05124_;
	assign _06337_ = _06336_ | _05120_;
	assign _06338_ = _06337_ | _05112_;
	assign _06339_ = _06338_ | _05109_;
	assign _06340_ = _06339_ | _05108_;
	assign _06341_ = _06340_ | _05104_;
	assign _06342_ = _06341_ | _05101_;
	assign _06343_ = _06342_ | _05098_;
	assign _06344_ = _06343_ | _05094_;
	assign _06345_ = _06344_ | _05088_;
	assign _06347_ = _06345_ | _05085_;
	assign _06348_ = _06347_ | _03071_;
	assign \mchip.val [1] = _06348_ | _02448_;
	assign _06349_ = _01472_ | _07758_;
	assign _06350_ = _01986_ & ~_06349_;
	assign _06351_ = _00681_ | \mchip.index [6];
	assign _06352_ = _06351_ | \mchip.index [7];
	assign _06353_ = _06352_ | \mchip.index [9];
	assign _06354_ = _01875_ & ~_06353_;
	assign _06355_ = _00329_ | \mchip.index [6];
	assign _06357_ = _06355_ | \mchip.index [7];
	assign _06358_ = _06357_ | _04648_;
	assign _06359_ = _06358_ | _07758_;
	assign _06360_ = _01875_ & ~_06359_;
	assign _06361_ = _04174_ | \mchip.index [8];
	assign _06362_ = _01875_ & ~_06361_;
	assign _06363_ = _02100_ | \mchip.index [9];
	assign _06364_ = \mchip.index [10] & ~_06363_;
	assign _06365_ = _07322_ | \mchip.index [9];
	assign _06366_ = \mchip.index [10] & ~_06365_;
	assign _06368_ = _02743_ | _02097_;
	assign _06369_ = _06368_ | _04648_;
	assign _06370_ = _01986_ & ~_06369_;
	assign _06371_ = _01290_ | _02984_;
	assign _06372_ = _06371_ | _02097_;
	assign _06373_ = _06372_ | \mchip.index [9];
	assign _06374_ = \mchip.index [10] & ~_06373_;
	assign _06375_ = _02031_ | _02097_;
	assign _06376_ = _06375_ | \mchip.index [8];
	assign _06377_ = \mchip.index [10] & ~_06376_;
	assign _06379_ = \mchip.index [10] & ~_03839_;
	assign _06380_ = _01189_ | \mchip.index [5];
	assign _06381_ = _06380_ | _02984_;
	assign _06382_ = _06381_ | \mchip.index [7];
	assign _06383_ = _06382_ | _01986_;
	assign _06384_ = \mchip.index [11] & ~_06383_;
	assign _06385_ = _05943_ | \mchip.index [9];
	assign _06386_ = \mchip.index [10] & ~_06385_;
	assign _06387_ = _03029_ | \mchip.index [5];
	assign _06388_ = _06387_ | _02984_;
	assign _06390_ = _06388_ | _01986_;
	assign _06391_ = \mchip.index [11] & ~_06390_;
	assign _06392_ = _01561_ | _02984_;
	assign _06393_ = _06392_ | \mchip.index [7];
	assign _06394_ = _06393_ | _04648_;
	assign _06395_ = _06394_ | \mchip.index [9];
	assign _06396_ = \mchip.index [10] & ~_06395_;
	assign _06397_ = _02819_ | _04648_;
	assign _06398_ = _01875_ & ~_06397_;
	assign _06399_ = _02943_ | \mchip.index [9];
	assign _06401_ = \mchip.index [11] & ~_06399_;
	assign _06402_ = _00781_ | _02097_;
	assign _06403_ = _06402_ | _04648_;
	assign _06404_ = _06403_ | \mchip.index [9];
	assign _06405_ = _01875_ & ~_06404_;
	assign _06406_ = _00352_ | _05424_;
	assign _06407_ = \mchip.index [7] & ~_06406_;
	assign _06408_ = _00415_ | \mchip.index [7];
	assign _06409_ = _06408_ | _04648_;
	assign _06410_ = _06409_ | \mchip.index [9];
	assign _06412_ = \mchip.index [10] & ~_06410_;
	assign _06413_ = _03165_ | \mchip.index [7];
	assign _06414_ = _06413_ | \mchip.index [9];
	assign _06415_ = \mchip.index [10] & ~_06414_;
	assign _06416_ = _04762_ | _02097_;
	assign _06417_ = _06416_ | \mchip.index [8];
	assign _06418_ = _07758_ & ~_06417_;
	assign _06419_ = _04143_ | _02984_;
	assign _06420_ = _06419_ | _02097_;
	assign _06421_ = _06420_ | _04648_;
	assign _06424_ = _06421_ | \mchip.index [9];
	assign _06425_ = \mchip.index [11] & ~_06424_;
	assign _06426_ = _07758_ & ~_02544_;
	assign _06427_ = _05434_ | _07758_;
	assign _06428_ = _01986_ & ~_06427_;
	assign _06429_ = _02696_ | \mchip.index [7];
	assign _06430_ = _06429_ | \mchip.index [8];
	assign _06431_ = _06430_ | \mchip.index [10];
	assign _06432_ = _01875_ & ~_06431_;
	assign _06433_ = _01152_ | _05424_;
	assign _06435_ = _06433_ | \mchip.index [7];
	assign _06436_ = _06435_ | _04648_;
	assign _06437_ = \mchip.index [11] & ~_06436_;
	assign _06438_ = _04741_ | _05424_;
	assign _06439_ = _06438_ | _02984_;
	assign _06440_ = _06439_ | \mchip.index [7];
	assign _06441_ = \mchip.index [10] & ~_06440_;
	assign _06442_ = _00703_ | _07758_;
	assign _06443_ = _01986_ & ~_06442_;
	assign _06444_ = _02810_ | _04648_;
	assign _06446_ = _07758_ & ~_06444_;
	assign _06447_ = \mchip.index [10] & ~_02721_;
	assign _06448_ = _01179_ | _02097_;
	assign _06449_ = _06448_ | _04648_;
	assign _06450_ = _01986_ & ~_06449_;
	assign _06451_ = _05957_ | \mchip.index [6];
	assign _06452_ = _06451_ | _02097_;
	assign _06453_ = _06452_ | \mchip.index [8];
	assign _06454_ = \mchip.index [11] & ~_06453_;
	assign _06455_ = _05059_ | _02097_;
	assign _06457_ = _06455_ | _04648_;
	assign _06458_ = _06457_ | \mchip.index [9];
	assign _06459_ = \mchip.index [10] & ~_06458_;
	assign _06460_ = _00587_ | _02097_;
	assign _06461_ = _06460_ | _04648_;
	assign _06462_ = _06461_ | \mchip.index [9];
	assign _06463_ = \mchip.index [10] & ~_06462_;
	assign _06464_ = _05494_ | _01986_;
	assign _06465_ = _01875_ & ~_06464_;
	assign _06466_ = _05451_ | _07758_;
	assign _06468_ = \mchip.index [10] & ~_06466_;
	assign _06469_ = _01359_ | \mchip.index [7];
	assign _06470_ = _06469_ | _07758_;
	assign _06471_ = _01875_ & ~_06470_;
	assign _06472_ = _00692_ | _07758_;
	assign _06473_ = \mchip.index [11] & ~_06472_;
	assign _06474_ = _03043_ | _01986_;
	assign _06475_ = \mchip.index [11] & ~_06474_;
	assign _06476_ = _02175_ | _02097_;
	assign _06477_ = _06476_ | \mchip.index [8];
	assign _06479_ = _06477_ | \mchip.index [9];
	assign _06480_ = \mchip.index [10] & ~_06479_;
	assign _06481_ = _00099_ | _05424_;
	assign _06482_ = _06481_ | _04648_;
	assign _06483_ = _06482_ | _01986_;
	assign _06484_ = _01875_ & ~_06483_;
	assign _06485_ = _04769_ | \mchip.index [9];
	assign _06486_ = _01986_ & ~_06485_;
	assign _06487_ = _06689_ | _05424_;
	assign _06488_ = _06487_ | \mchip.index [6];
	assign _06490_ = _06488_ | \mchip.index [7];
	assign _06491_ = _06490_ | _01986_;
	assign _06492_ = \mchip.index [11] & ~_06491_;
	assign _06493_ = _01819_ | \mchip.index [9];
	assign _06494_ = \mchip.index [10] & ~_06493_;
	assign _06495_ = _03998_ | _04648_;
	assign _06496_ = _01986_ & ~_06495_;
	assign _06497_ = _03200_ | _02097_;
	assign _06498_ = _06497_ | \mchip.index [10];
	assign _06499_ = \mchip.index [11] & ~_06498_;
	assign _06501_ = _01986_ & ~_03476_;
	assign _06502_ = _03651_ | _07758_;
	assign _06503_ = _01986_ & ~_06502_;
	assign _06504_ = _01535_ | _02097_;
	assign _06505_ = \mchip.index [9] & ~_06504_;
	assign _06506_ = \mchip.index [10] & ~_04440_;
	assign _06507_ = _01099_ | \mchip.index [7];
	assign _06508_ = _06507_ | _04648_;
	assign _06509_ = _06508_ | _07758_;
	assign _06510_ = _06509_ | \mchip.index [10];
	assign _06512_ = _01875_ & ~_06510_;
	assign _06513_ = _02016_ | \mchip.index [8];
	assign _06514_ = \mchip.index [9] & ~_06513_;
	assign _06515_ = _00299_ | _02984_;
	assign _06516_ = _06515_ | _04648_;
	assign _06517_ = _07758_ & ~_06516_;
	assign _06518_ = _03291_ | \mchip.index [8];
	assign _06519_ = \mchip.index [9] & ~_06518_;
	assign _06520_ = _01364_ | \mchip.index [8];
	assign _06521_ = \mchip.index [9] & ~_06520_;
	assign _06523_ = _01966_ | \mchip.index [9];
	assign _06524_ = \mchip.index [11] & ~_06523_;
	assign _06525_ = _03260_ | _04648_;
	assign _06526_ = _06525_ | \mchip.index [10];
	assign _06527_ = \mchip.index [11] & ~_06526_;
	assign _06528_ = _01970_ | \mchip.index [8];
	assign _06529_ = _06528_ | \mchip.index [9];
	assign _06530_ = \mchip.index [11] & ~_06529_;
	assign _06531_ = _01986_ & ~_04513_;
	assign _06532_ = _04628_ | _07758_;
	assign _06535_ = _01986_ & ~_06532_;
	assign _06536_ = _02897_ | \mchip.index [8];
	assign _06537_ = \mchip.index [10] & ~_06536_;
	assign _06538_ = _05628_ | _04648_;
	assign _06539_ = _06538_ | _07758_;
	assign _06540_ = _06539_ | _01986_;
	assign _06541_ = _01875_ & ~_06540_;
	assign _06542_ = _05964_ | _07758_;
	assign _06543_ = _06542_ | \mchip.index [10];
	assign _06544_ = _01875_ & ~_06543_;
	assign _06546_ = _03877_ | \mchip.index [7];
	assign _06547_ = _06546_ | \mchip.index [8];
	assign _06548_ = _06547_ | \mchip.index [9];
	assign _06549_ = \mchip.index [10] & ~_06548_;
	assign _06550_ = _02966_ | \mchip.index [8];
	assign _06551_ = \mchip.index [11] & ~_06550_;
	assign _06552_ = _01196_ | \mchip.index [6];
	assign _06553_ = _06552_ | \mchip.index [8];
	assign _06554_ = _06553_ | _07758_;
	assign _06555_ = \mchip.index [11] & ~_06554_;
	assign _06557_ = _01774_ | _02097_;
	assign _06558_ = _06557_ | \mchip.index [9];
	assign _06559_ = _01986_ & ~_06558_;
	assign _06560_ = _07720_ | \mchip.index [8];
	assign _06561_ = _06560_ | _07758_;
	assign _06562_ = _06561_ | \mchip.index [10];
	assign _06563_ = _01875_ & ~_06562_;
	assign _06564_ = _01387_ | _04648_;
	assign _06565_ = _06564_ | \mchip.index [9];
	assign _06566_ = _01875_ & ~_06565_;
	assign _06568_ = _01647_ | _04648_;
	assign _06569_ = _06568_ | _07758_;
	assign _06570_ = \mchip.index [10] & ~_06569_;
	assign _06571_ = _01320_ | \mchip.index [6];
	assign _06572_ = _06571_ | \mchip.index [8];
	assign _06573_ = _06572_ | _07758_;
	assign _06574_ = _06573_ | \mchip.index [10];
	assign _06575_ = _01875_ & ~_06574_;
	assign _06576_ = _01717_ | _07758_;
	assign _06577_ = _01986_ & ~_06576_;
	assign _06579_ = _00530_ | _02097_;
	assign _06580_ = _06579_ | _01986_;
	assign _06581_ = \mchip.index [11] & ~_06580_;
	assign _06582_ = _02320_ | _02984_;
	assign _06583_ = _06582_ | \mchip.index [9];
	assign _06584_ = \mchip.index [11] & ~_06583_;
	assign _06585_ = _00422_ | _04648_;
	assign _06586_ = _06585_ | \mchip.index [9];
	assign _06587_ = \mchip.index [10] & ~_06586_;
	assign _06588_ = _01618_ | \mchip.index [6];
	assign _06590_ = _06588_ | _02097_;
	assign _06591_ = _06590_ | \mchip.index [8];
	assign _06592_ = \mchip.index [9] & ~_06591_;
	assign _06593_ = _03209_ | \mchip.index [8];
	assign _06594_ = \mchip.index [11] & ~_06593_;
	assign _06595_ = _01451_ | _04648_;
	assign _06596_ = _01875_ & ~_06595_;
	assign _06597_ = _01791_ | \mchip.index [9];
	assign _06598_ = _06597_ | \mchip.index [10];
	assign _06599_ = _01875_ & ~_06598_;
	assign _06601_ = _03923_ | _07758_;
	assign _06602_ = _01986_ & ~_06601_;
	assign _06603_ = _01337_ | _04648_;
	assign _06604_ = _06603_ | _07758_;
	assign _06605_ = _01986_ & ~_06604_;
	assign _06606_ = _01230_ | \mchip.index [7];
	assign _06607_ = _06606_ | \mchip.index [8];
	assign _06608_ = _06607_ | \mchip.index [10];
	assign _06609_ = _01875_ & ~_06608_;
	assign _06610_ = _00771_ | \mchip.index [10];
	assign _06612_ = _01875_ & ~_06610_;
	assign _06613_ = _05445_ | \mchip.index [6];
	assign _06614_ = _06613_ | _02097_;
	assign _06615_ = _06614_ | \mchip.index [8];
	assign _06616_ = _06615_ | \mchip.index [9];
	assign _06617_ = \mchip.index [10] & ~_06616_;
	assign _06618_ = _03371_ | \mchip.index [8];
	assign _06619_ = _06618_ | _07758_;
	assign _06620_ = \mchip.index [10] & ~_06619_;
	assign _06621_ = _07720_ | \mchip.index [5];
	assign _06623_ = _06621_ | \mchip.index [6];
	assign _06624_ = _06623_ | \mchip.index [7];
	assign _06625_ = _06624_ | \mchip.index [8];
	assign _06626_ = _06625_ | _07758_;
	assign _06627_ = \mchip.index [11] & ~_06626_;
	assign _06628_ = _01986_ & ~_03326_;
	assign _06629_ = _04577_ | \mchip.index [7];
	assign _06630_ = _06629_ | \mchip.index [8];
	assign _06631_ = \mchip.index [10] & ~_06630_;
	assign _06632_ = _05354_ | _07758_;
	assign _06634_ = \mchip.index [10] & ~_06632_;
	assign _06635_ = _00318_ | _01098_;
	assign _06636_ = _06635_ | _02984_;
	assign _06637_ = _06636_ | \mchip.index [7];
	assign _06638_ = _06637_ | \mchip.index [8];
	assign _06639_ = _06638_ | \mchip.index [9];
	assign _06640_ = \mchip.index [10] & ~_06639_;
	assign _06641_ = _00662_ | \mchip.index [5];
	assign _06642_ = _06641_ | _02984_;
	assign _06643_ = _06642_ | _07758_;
	assign _06646_ = _06643_ | \mchip.index [10];
	assign _06647_ = _01875_ & ~_06646_;
	assign _06648_ = _04131_ | _04648_;
	assign _06649_ = _06648_ | \mchip.index [10];
	assign _06650_ = \mchip.index [11] & ~_06649_;
	assign _06651_ = _01220_ | \mchip.index [10];
	assign _06652_ = _01875_ & ~_06651_;
	assign _06653_ = _03057_ | \mchip.index [7];
	assign _06654_ = _06653_ | \mchip.index [8];
	assign _06655_ = \mchip.index [9] & ~_06654_;
	assign _06657_ = _00351_ | \mchip.index [7];
	assign _06658_ = _06657_ | \mchip.index [8];
	assign _06659_ = _06658_ | _07758_;
	assign _06660_ = _06659_ | \mchip.index [10];
	assign _06661_ = \mchip.index [11] & ~_06660_;
	assign _06662_ = _07199_ | \mchip.index [5];
	assign _06663_ = _06662_ | \mchip.index [7];
	assign _06664_ = _06663_ | \mchip.index [9];
	assign _06665_ = \mchip.index [11] & ~_06664_;
	assign _06666_ = _05880_ | \mchip.index [8];
	assign _06668_ = _06666_ | _07758_;
	assign _06669_ = _01986_ & ~_06668_;
	assign _06670_ = _02595_ | _01986_;
	assign _06671_ = _01875_ & ~_06670_;
	assign _06672_ = _00380_ | _05424_;
	assign _06673_ = _06672_ | \mchip.index [6];
	assign _06674_ = _06673_ | _01986_;
	assign _06675_ = \mchip.index [11] & ~_06674_;
	assign _06676_ = _06515_ | \mchip.index [7];
	assign _06677_ = _06676_ | _04648_;
	assign _06679_ = _06677_ | _01986_;
	assign _06680_ = _01875_ & ~_06679_;
	assign _06681_ = _01528_ | _02097_;
	assign _06682_ = _06681_ | \mchip.index [8];
	assign _06683_ = _06682_ | \mchip.index [10];
	assign _06684_ = \mchip.index [11] & ~_06683_;
	assign _06685_ = _01244_ | _02097_;
	assign _06686_ = _06685_ | _04648_;
	assign _06687_ = _06686_ | _07758_;
	assign _06688_ = \mchip.index [10] & ~_06687_;
	assign _06690_ = _02320_ | \mchip.index [7];
	assign _06691_ = _06690_ | \mchip.index [8];
	assign _06692_ = _06691_ | \mchip.index [9];
	assign _06693_ = \mchip.index [11] & ~_06692_;
	assign _06694_ = _04399_ | \mchip.index [8];
	assign _06695_ = _06694_ | _07758_;
	assign _06696_ = \mchip.index [10] & ~_06695_;
	assign _06697_ = _02021_ | \mchip.index [8];
	assign _06698_ = \mchip.index [11] & ~_06697_;
	assign _06699_ = _02231_ | _04648_;
	assign _06701_ = \mchip.index [9] & ~_06699_;
	assign _06702_ = _04449_ | _02097_;
	assign _06703_ = _06702_ | \mchip.index [8];
	assign _06704_ = \mchip.index [10] & ~_06703_;
	assign _06705_ = _01925_ | \mchip.index [8];
	assign _06706_ = _06705_ | _07758_;
	assign _06707_ = \mchip.index [10] & ~_06706_;
	assign _06708_ = _01380_ | _04648_;
	assign _06709_ = \mchip.index [11] & ~_06708_;
	assign _06710_ = _06635_ | \mchip.index [5];
	assign _06712_ = _06710_ | _02984_;
	assign _06713_ = _06712_ | _02097_;
	assign _06714_ = _06713_ | _04648_;
	assign _06715_ = _06714_ | _01986_;
	assign _06716_ = _01875_ & ~_06715_;
	assign _06717_ = _04449_ | \mchip.index [8];
	assign _06718_ = _06717_ | _07758_;
	assign _06719_ = \mchip.index [10] & ~_06718_;
	assign _06720_ = _01427_ | \mchip.index [8];
	assign _06721_ = _06720_ | \mchip.index [10];
	assign _06723_ = _01875_ & ~_06721_;
	assign _06724_ = _00000_ | \mchip.index [8];
	assign _06725_ = _06724_ | _07758_;
	assign _06726_ = _06725_ | \mchip.index [10];
	assign _06727_ = _01875_ & ~_06726_;
	assign _06728_ = _02975_ | \mchip.index [6];
	assign _06729_ = _06728_ | _04648_;
	assign _06730_ = _06729_ | _01986_;
	assign _06731_ = _01875_ & ~_06730_;
	assign _06732_ = _01359_ | _04648_;
	assign _06734_ = _06732_ | \mchip.index [10];
	assign _06735_ = _01875_ & ~_06734_;
	assign _06736_ = _01986_ & ~_05102_;
	assign _06737_ = _06090_ | _02097_;
	assign _06738_ = _06737_ | \mchip.index [8];
	assign _06739_ = _06738_ | \mchip.index [9];
	assign _06740_ = _01875_ & ~_06739_;
	assign _06741_ = _00541_ | \mchip.index [6];
	assign _06742_ = _06741_ | \mchip.index [7];
	assign _06743_ = _06742_ | _04648_;
	assign _06745_ = _06743_ | \mchip.index [10];
	assign _06746_ = \mchip.index [11] & ~_06745_;
	assign _06747_ = _00311_ | _02984_;
	assign _06748_ = _06747_ | _02097_;
	assign _06749_ = _06748_ | \mchip.index [8];
	assign _06750_ = _06749_ | _07758_;
	assign _06751_ = \mchip.index [10] & ~_06750_;
	assign _06752_ = _07714_ | \mchip.index [6];
	assign _06753_ = _06752_ | _02097_;
	assign _06754_ = _06753_ | _04648_;
	assign _06757_ = _06754_ | \mchip.index [9];
	assign _06758_ = _06757_ | \mchip.index [10];
	assign _06759_ = _01875_ & ~_06758_;
	assign _06760_ = _04310_ | \mchip.index [8];
	assign _06761_ = \mchip.index [11] & ~_06760_;
	assign _06762_ = _00267_ | _02984_;
	assign _06763_ = _06762_ | _02097_;
	assign _06764_ = _06763_ | _04648_;
	assign _06765_ = _06764_ | \mchip.index [9];
	assign _06766_ = \mchip.index [11] & ~_06765_;
	assign _06768_ = _02122_ | \mchip.index [7];
	assign _06769_ = _06768_ | _07758_;
	assign _06770_ = _06769_ | _01986_;
	assign _06771_ = _01875_ & ~_06770_;
	assign _06772_ = _06578_ | _05424_;
	assign _06773_ = _06772_ | _02984_;
	assign _06774_ = \mchip.index [11] & ~_06773_;
	assign _06775_ = _03212_ | _04648_;
	assign _06776_ = _06775_ | \mchip.index [9];
	assign _06777_ = \mchip.index [11] & ~_06776_;
	assign _06779_ = _04744_ | \mchip.index [8];
	assign _06780_ = _06779_ | \mchip.index [9];
	assign _06781_ = _01986_ & ~_06780_;
	assign _06782_ = _02884_ | \mchip.index [7];
	assign _06783_ = _06782_ | _04648_;
	assign _06784_ = _06783_ | _07758_;
	assign _06785_ = _01875_ & ~_06784_;
	assign _06786_ = _01620_ | _05424_;
	assign _06787_ = _06786_ | _02984_;
	assign _06788_ = _06787_ | _02097_;
	assign _06790_ = _06788_ | _04648_;
	assign _06791_ = _06790_ | _01986_;
	assign _06792_ = _01875_ & ~_06791_;
	assign _06793_ = _06585_ | _07758_;
	assign _06794_ = _01986_ & ~_06793_;
	assign _06795_ = _03960_ | _02984_;
	assign _06796_ = _06795_ | _02097_;
	assign _06797_ = _06796_ | \mchip.index [8];
	assign _06798_ = _06797_ | \mchip.index [9];
	assign _06799_ = \mchip.index [11] & ~_06798_;
	assign _06801_ = _07677_ | _02097_;
	assign _06802_ = _06801_ | _07758_;
	assign _06803_ = _01986_ & ~_06802_;
	assign _06804_ = _03739_ | _02097_;
	assign _06805_ = _06804_ | _04648_;
	assign _06806_ = _06805_ | \mchip.index [9];
	assign _06807_ = _06806_ | \mchip.index [10];
	assign _06808_ = _01875_ & ~_06807_;
	assign _06809_ = _05246_ | \mchip.index [6];
	assign _06810_ = _06809_ | _02097_;
	assign _06812_ = _06810_ | \mchip.index [8];
	assign _06813_ = _06812_ | \mchip.index [9];
	assign _06814_ = \mchip.index [11] & ~_06813_;
	assign _06815_ = _01111_ | \mchip.index [7];
	assign _06816_ = _06815_ | _04648_;
	assign _06817_ = _06816_ | _01986_;
	assign _06818_ = _01875_ & ~_06817_;
	assign _06819_ = _01207_ | _04648_;
	assign _06820_ = _06819_ | \mchip.index [9];
	assign _06821_ = _06820_ | \mchip.index [10];
	assign _06823_ = _01875_ & ~_06821_;
	assign _06824_ = _02154_ | _01986_;
	assign _06825_ = _01875_ & ~_06824_;
	assign _06826_ = _01938_ | _04648_;
	assign _06827_ = _06826_ | _07758_;
	assign _06828_ = _06827_ | _01986_;
	assign _06829_ = _01875_ & ~_06828_;
	assign _06830_ = _02481_ | \mchip.index [8];
	assign _06831_ = _06830_ | \mchip.index [9];
	assign _06832_ = _01986_ & ~_06831_;
	assign _06834_ = _01875_ & ~_05416_;
	assign _06835_ = _07758_ & ~_01273_;
	assign _06836_ = _02034_ | \mchip.index [7];
	assign _06837_ = \mchip.index [11] & ~_06836_;
	assign _06838_ = _07588_ | _02984_;
	assign _06839_ = _06838_ | \mchip.index [7];
	assign _06840_ = _06839_ | \mchip.index [9];
	assign _06841_ = \mchip.index [11] & ~_06840_;
	assign _06842_ = _01908_ | _02984_;
	assign _06843_ = _06842_ | \mchip.index [8];
	assign _06845_ = _06843_ | \mchip.index [9];
	assign _06846_ = \mchip.index [11] & ~_06845_;
	assign _06847_ = _01986_ & ~_04554_;
	assign _06848_ = _02479_ | _07758_;
	assign _06849_ = _01875_ & ~_06848_;
	assign _06850_ = _07758_ & ~_01478_;
	assign _06851_ = _00631_ | _02097_;
	assign _06852_ = _06851_ | \mchip.index [8];
	assign _06853_ = _06852_ | _07758_;
	assign _06854_ = _01875_ & ~_06853_;
	assign _06856_ = _07821_ | _05424_;
	assign _06857_ = _02984_ & ~_06856_;
	assign _06858_ = _04310_ | \mchip.index [7];
	assign _06859_ = _07758_ & ~_06858_;
	assign _06860_ = \mchip.index [11] & ~_02880_;
	assign _06861_ = _01347_ | _02097_;
	assign _06862_ = _06861_ | _01986_;
	assign _06863_ = \mchip.index [11] & ~_06862_;
	assign _06864_ = _06635_ | \mchip.index [6];
	assign _06865_ = _06864_ | \mchip.index [7];
	assign _06868_ = _06865_ | \mchip.index [8];
	assign _06869_ = _06868_ | _07758_;
	assign _06870_ = \mchip.index [10] & ~_06869_;
	assign _06871_ = _01875_ & ~_05840_;
	assign _06872_ = _07783_ | \mchip.index [9];
	assign _06873_ = _06872_ | \mchip.index [10];
	assign _06874_ = _01875_ & ~_06873_;
	assign _06875_ = _05302_ | _02097_;
	assign _06876_ = _06875_ | _04648_;
	assign _06877_ = _06876_ | _07758_;
	assign _06879_ = _01875_ & ~_06877_;
	assign _06880_ = _01958_ | _02097_;
	assign _06881_ = _06880_ | \mchip.index [9];
	assign _06882_ = _06881_ | _01986_;
	assign _06883_ = _01875_ & ~_06882_;
	assign _06884_ = \mchip.index [10] & ~_06005_;
	assign _06885_ = _01462_ | _02097_;
	assign _06886_ = _06885_ | _04648_;
	assign _06887_ = _06886_ | \mchip.index [9];
	assign _06888_ = _01875_ & ~_06887_;
	assign _06890_ = _00879_ | _05424_;
	assign _06891_ = _06890_ | \mchip.index [8];
	assign _06892_ = \mchip.index [9] & ~_06891_;
	assign _06893_ = _04639_ | _04648_;
	assign _06894_ = _06893_ | \mchip.index [9];
	assign _06895_ = _06894_ | \mchip.index [10];
	assign _06896_ = _01875_ & ~_06895_;
	assign _06897_ = _04572_ | _01986_;
	assign _06898_ = \mchip.index [11] & ~_06897_;
	assign _06899_ = _00688_ | _07758_;
	assign _06901_ = \mchip.index [11] & ~_06899_;
	assign _06902_ = _04549_ | \mchip.index [8];
	assign _06903_ = _06902_ | _07758_;
	assign _06904_ = \mchip.index [11] & ~_06903_;
	assign _06905_ = _03628_ | \mchip.index [7];
	assign _06906_ = _06905_ | _07758_;
	assign _06907_ = _01875_ & ~_06906_;
	assign _06908_ = _00435_ & ~\mchip.index [11];
	assign _06909_ = _01814_ | \mchip.index [8];
	assign _06910_ = _06909_ | \mchip.index [9];
	assign _06912_ = \mchip.index [10] & ~_06910_;
	assign _06913_ = _06589_ | _04648_;
	assign _06914_ = _06913_ | \mchip.index [9];
	assign _06915_ = _06914_ | \mchip.index [10];
	assign _06916_ = _01875_ & ~_06915_;
	assign _06917_ = _01797_ | \mchip.index [7];
	assign _06918_ = _06917_ | _01986_;
	assign _06919_ = \mchip.index [11] & ~_06918_;
	assign _06920_ = _00209_ | \mchip.index [6];
	assign _06921_ = _06920_ | \mchip.index [7];
	assign _06923_ = _06921_ | \mchip.index [8];
	assign _06924_ = _07758_ & ~_06923_;
	assign _06925_ = _06641_ | _02097_;
	assign _06926_ = _06925_ | \mchip.index [9];
	assign _06927_ = \mchip.index [11] & ~_06926_;
	assign _06928_ = _07646_ | _02097_;
	assign _06929_ = _06928_ | _04648_;
	assign _06930_ = _06929_ | \mchip.index [9];
	assign _06931_ = \mchip.index [11] & ~_06930_;
	assign _06932_ = _04460_ | _07758_;
	assign _06934_ = \mchip.index [11] & ~_06932_;
	assign _06935_ = _07310_ | \mchip.index [6];
	assign _06936_ = _06935_ | \mchip.index [7];
	assign _06937_ = _04648_ & ~_06936_;
	assign _06938_ = _02191_ | _02097_;
	assign _06939_ = _06938_ | \mchip.index [9];
	assign _06940_ = _06939_ | \mchip.index [10];
	assign _06941_ = _01875_ & ~_06940_;
	assign _06942_ = _02231_ | \mchip.index [10];
	assign _06943_ = _01875_ & ~_06942_;
	assign _06945_ = _06301_ | \mchip.index [8];
	assign _06946_ = _06945_ | \mchip.index [10];
	assign _06947_ = _01875_ & ~_06946_;
	assign _06948_ = _06756_ | _02097_;
	assign _06949_ = _06948_ | _07758_;
	assign _06950_ = \mchip.index [10] & ~_06949_;
	assign _06951_ = _03439_ | \mchip.index [8];
	assign _06952_ = _06951_ | _07758_;
	assign _06953_ = \mchip.index [10] & ~_06952_;
	assign _06954_ = _02990_ | _07758_;
	assign _06956_ = \mchip.index [11] & ~_06954_;
	assign _06957_ = _01569_ | _02097_;
	assign _06958_ = _06957_ | _04648_;
	assign _06959_ = _06958_ | _07758_;
	assign _06960_ = _01875_ & ~_06959_;
	assign _06961_ = _04249_ | _01098_;
	assign _06962_ = _06961_ | _02097_;
	assign _06963_ = _06962_ | _07758_;
	assign _06964_ = _06963_ | \mchip.index [10];
	assign _06965_ = \mchip.index [11] & ~_06964_;
	assign _06967_ = _07588_ | \mchip.index [5];
	assign _06968_ = _06967_ | \mchip.index [6];
	assign _06969_ = _06968_ | _02097_;
	assign _06970_ = _06969_ | \mchip.index [9];
	assign _06971_ = \mchip.index [10] & ~_06970_;
	assign _06972_ = _06582_ | \mchip.index [7];
	assign _06973_ = _06972_ | \mchip.index [8];
	assign _06974_ = \mchip.index [10] & ~_06973_;
	assign _06975_ = _01986_ & ~_02544_;
	assign _06976_ = _05529_ | _01986_;
	assign _06979_ = _01875_ & ~_06976_;
	assign _06980_ = \mchip.index [11] & ~_04684_;
	assign _06981_ = _01681_ | \mchip.index [9];
	assign _06982_ = \mchip.index [10] & ~_06981_;
	assign _06983_ = _04712_ | _02097_;
	assign _06984_ = _06983_ | _04648_;
	assign _06985_ = _06984_ | \mchip.index [9];
	assign _06986_ = _06985_ | \mchip.index [10];
	assign _06987_ = _01875_ & ~_06986_;
	assign _06988_ = _01523_ | \mchip.index [8];
	assign _06990_ = \mchip.index [11] & ~_06988_;
	assign _06991_ = _01869_ | _04648_;
	assign _06992_ = _06991_ | _07758_;
	assign _06993_ = _06992_ | _01986_;
	assign _06994_ = _01875_ & ~_06993_;
	assign _06995_ = _04741_ | \mchip.index [6];
	assign _06996_ = _06995_ | \mchip.index [7];
	assign _06997_ = _06996_ | _04648_;
	assign _06998_ = _06997_ | \mchip.index [9];
	assign _06999_ = _06998_ | \mchip.index [10];
	assign _07001_ = _01875_ & ~_06999_;
	assign _07002_ = _00514_ | \mchip.index [6];
	assign _07003_ = _07002_ | _01986_;
	assign _07004_ = \mchip.index [11] & ~_07003_;
	assign _07005_ = _04648_ & ~_06836_;
	assign _07006_ = _01172_ | _04648_;
	assign _07007_ = _07006_ | \mchip.index [10];
	assign _07008_ = _01875_ & ~_07007_;
	assign _07009_ = _00838_ | _07758_;
	assign _07010_ = _01986_ & ~_07009_;
	assign _07012_ = _01263_ | _04648_;
	assign _07013_ = _07012_ | _07758_;
	assign _07014_ = _01986_ & ~_07013_;
	assign _07015_ = _00796_ | _02984_;
	assign _07016_ = _07015_ | \mchip.index [7];
	assign _07017_ = _07016_ | \mchip.index [8];
	assign _07018_ = _07017_ | \mchip.index [9];
	assign _07019_ = \mchip.index [11] & ~_07018_;
	assign _07020_ = _07780_ | \mchip.index [7];
	assign _07021_ = _07020_ | \mchip.index [8];
	assign _07023_ = _07021_ | \mchip.index [10];
	assign _07024_ = _01875_ & ~_07023_;
	assign _07025_ = _04116_ | _04648_;
	assign _07026_ = _07025_ | \mchip.index [9];
	assign _07027_ = _07026_ | \mchip.index [10];
	assign _07028_ = _01875_ & ~_07027_;
	assign _07029_ = _01133_ | _04648_;
	assign _07030_ = _07029_ | _07758_;
	assign _07031_ = _01986_ & ~_07030_;
	assign _07032_ = _01839_ | _04648_;
	assign _07034_ = _07032_ | \mchip.index [9];
	assign _07035_ = \mchip.index [11] & ~_07034_;
	assign _07036_ = _04204_ | \mchip.index [6];
	assign _07037_ = _07036_ | _02097_;
	assign _07038_ = _07037_ | _04648_;
	assign _07039_ = _07038_ | \mchip.index [9];
	assign _07040_ = \mchip.index [10] & ~_07039_;
	assign _07041_ = _05520_ | \mchip.index [7];
	assign _07042_ = _07041_ | _04648_;
	assign _07043_ = _07758_ & ~_07042_;
	assign _07045_ = _01442_ | _01986_;
	assign _07046_ = \mchip.index [11] & ~_07045_;
	assign _07047_ = _00837_ | \mchip.index [5];
	assign _07048_ = _07047_ | \mchip.index [7];
	assign _07049_ = _07048_ | \mchip.index [8];
	assign _07050_ = _01875_ & ~_07049_;
	assign _07051_ = _00501_ | _02984_;
	assign _07052_ = _07051_ | _02097_;
	assign _07053_ = _07052_ | _04648_;
	assign _07054_ = _07053_ | _07758_;
	assign _07056_ = _07054_ | _01986_;
	assign _07057_ = _01875_ & ~_07056_;
	assign _07058_ = _01842_ | \mchip.index [7];
	assign _07059_ = _07058_ | _04648_;
	assign _07060_ = _07059_ | \mchip.index [9];
	assign _07061_ = _07060_ | \mchip.index [10];
	assign _07062_ = _01875_ & ~_07061_;
	assign _07063_ = _05166_ | \mchip.index [9];
	assign _07064_ = _07063_ | \mchip.index [10];
	assign _07065_ = \mchip.index [11] & ~_07064_;
	assign _07067_ = _02445_ | _01986_;
	assign _07068_ = \mchip.index [11] & ~_07067_;
	assign _07069_ = _06768_ | \mchip.index [10];
	assign _07070_ = \mchip.index [11] & ~_07069_;
	assign _07071_ = _04204_ | _02984_;
	assign _07072_ = _07071_ | _02097_;
	assign _07073_ = _07072_ | \mchip.index [8];
	assign _07074_ = _07073_ | _07758_;
	assign _07075_ = \mchip.index [10] & ~_07074_;
	assign _07076_ = _04135_ | \mchip.index [8];
	assign _07078_ = _07076_ | _07758_;
	assign _07079_ = _07078_ | \mchip.index [10];
	assign _07080_ = _01875_ & ~_07079_;
	assign _07081_ = _00022_ | _01986_;
	assign _07082_ = \mchip.index [11] & ~_07081_;
	assign _07083_ = _05433_ | \mchip.index [6];
	assign _07084_ = _07083_ | \mchip.index [9];
	assign _07085_ = \mchip.index [10] & ~_07084_;
	assign _07086_ = _04680_ | \mchip.index [8];
	assign _07087_ = _07086_ | \mchip.index [9];
	assign _07090_ = _01875_ & ~_07087_;
	assign _07091_ = _01120_ | _02984_;
	assign _07092_ = _07091_ | _04648_;
	assign _07093_ = _07092_ | _01986_;
	assign _07094_ = _01875_ & ~_07093_;
	assign _07095_ = _04071_ | _04648_;
	assign _07096_ = _07095_ | _07758_;
	assign _07097_ = \mchip.index [10] & ~_07096_;
	assign _07098_ = _01889_ | \mchip.index [8];
	assign _07099_ = _07098_ | _07758_;
	assign _07101_ = \mchip.index [11] & ~_07099_;
	assign _07102_ = _01231_ | \mchip.index [8];
	assign _07103_ = _07102_ | \mchip.index [10];
	assign _07104_ = _01875_ & ~_07103_;
	assign _07105_ = _01748_ | _04648_;
	assign _07106_ = _07105_ | \mchip.index [9];
	assign _07107_ = \mchip.index [10] & ~_07106_;
	assign _07108_ = \mchip.index [11] & ~_06349_;
	assign _07109_ = _02441_ | _07758_;
	assign _07110_ = _01986_ & ~_07109_;
	assign _07112_ = _01899_ | _02984_;
	assign _07113_ = _07112_ | \mchip.index [8];
	assign _07114_ = _07113_ | \mchip.index [10];
	assign _07115_ = _01875_ & ~_07114_;
	assign _07116_ = _03985_ | \mchip.index [8];
	assign _07117_ = _07116_ | \mchip.index [9];
	assign _07118_ = \mchip.index [11] & ~_07117_;
	assign _07119_ = _00754_ | \mchip.index [7];
	assign _07120_ = _07119_ | \mchip.index [8];
	assign _07121_ = _07120_ | \mchip.index [9];
	assign _07123_ = \mchip.index [10] & ~_07121_;
	assign _07124_ = \mchip.index [11] & ~_03302_;
	assign _07125_ = _01376_ | \mchip.index [5];
	assign _07126_ = _07125_ | _02984_;
	assign _07127_ = _07126_ | _02097_;
	assign _07128_ = _07127_ | _04648_;
	assign _07129_ = _07128_ | \mchip.index [10];
	assign _07130_ = _01875_ & ~_07129_;
	assign _07131_ = _01619_ | \mchip.index [7];
	assign _07132_ = _07131_ | \mchip.index [8];
	assign _07134_ = \mchip.index [10] & ~_07132_;
	assign _07135_ = _02531_ | \mchip.index [10];
	assign _07136_ = _01875_ & ~_07135_;
	assign _07137_ = _02064_ | _02097_;
	assign _07138_ = _07137_ | _04648_;
	assign _07139_ = _07138_ | \mchip.index [9];
	assign _07140_ = \mchip.index [11] & ~_07139_;
	assign _07141_ = _01875_ & ~_05290_;
	assign _07142_ = _07599_ | _04648_;
	assign _07143_ = _07142_ | _07758_;
	assign _07145_ = _07143_ | _01986_;
	assign _07146_ = _01875_ & ~_07145_;
	assign _07147_ = _01869_ | _02097_;
	assign _07148_ = _07147_ | \mchip.index [9];
	assign _07149_ = \mchip.index [10] & ~_07148_;
	assign _07150_ = _02088_ | \mchip.index [7];
	assign _07151_ = _07150_ | \mchip.index [8];
	assign _07152_ = _01875_ & ~_07151_;
	assign _07153_ = _01893_ | _02097_;
	assign _07154_ = _07153_ | _07758_;
	assign _07156_ = _01875_ & ~_07154_;
	assign _07157_ = _04548_ | _02097_;
	assign _07158_ = _07157_ | _04648_;
	assign _07159_ = _07158_ | \mchip.index [9];
	assign _07160_ = \mchip.index [10] & ~_07159_;
	assign _07161_ = _07690_ | _02097_;
	assign _07162_ = _07161_ | _04648_;
	assign _07163_ = \mchip.index [11] & ~_07162_;
	assign _07164_ = _01748_ | \mchip.index [8];
	assign _07165_ = _07164_ | _07758_;
	assign _07167_ = \mchip.index [11] & ~_07165_;
	assign _07168_ = \mchip.index [10] & ~_03182_;
	assign _07169_ = _02486_ | \mchip.index [8];
	assign _07170_ = _07169_ | \mchip.index [9];
	assign _07171_ = \mchip.index [10] & ~_07170_;
	assign _07172_ = _03357_ | _07758_;
	assign _07173_ = _07172_ | _01986_;
	assign _07174_ = _01875_ & ~_07173_;
	assign _07175_ = _02474_ | _02097_;
	assign _07176_ = _07175_ | _07758_;
	assign _07178_ = _07176_ | \mchip.index [10];
	assign _07179_ = \mchip.index [11] & ~_07178_;
	assign _07180_ = _06235_ | _05424_;
	assign _07181_ = _02097_ & ~_07180_;
	assign _07182_ = _05162_ | \mchip.index [7];
	assign _07183_ = _07182_ | _04648_;
	assign _07184_ = _07183_ | \mchip.index [10];
	assign _07185_ = \mchip.index [11] & ~_07184_;
	assign _07186_ = _04631_ | _04648_;
	assign _07187_ = _07186_ | _07758_;
	assign _07189_ = _07187_ | _01986_;
	assign _07190_ = _01875_ & ~_07189_;
	assign _07191_ = _00268_ | _02097_;
	assign _07192_ = _07191_ | _07758_;
	assign _07193_ = _07192_ | \mchip.index [10];
	assign _07194_ = \mchip.index [11] & ~_07193_;
	assign _07195_ = _03540_ | \mchip.index [6];
	assign _07196_ = _07195_ | _02097_;
	assign _07197_ = _07196_ | _04648_;
	assign _07198_ = _07197_ | _07758_;
	assign _07201_ = _07198_ | _01986_;
	assign _07202_ = _01875_ & ~_07201_;
	assign _07203_ = _01710_ | _04648_;
	assign _07204_ = _07203_ | _07758_;
	assign _07205_ = _07204_ | _01986_;
	assign _07206_ = \mchip.index [11] & ~_07205_;
	assign _07207_ = _00765_ | \mchip.index [9];
	assign _07208_ = \mchip.index [10] & ~_07207_;
	assign _07209_ = _05946_ | _02984_;
	assign _07210_ = _07209_ | _02097_;
	assign _07212_ = _07210_ | \mchip.index [9];
	assign _07213_ = \mchip.index [11] & ~_07212_;
	assign _07214_ = _04143_ | \mchip.index [6];
	assign _07215_ = _07214_ | _02097_;
	assign _07216_ = _07215_ | \mchip.index [8];
	assign _07217_ = _07216_ | _07758_;
	assign _07218_ = _01986_ & ~_07217_;
	assign _07219_ = _01949_ | _02097_;
	assign _07220_ = _07219_ | _04648_;
	assign _07221_ = _07220_ | \mchip.index [9];
	assign _07223_ = _07221_ | \mchip.index [10];
	assign _07224_ = _01875_ & ~_07223_;
	assign _07225_ = _06618_ | \mchip.index [9];
	assign _07226_ = \mchip.index [11] & ~_07225_;
	assign _07227_ = _00329_ | _02984_;
	assign _07228_ = _07227_ | \mchip.index [7];
	assign _07229_ = _07228_ | _04648_;
	assign _07230_ = _07229_ | _07758_;
	assign _07231_ = _07230_ | _01986_;
	assign _07232_ = \mchip.index [11] & ~_07231_;
	assign _07234_ = _00791_ | \mchip.index [6];
	assign _07235_ = _07234_ | _02097_;
	assign _07236_ = _07235_ | _04648_;
	assign _07237_ = _07236_ | _07758_;
	assign _07238_ = _07237_ | _01986_;
	assign _07239_ = _01875_ & ~_07238_;
	assign _07240_ = _02109_ | _02984_;
	assign _07241_ = _07240_ | \mchip.index [7];
	assign _07242_ = _07241_ | \mchip.index [8];
	assign _07243_ = \mchip.index [9] & ~_07242_;
	assign _07245_ = _01491_ | \mchip.index [6];
	assign _07246_ = _07245_ | \mchip.index [8];
	assign _07247_ = _07246_ | _07758_;
	assign _07248_ = _07247_ | \mchip.index [10];
	assign _07249_ = _01875_ & ~_07248_;
	assign _07250_ = _07736_ | \mchip.index [8];
	assign _07251_ = _07250_ | \mchip.index [9];
	assign _07252_ = \mchip.index [10] & ~_07251_;
	assign _07253_ = _00600_ | \mchip.index [7];
	assign _07254_ = _07253_ | _04648_;
	assign _07256_ = _07254_ | \mchip.index [9];
	assign _07257_ = _07256_ | \mchip.index [10];
	assign _07258_ = _01875_ & ~_07257_;
	assign _07259_ = _01986_ & ~_07641_;
	assign _07260_ = _04017_ | \mchip.index [8];
	assign _07261_ = _07260_ | _07758_;
	assign _07262_ = \mchip.index [10] & ~_07261_;
	assign _07263_ = _00703_ | \mchip.index [8];
	assign _07264_ = _07758_ & ~_07263_;
	assign _07265_ = _05273_ | \mchip.index [7];
	assign _07267_ = \mchip.index [11] & ~_07265_;
	assign _07268_ = _03954_ | _02984_;
	assign _07269_ = _07268_ | _02097_;
	assign _07270_ = _07269_ | _01986_;
	assign _07271_ = _01875_ & ~_07270_;
	assign _07272_ = _04291_ | _02984_;
	assign _07273_ = _07272_ | \mchip.index [7];
	assign _07274_ = _07273_ | _01986_;
	assign _07275_ = \mchip.index [11] & ~_07274_;
	assign _07276_ = _03239_ | \mchip.index [10];
	assign _07278_ = \mchip.index [11] & ~_07276_;
	assign _07279_ = _05222_ | _02097_;
	assign _07280_ = _07279_ | \mchip.index [8];
	assign _07281_ = _07280_ | \mchip.index [9];
	assign _07282_ = _07281_ | _01986_;
	assign _07283_ = _01875_ & ~_07282_;
	assign _07284_ = _00263_ | _02984_;
	assign _07285_ = _07284_ | _02097_;
	assign _07286_ = _07285_ | _04648_;
	assign _07287_ = _07286_ | \mchip.index [10];
	assign _07289_ = \mchip.index [11] & ~_07287_;
	assign _07290_ = _05193_ | _07758_;
	assign _07291_ = \mchip.index [10] & ~_07290_;
	assign _07292_ = _01429_ | _04648_;
	assign _07293_ = _07292_ | \mchip.index [9];
	assign _07294_ = \mchip.index [10] & ~_07293_;
	assign _07295_ = _04648_ & ~_07083_;
	assign _07296_ = _02707_ | _02097_;
	assign _07297_ = _07296_ | \mchip.index [9];
	assign _07298_ = _07297_ | \mchip.index [10];
	assign _07300_ = _01875_ & ~_07298_;
	assign _07301_ = _02220_ | _04648_;
	assign _07302_ = _07301_ | \mchip.index [9];
	assign _07303_ = \mchip.index [10] & ~_07302_;
	assign _07304_ = _00884_ | _02984_;
	assign _07305_ = _07304_ | _02097_;
	assign _07306_ = _07305_ | \mchip.index [8];
	assign _07307_ = \mchip.index [10] & ~_07306_;
	assign _07308_ = _03010_ | \mchip.index [6];
	assign _07309_ = _02097_ & ~_07308_;
	assign _07312_ = _05115_ | \mchip.index [6];
	assign _07313_ = _07312_ | _02097_;
	assign _07314_ = _07313_ | _07758_;
	assign _07315_ = _07314_ | \mchip.index [10];
	assign _07316_ = _01875_ & ~_07315_;
	assign _07317_ = _01190_ | \mchip.index [8];
	assign _07318_ = \mchip.index [10] & ~_07317_;
	assign _07319_ = _07318_ | _07316_;
	assign _07320_ = _07319_ | _07309_;
	assign _07321_ = _07320_ | _07307_;
	assign _07323_ = _07321_ | _07303_;
	assign _07324_ = _07323_ | _07300_;
	assign _07325_ = _07324_ | _07295_;
	assign _07326_ = _07325_ | _07294_;
	assign _07327_ = _07326_ | _07291_;
	assign _07328_ = _07327_ | _07289_;
	assign _07329_ = _07328_ | _07283_;
	assign _07330_ = _07329_ | _07278_;
	assign _07331_ = _07330_ | _07275_;
	assign _07332_ = _07331_ | _07271_;
	assign _07334_ = _07332_ | _07267_;
	assign _07335_ = _07334_ | _07264_;
	assign _07336_ = _07335_ | _07262_;
	assign _07337_ = _07336_ | _07259_;
	assign _07338_ = _07337_ | _07258_;
	assign _07339_ = _07338_ | _07252_;
	assign _07340_ = _07339_ | _07249_;
	assign _07341_ = _07340_ | _07243_;
	assign _07342_ = _07341_ | _07239_;
	assign _07343_ = _07342_ | _07232_;
	assign _07345_ = _07343_ | _07226_;
	assign _07346_ = _07345_ | _07224_;
	assign _07347_ = _07346_ | _07218_;
	assign _07348_ = _07347_ | _07213_;
	assign _07349_ = _07348_ | _07208_;
	assign _07350_ = _07349_ | _07206_;
	assign _07351_ = _07350_ | _07202_;
	assign _07352_ = _07351_ | _07194_;
	assign _07353_ = _07352_ | _07190_;
	assign _07354_ = _07353_ | _07185_;
	assign _07356_ = _07354_ | _07181_;
	assign _07357_ = _07356_ | _07179_;
	assign _07358_ = _07357_ | _07174_;
	assign _07359_ = _07358_ | _07171_;
	assign _07360_ = _07359_ | _07168_;
	assign _07361_ = _07360_ | _07167_;
	assign _07362_ = _07361_ | _07163_;
	assign _07363_ = _07362_ | _07160_;
	assign _07364_ = _07363_ | _07156_;
	assign _07365_ = _07364_ | _07152_;
	assign _07367_ = _07365_ | _07149_;
	assign _07368_ = _07367_ | _07146_;
	assign _07369_ = _07368_ | _07141_;
	assign _07370_ = _07369_ | _07140_;
	assign _07371_ = _07370_ | _07136_;
	assign _07372_ = _07371_ | _07134_;
	assign _07373_ = _07372_ | _07130_;
	assign _07374_ = _07373_ | _07124_;
	assign _07375_ = _07374_ | _07123_;
	assign _07376_ = _07375_ | _07118_;
	assign _07378_ = _07376_ | _07115_;
	assign _07379_ = _07378_ | _07110_;
	assign _07380_ = _07379_ | _07108_;
	assign _07381_ = _07380_ | _07107_;
	assign _07382_ = _07381_ | _07104_;
	assign _07383_ = _07382_ | _07101_;
	assign _07384_ = _07383_ | _07097_;
	assign _07385_ = _07384_ | _07094_;
	assign _07386_ = _07385_ | _07090_;
	assign _07387_ = _07386_ | _07085_;
	assign _07389_ = _07387_ | _07082_;
	assign _07390_ = _07389_ | _07080_;
	assign _07391_ = _07390_ | _07075_;
	assign _07392_ = _07391_ | _07070_;
	assign _07393_ = _07392_ | _07068_;
	assign _07394_ = _07393_ | _07065_;
	assign _07395_ = _07394_ | _07062_;
	assign _07396_ = _07395_ | _07057_;
	assign _07397_ = _07396_ | _07050_;
	assign _07398_ = _07397_ | _07046_;
	assign _07400_ = _07398_ | _07043_;
	assign _07401_ = _07400_ | _07040_;
	assign _07402_ = _07401_ | _07035_;
	assign _07403_ = _07402_ | _07031_;
	assign _07404_ = _07403_ | _07028_;
	assign _07405_ = _07404_ | _07024_;
	assign _07406_ = _07405_ | _07019_;
	assign _07407_ = _07406_ | _07014_;
	assign _07408_ = _07407_ | _07010_;
	assign _07409_ = _07408_ | _07008_;
	assign _07411_ = _07409_ | _07005_;
	assign _07412_ = _07411_ | _07004_;
	assign _07413_ = _07412_ | _07001_;
	assign _07414_ = _07413_ | _06994_;
	assign _07415_ = _07414_ | _06990_;
	assign _07416_ = _07415_ | _06987_;
	assign _07417_ = _07416_ | _05796_;
	assign _07418_ = _07417_ | _06982_;
	assign _07419_ = _07418_ | _06980_;
	assign _07420_ = _07419_ | _06979_;
	assign _07423_ = _07420_ | _06975_;
	assign _07424_ = _07423_ | _06974_;
	assign _07425_ = _07424_ | _06971_;
	assign _07426_ = _07425_ | _06965_;
	assign _07427_ = _07426_ | _06960_;
	assign _07428_ = _07427_ | _06956_;
	assign _07429_ = _07428_ | _06953_;
	assign _07430_ = _07429_ | _06950_;
	assign _07431_ = _07430_ | _06947_;
	assign _07432_ = _07431_ | _06943_;
	assign _07434_ = _07432_ | _06941_;
	assign _07435_ = _07434_ | _06937_;
	assign _07436_ = _07435_ | _06934_;
	assign _07437_ = _07436_ | _06931_;
	assign _07438_ = _07437_ | _04352_;
	assign _07439_ = _07438_ | _06927_;
	assign _07440_ = _07439_ | _06924_;
	assign _07441_ = _07440_ | _06919_;
	assign _07442_ = _07441_ | _06916_;
	assign _07443_ = _07442_ | _06912_;
	assign _07445_ = _07443_ | _06908_;
	assign _07446_ = _07445_ | _06907_;
	assign _07447_ = _07446_ | _06904_;
	assign _07448_ = _07447_ | _06901_;
	assign _07449_ = _07448_ | _06898_;
	assign _07450_ = _07449_ | _06896_;
	assign _07451_ = _07450_ | _06892_;
	assign _07452_ = _07451_ | _06888_;
	assign _07453_ = _07452_ | _06884_;
	assign _07454_ = _07453_ | _06883_;
	assign _07456_ = _07454_ | _06879_;
	assign _07457_ = _07456_ | _06874_;
	assign _07458_ = _07457_ | _06871_;
	assign _07459_ = _07458_ | _06870_;
	assign _07460_ = _07459_ | _06863_;
	assign _07461_ = _07460_ | _06860_;
	assign _07462_ = _07461_ | _06859_;
	assign _07463_ = _07462_ | _06857_;
	assign _07464_ = _07463_ | _06854_;
	assign _07465_ = _07464_ | _06850_;
	assign _07467_ = _07465_ | _06849_;
	assign _07468_ = _07467_ | _06847_;
	assign _07469_ = _07468_ | _04248_;
	assign _07470_ = _07469_ | _06846_;
	assign _07471_ = _07470_ | _06841_;
	assign _07472_ = _07471_ | _06837_;
	assign _07473_ = _07472_ | _06835_;
	assign _07474_ = _07473_ | _06834_;
	assign _07475_ = _07474_ | _06832_;
	assign _07476_ = _07475_ | _06829_;
	assign _07478_ = _07476_ | _06825_;
	assign _07479_ = _07478_ | _04221_;
	assign _07480_ = _07479_ | _06823_;
	assign _07481_ = _07480_ | _06818_;
	assign _07482_ = _07481_ | _06814_;
	assign _07483_ = _07482_ | _06808_;
	assign _07484_ = _07483_ | _06803_;
	assign _07485_ = _07484_ | _06799_;
	assign _07486_ = _07485_ | _06794_;
	assign _07487_ = _07486_ | _06792_;
	assign _07489_ = _07487_ | _06785_;
	assign _07490_ = _07489_ | _06781_;
	assign _07491_ = _07490_ | _06777_;
	assign _07492_ = _07491_ | _06774_;
	assign _07493_ = _07492_ | _06771_;
	assign _07494_ = _07493_ | _06766_;
	assign _07495_ = _07494_ | _06761_;
	assign _07496_ = _07495_ | _06759_;
	assign _07497_ = _07496_ | _06751_;
	assign _07498_ = _07497_ | _06746_;
	assign _07500_ = _07498_ | _06740_;
	assign _07501_ = _07500_ | _01488_;
	assign _07502_ = _07501_ | _06736_;
	assign _07503_ = _07502_ | _06735_;
	assign _07504_ = _07503_ | _06731_;
	assign _07505_ = _07504_ | _06727_;
	assign _07506_ = _07505_ | _06723_;
	assign _07507_ = _07506_ | _06719_;
	assign _07508_ = _07507_ | _06716_;
	assign _07509_ = _07508_ | _06709_;
	assign _07511_ = _07509_ | _06707_;
	assign _07512_ = _07511_ | _06704_;
	assign _07513_ = _07512_ | _06701_;
	assign _07514_ = _07513_ | _06698_;
	assign _07515_ = _07514_ | _06696_;
	assign _07516_ = _07515_ | _06693_;
	assign _07517_ = _07516_ | _06688_;
	assign _07518_ = _07517_ | _06684_;
	assign _07519_ = _07518_ | _06680_;
	assign _07520_ = _07519_ | _06675_;
	assign _07522_ = _07520_ | _06671_;
	assign _07523_ = _07522_ | _06669_;
	assign _07524_ = _07523_ | _06665_;
	assign _07525_ = _07524_ | _06661_;
	assign _07526_ = _07525_ | _06655_;
	assign _07527_ = _07526_ | _06652_;
	assign _07528_ = _07527_ | _06650_;
	assign _07529_ = _07528_ | _06647_;
	assign _07530_ = _07529_ | _06640_;
	assign _07531_ = _07530_ | _06634_;
	assign _07534_ = _07531_ | _06631_;
	assign _07535_ = _07534_ | _06628_;
	assign _07536_ = _07535_ | _06627_;
	assign _07537_ = _07536_ | _06620_;
	assign _07538_ = _07537_ | _06617_;
	assign _07539_ = _07538_ | _06612_;
	assign _07540_ = _07539_ | _06609_;
	assign _07541_ = _07540_ | _06605_;
	assign _07542_ = _07541_ | _02690_;
	assign _07543_ = _07542_ | _06602_;
	assign _07545_ = _07543_ | _06599_;
	assign _07546_ = _07545_ | _06596_;
	assign _07547_ = _07546_ | _06594_;
	assign _07548_ = _07547_ | _06592_;
	assign _07549_ = _07548_ | _06587_;
	assign _07550_ = _07549_ | _06584_;
	assign _07551_ = _07550_ | _04076_;
	assign _07552_ = _07551_ | _06581_;
	assign _07553_ = _07552_ | _06577_;
	assign _07554_ = _07553_ | _06575_;
	assign _07556_ = _07554_ | _06570_;
	assign _07557_ = _07556_ | _06566_;
	assign _07558_ = _07557_ | _06563_;
	assign _07559_ = _07558_ | _06559_;
	assign _07560_ = _07559_ | _06555_;
	assign _07561_ = _07560_ | _06551_;
	assign _07562_ = _07561_ | _06549_;
	assign _07563_ = _07562_ | _06544_;
	assign _07564_ = _07563_ | _05297_;
	assign _07565_ = _07564_ | _06541_;
	assign _07567_ = _07565_ | _06537_;
	assign _07568_ = _07567_ | _06535_;
	assign _07569_ = _07568_ | _06531_;
	assign _07570_ = _07569_ | _06530_;
	assign _07571_ = _07570_ | _06527_;
	assign _07572_ = _07571_ | _06524_;
	assign _07573_ = _07572_ | _06521_;
	assign _07574_ = _07573_ | _06519_;
	assign _07575_ = _07574_ | _06517_;
	assign _07576_ = _07575_ | _03965_;
	assign _07578_ = _07576_ | _06514_;
	assign _07579_ = _07578_ | _01346_;
	assign _07580_ = _07579_ | _06512_;
	assign _07581_ = _07580_ | _06506_;
	assign _07582_ = _07581_ | _06505_;
	assign _07583_ = _07582_ | _06503_;
	assign _07584_ = _07583_ | _06501_;
	assign _07585_ = _07584_ | _06499_;
	assign _07586_ = _07585_ | _06496_;
	assign _07587_ = _07586_ | _06494_;
	assign _07589_ = _07587_ | _06492_;
	assign _07590_ = _07589_ | _06486_;
	assign _07591_ = _07590_ | _06484_;
	assign _07592_ = _07591_ | _06480_;
	assign _07593_ = _07592_ | _06475_;
	assign _07594_ = _07593_ | _06473_;
	assign _07595_ = _07594_ | _06471_;
	assign _07596_ = _07595_ | _06468_;
	assign _07597_ = _07596_ | _06465_;
	assign _07598_ = _07597_ | _06463_;
	assign _07600_ = _07598_ | _06459_;
	assign _07601_ = _07600_ | _06454_;
	assign _07602_ = _07601_ | _06450_;
	assign _07603_ = _07602_ | _06447_;
	assign _07604_ = _07603_ | _06446_;
	assign _07605_ = _07604_ | _06443_;
	assign _07606_ = _07605_ | _06441_;
	assign _07607_ = _07606_ | _06437_;
	assign _07608_ = _07607_ | _06432_;
	assign _07609_ = _07608_ | _06428_;
	assign _07611_ = _07609_ | _06426_;
	assign _07612_ = _07611_ | _06425_;
	assign _07613_ = _07612_ | _06418_;
	assign _07614_ = _07613_ | _06415_;
	assign _07615_ = _07614_ | _06412_;
	assign _07616_ = _07615_ | _06407_;
	assign _07617_ = _07616_ | _06405_;
	assign _07618_ = _07617_ | _06401_;
	assign _07619_ = _07618_ | _01151_;
	assign _07620_ = _07619_ | _06398_;
	assign _07622_ = _07620_ | _06396_;
	assign _07623_ = _07622_ | _06391_;
	assign _07624_ = _07623_ | _06386_;
	assign _07625_ = _07624_ | _06384_;
	assign _07626_ = _07625_ | _06379_;
	assign _07627_ = _07626_ | _06377_;
	assign _07628_ = _07627_ | _06374_;
	assign _07629_ = _07628_ | _06370_;
	assign _07630_ = _07629_ | _06366_;
	assign _07631_ = _07630_ | _06364_;
	assign _07633_ = _07631_ | _06362_;
	assign _07634_ = _07633_ | _06360_;
	assign _07635_ = _07634_ | _02443_;
	assign _07636_ = _07635_ | _06354_;
	assign \mchip.val [0] = _07636_ | _06350_;
	always @(posedge io_in[12]) \mchip.index [0] <= io_in[0];
	always @(posedge io_in[12]) \mchip.index [1] <= io_in[1];
	always @(posedge io_in[12]) \mchip.index [2] <= io_in[2];
	always @(posedge io_in[12]) \mchip.index [3] <= io_in[3];
	always @(posedge io_in[12]) \mchip.index [4] <= io_in[4];
	always @(posedge io_in[12]) \mchip.index [5] <= io_in[5];
	always @(posedge io_in[12]) \mchip.index [6] <= io_in[6];
	always @(posedge io_in[12]) \mchip.index [7] <= io_in[7];
	always @(posedge io_in[12]) \mchip.index [8] <= io_in[8];
	always @(posedge io_in[12]) \mchip.index [9] <= io_in[9];
	always @(posedge io_in[12]) \mchip.index [10] <= io_in[10];
	always @(posedge io_in[12]) \mchip.index [11] <= io_in[11];
	reg \mchip.io_out_reg[0] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[0]  <= \mchip.val [0];
	assign \mchip.io_out [0] = \mchip.io_out_reg[0] ;
	reg \mchip.io_out_reg[1] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[1]  <= \mchip.val [1];
	assign \mchip.io_out [1] = \mchip.io_out_reg[1] ;
	reg \mchip.io_out_reg[2] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[2]  <= \mchip.val [2];
	assign \mchip.io_out [2] = \mchip.io_out_reg[2] ;
	reg \mchip.io_out_reg[3] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[3]  <= \mchip.val [3];
	assign \mchip.io_out [3] = \mchip.io_out_reg[3] ;
	reg \mchip.io_out_reg[4] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[4]  <= \mchip.val [4];
	assign \mchip.io_out [4] = \mchip.io_out_reg[4] ;
	reg \mchip.io_out_reg[5] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[5]  <= \mchip.val [5];
	assign \mchip.io_out [5] = \mchip.io_out_reg[5] ;
	reg \mchip.io_out_reg[6] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[6]  <= \mchip.val [6];
	assign \mchip.io_out [6] = \mchip.io_out_reg[6] ;
	assign io_out = {7'h00, \mchip.io_out [6:0]};
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out [11:7] = 5'h00;
	assign \mchip.reset  = io_in[13];
	assign \mchip.val [7] = 1'h0;
endmodule
`default_nettype none
module multiplexer (
	io_in,
	io_out,
	des_sel,
	hold_if_not_sel,
	sync_inputs,
	des_io_in,
	des_reset,
	des_io_out,
	clock,
	reset
);
	input wire [11:0] io_in;
	output reg [11:0] io_out;
	input wire [5:0] des_sel;
	input wire hold_if_not_sel;
	input wire sync_inputs;
	output reg [767:0] des_io_in;
	output reg [0:63] des_reset;
	input wire [767:0] des_io_out;
	input wire clock;
	input wire reset;
	reg [12:0] io_in_sync1;
	reg [12:0] io_in_sync2;
	reg [12:0] io_in_sync3;
	reg [63:0] des_sel_dec;
	always @(posedge clock) begin
		des_sel_dec <= 1'sb0;
		des_sel_dec[des_sel] <= 1;
		io_in_sync3 <= io_in_sync2;
		io_in_sync2 <= io_in_sync1;
		io_in_sync1 <= {reset, io_in};
	end
	integer i;
	always @(*) begin
		io_out = 1'sb0;
		for (i = 0; i < 64; i = i + 1)
			begin
				if (des_sel_dec[i])
					io_out = des_io_out[(63 - i) * 12+:12];
				if (hold_if_not_sel && !des_sel_dec[i]) begin
					des_io_in[(63 - i) * 12+:12] = 1'sb0;
					des_reset[i] = 1'sb1;
				end
				else begin
					des_io_in[(63 - i) * 12+:12] = (sync_inputs ? io_in_sync3[11:0] : io_in);
					des_reset[i] = (sync_inputs ? io_in_sync3[12] : reset);
				end
			end
	end
endmodule
`default_nettype none
module design_instantiations (
	io_in,
	io_out,
	des_sel,
	hold_if_not_sel,
	sync_inputs,
	clock,
	reset
);
	input wire [11:0] io_in;
	output wire [11:0] io_out;
	input wire [5:0] des_sel;
	input wire hold_if_not_sel;
	input wire sync_inputs;
	input wire clock;
	input wire reset;
	wire [767:0] des_io_in;
	wire [767:0] des_io_out;
	wire [0:63] des_reset;
	multiplexer mux(
		.io_in(io_in),
		.io_out(io_out),
		.des_sel(des_sel),
		.hold_if_not_sel(hold_if_not_sel),
		.sync_inputs(sync_inputs),
		.des_io_in(des_io_in),
		.des_reset(des_reset),
		.des_io_out(des_io_out),
		.clock(clock),
		.reset(reset)
	);
	assign des_io_out[756+:12] = 12'h000;
	d01_example_adder inst1(
		.io_in({des_reset[1], clock, des_io_in[744+:12]}),
		.io_out(des_io_out[744+:12])
	);
	d02_example_counter inst2(
		.io_in({des_reset[2], clock, des_io_in[732+:12]}),
		.io_out(des_io_out[732+:12])
	);
	assign des_io_out[720+:12] = 12'h000;
	assign des_io_out[708+:12] = 12'h000;
	d05_meta_info inst5(
		.io_in({des_reset[5], clock, des_io_in[696+:12]}),
		.io_out(des_io_out[696+:12])
	);
	assign des_io_out[684+:12] = 12'h000;
	assign des_io_out[672+:12] = 12'h000;
	assign des_io_out[660+:12] = 12'h000;
	assign des_io_out[648+:12] = 12'h000;
	assign des_io_out[636+:12] = 12'h000;
	assign des_io_out[624+:12] = 12'h000;
	assign des_io_out[612+:12] = 12'h000;
	assign des_io_out[600+:12] = 12'h000;
	assign des_io_out[588+:12] = 12'h000;
	assign des_io_out[576+:12] = 12'h000;
	assign des_io_out[564+:12] = 12'h000;
	assign des_io_out[552+:12] = 12'h000;
	assign des_io_out[540+:12] = 12'h000;
	assign des_io_out[528+:12] = 12'h000;
	assign des_io_out[516+:12] = 12'h000;
	assign des_io_out[504+:12] = 12'h000;
	assign des_io_out[492+:12] = 12'h000;
	assign des_io_out[480+:12] = 12'h000;
	assign des_io_out[468+:12] = 12'h000;
	assign des_io_out[456+:12] = 12'h000;
	assign des_io_out[444+:12] = 12'h000;
	assign des_io_out[432+:12] = 12'h000;
	assign des_io_out[420+:12] = 12'h000;
	assign des_io_out[408+:12] = 12'h000;
	assign des_io_out[396+:12] = 12'h000;
	assign des_io_out[384+:12] = 12'h000;
	assign des_io_out[372+:12] = 12'h000;
	assign des_io_out[360+:12] = 12'h000;
	assign des_io_out[348+:12] = 12'h000;
	assign des_io_out[336+:12] = 12'h000;
	assign des_io_out[324+:12] = 12'h000;
	assign des_io_out[312+:12] = 12'h000;
	assign des_io_out[300+:12] = 12'h000;
	assign des_io_out[288+:12] = 12'h000;
	assign des_io_out[276+:12] = 12'h000;
	assign des_io_out[264+:12] = 12'h000;
	assign des_io_out[252+:12] = 12'h000;
	assign des_io_out[240+:12] = 12'h000;
	assign des_io_out[228+:12] = 12'h000;
	assign des_io_out[216+:12] = 12'h000;
	assign des_io_out[204+:12] = 12'h000;
	assign des_io_out[192+:12] = 12'h000;
	assign des_io_out[180+:12] = 12'h000;
	assign des_io_out[168+:12] = 12'h000;
	assign des_io_out[156+:12] = 12'h000;
	assign des_io_out[144+:12] = 12'h000;
	assign des_io_out[132+:12] = 12'h000;
	assign des_io_out[120+:12] = 12'h000;
	assign des_io_out[108+:12] = 12'h000;
	assign des_io_out[96+:12] = 12'h000;
	assign des_io_out[84+:12] = 12'h000;
	assign des_io_out[72+:12] = 12'h000;
	assign des_io_out[60+:12] = 12'h000;
	assign des_io_out[48+:12] = 12'h000;
	assign des_io_out[36+:12] = 12'h000;
	assign des_io_out[24+:12] = 12'h000;
	assign des_io_out[12+:12] = 12'h000;
	assign des_io_out[0+:12] = 12'h000;
endmodule
